module testbench();
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    reg [31:0] src16;
    reg [31:0] src17;
    reg [31:0] src18;
    reg [31:0] src19;
    reg [31:0] src20;
    reg [31:0] src21;
    reg [31:0] src22;
    reg [31:0] src23;
    reg [31:0] src24;
    reg [31:0] src25;
    reg [31:0] src26;
    reg [31:0] src27;
    reg [31:0] src28;
    reg [31:0] src29;
    reg [31:0] src30;
    reg [31:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [36:0] srcsum;
    wire [36:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6407c9b3e1030cf3164d10ea5d38e795b884d627d59ab7f7fb73b8882f40338b7da219f40231063b6baf62af61366ddf25f29ebb9e69caaccb904d7dc4de007987952531b9593c9bf00ac67a11d556b0ee842627d7ad0bb239d0ad9f99155fb4850c8460b01c17d852571beae8ab73e9f81499c7f50dc4e935f35a5b0c721863;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e5f9debe34ab6e80f9093267f438267b36dd8785371faafc62f141bf258bf278bed281d49a4f638692b5e815f162d53bc1b26be5e426f43c86c05fdbd05c24ce8e252988970b3974a021c0a1d51555fccf186bc83c22e96c02de486d1ba6015b032fe230c213b2414d424520be54fe61ddc3dabddedfb175f93d79f8bf47556;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a9e828ca38a6e42a0884064773db1e8f206827c3bca855e5cb39f1d845cf5fa3cd938d7db9ad3dd35d3107e883c21fbb425e0dde4a60b23fd873595a7f6dd6f118dae224c3a7d0351af5d1d611e683752b1e4eef65a176fd733acf7470675e4c93630992b0f51dec8915c97ec264c052fdfce060b0ce41ee0df9e0990a61820;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f2d583c51df2bb16294b831b6784827e3b3b2c4f2fe40bcb9e6b22151776b370f1c8e6f59f3934c38bea95571cddfc58efeea95b9f89163f5bdd649544b5d68ff83c422a31266d45ff66f4e8095b4a670e079f9c31afdcb118bb56ce426cd21fb05f3d0310f7bfca9bb9202f72e5de9918c05875562faf1b8b2d918d3b92e11;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb328e5c14374a02599077ca534ed589d7bab454114b29d12f53dfca651fe3c8ca45babdd83dd3234809f898c06ac0baeb13c7ef7842d18a2c12649d769dd6d091d95ee52c9fa4aed8220b378c42cd5083b3da6b095f931c2851376012a3cd7c5303db3d23c8c23caed8f1c738214d104a6a1aff24607cb8c574fde74a099f8fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a54e6efd6421836ee636ea70952997d72d360903266b44f8dea06a4a0c5a8fba885406b4f28912bf18ce55513bf077c7cdba799f99889f75409d32d63eac5b359c8c719b83472508e2aaa7a0d70a5fdad1ad3cd7ba6afcffdb38425ecdbc8c11a99693188ab300141b763ada0bfdaa41cff34f83a55519e9f0e37cb9b8eb6f4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb55bba6ed317553808dd58f29eafad1f9f42e05d98b85759fe90640c5d120270305f692c335a9fdde148f6b4892e9504c22b92be8d85cdbc42a8e49703ede1da5006be9653ebc7c5be6bec89753526f8ea28523c0fc63eece3c5eb4a25376cc84cb930be8f50629a52acf42280ea3fe1ddecf1bf7d995d005969c6d70c4a3d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2b1d2f218a509b6023eac835e10e57684f69d659b1b576ea0578f59fe0f4ab62cf3ef15186a2743a3d3a0b31aa1db16668b790d8c7d8193086a307bfd46ade56155269c39be66399674dbab9e966010913b533a063692e3f1965cd5b9e6597973dfebb80c53f5fd1b7ab816817c3883890a2a28ae52b5e73b787e7996dfb58d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h572624d427c8f1c9a784cb942f018765cac461ab482e258134038d0e1bcc9b8fe85dd611cb228797cc88bba0f8b85118249a273b010efddf83d6cd63c9f91c18a9cad10077b41adf7b8f39d29a1b3b9af252497e45820bfa3a77dad176d1134ef80281a9616c316f7403c2d6a964332ca991d4d1689c11a03a753b3f026cb74a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a3e3d387a7158e99f0a395ac3b4f20fd2f1382c6618bea1ee4230857412ffc00e6c2a93ca4151b1252664ae8732ef7f1e99615f92b6d95b232296dcf5ddef9f14ab3e4a799e8e0ce6d953e2ab95fc6c1543dc3534c5ef653d76b3bb1a901907fa128b22a222f2dc3cb4b7dc818d5b4975f07174bb25a6300d43feaf1dfe8a70;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ebef178195ef07e1e37b4c6238af83f91345913580b9df9d46c49673ed0aa6e27601e41d44b66682609d52b1a8666611caa972c33e8ff056a6cbdbc4076e5abbf6a3a04776db5a16b6490312fcc5d5ee57d86dea30bf599b725c69ddb7f275914ed6de4a995fe3f178e8042d09fa1e1338cffabe2c8e0fb63c0e9adb45d9bcc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34b859b9377ca265ab3d9e2c42444bec4ac2ef2ed10f85d83cd1edd88d125c22bf557ccabc80687690eb3842c87d2ceb6c5433a8c5967f6dc9b6062f3c071fae458f67ab1ac1af5a2ee9af839b788764887896556d592d3a90ad231c5f96285a71cffc8ee333fce434824ee75088021f2970219e5b47f8fbc81916f718691a2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4659347916fdcbffcf9bfa1f09b54189464126d243e27182b6ae2b8a272c8f1d542f676d49bc7b4a06dd7b4df631391640ea1df014b40a1deade0010381df1986671be2954500437d29a7d46c18a4c5af905da88c77c463b822dc506477e8d3a994f0481d4988c1bf315c177e2e9bd357708e5ae59497e9a2c832339274384d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'habe40c85d933a97d4f20aabae035844ae858e26bea55b77438c2e872cebdb10c568e545ed24b8c05a26c6afe5f8ebec4480adaa8051c4f8834925d5b1a7ae29db3fa8a84acd27ea385ae41556783974ccc81f276b7f0322f13881e1a6bbfb522a27ae26f9c5e642c02c58cf9d2cf079098e7c22532577a88d6ae7c36329cf441;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62a5d7a0b4eb20d6952723d427224b534d31d14bd9219b5d0c949422c9b0480e065c729e9f7ac47d4e09129e1c48298e5a614081c31e5f6417823d76d6bd9e1eb9a7c9daae8dd90c2f357757c3c9292c7f578fb17f45b0a1721f4284c824f7e78c707112fa6b5de28a28e94fa65b532cbe738a9389fad2c3e58622c496911667;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h842d2847b54068b5ee00caedebbefbe270f3a69316ddfc0aea9877a797ffc0f8d779602b35aacbee99d04fb534cc0856362c8aee56615d015b8b9f8f83987a564c71c400407ea4b90a3e74bb8af60bed57d855be033bc2b223a3c8301349ec53f08f41ddb92fb91ae6f208de480def31be1a73ee031532fa70f8922f40166141;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfcffe57df7221cb56f270f1ad31df002a98313a5e1211fce00e3019e5a18ae0218c84123b39f553eb173555b00b6750d1b40114b6118eab9e0b4850529a8d68bcb0d55db8596aab5967385dcbc83261dfbc24ccf3a0ab4d7bec13c091cc35e648600ef79cf99bf92254071c1d3e33375fb74d17cf1563e9c242c545467f6d194;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85c797f62d8f214310706a9e62df1fe08c478dcf98f008578b190bd1f7b02f7b05dcf6404b20d6be2f4a4db39aa8fe231578a14ca6cb03d33d940183dd104676d7f2e6293e65be2d9fe648450cc2997a0a3a8bbb2f02d2ba150a52b7925cd334509f9c62a8e7f376414097400378be51dfeb109d7d527306a52e1a3c35521b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4a4883898f634d8eaec2317fc345e221acc1937738382ed8a9fb4365ff285b3f787d780b1c3e82652a5248c4f823739b9995e536232ad57708409e44cf34968799a27efe4e5fec9c023df5824facc5c2fabdef53eecfaa434cac20114ed457f9ea07bba32b14e0f3fd293f4baa6fd8c4ed0c6ce0a277138aeb85f82bfefaee0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54a184a40db9bb82f4c3351c04aa0bc9e318a0fcfe3a6ec8ad65ad91f521e135a144df94b04a108bca2bb6ae5be4acaaa17c65534bac506ae2197452db643500fad7520f9b51cffef25225088d1cbf920bd1962010ad9cadbde74552df734ceacd60410033f5b1762e54d9bcad7741438af58aea930f85d778838c144c7bfda7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc31526194e371cadb96d01bb01a78dcd894beed820dfb1c1e2734e583475a8468f96e76ed1d346e65798b849234f2b977c5e66a179dc32440975ad66cfde67567bebd1381c5a74c6bb965858a22734c1593f5c1d7f3ea869d9c1ccb62b84c01a7a1701961d9b9c9c766ae506b1631661da087fa9e238b3b7da532c752f3eee0d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86b57ca6733b1da5fb1bab483a1ce084d12a7de10e67a232accc032b52e7e857c851f183e8cecee4c69044f14289803f8547d89b78069ed1cc82223e61a3e64450add1b91830689d6f94d42743af159ade101bf5319b666a6c6988fdd3a52e782579258bfcb3d11e2a10c0f3fe853bb6c9e78866107b10fb431520f5fcd634e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h956486ec8ef8737ed5c12e17f4c062c08365b1c1466634062553a0ba15caad5b8125f949677013e07dd796bbbb607b7b20b895611c2199c211996c47dbc3f2b3106af2e04e3695e6db4ba022a41931760eec736045459216e562d528172335a601aa4e4374b22132340478069b48221705e1e3a5fdad9c64a2f231cb00377ea0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46fc7873b12fe90a367a1dd852299c401daa8b3d765fcba714688c634a3c3f5e88f64ed7eb3a84b162bbee287eccb6384307fd5c101024079470fc4cea4c4c183218d3e3f99aa235752574fa34d569cdadfdd4ae8af294cde765fb7f968815985f3ef49af544416ddaf31e0177eff9ef8fcb7df3b29210bf8d612e6b8dba0719;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h583ce894b4d54dd419b0e74438aa2d389638fda1a859b4c0742bf61a2281ad12afb4963667fe79997d35f3f12a6c5259daa03147fc98f72d69ad78b080e35628096e8672674929172d9e196209b9f0d7f9ae93b00bc9cb4e26a1ffecde7d731b701c0c1b1e2483b59e6bd9c28e88ad2ac5ca78174cc3f6c0251b68823f02d5de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f2f475714527197625f88bfc5b36c6e58101df25828093782236f2532523b040737d81e45b3e4ef90d001ae8ca2c08b31b62286344dbe56b893804135b61c680542abf1861ee1bb79a7646f682f78c9a8f14ef469af13365003676fb659933188deedbb019d648fe214259d1439bfcc8fecba83cce6b82ad9100220504b8a2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc35fe8e05243f6ce2b9b894dbec642893b6ae6e4f96e72d674823aef74ecd898740b52b2fb0f8e0a846e35a460178a11604595098b93fe365ca9dc12939f9478bf4a008b932d932cf908b751b860298e8f5ad3c6cef988ab08b6c1b083743e16e6dcb146889f59bc567b4de02ce2cecad55797e1fc6ea52bd1f670bfd678c5f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21baa420d2aa7779a71487dd0fb9f63ac09863224e6213a2daa896732ced0fef0a60354409253a3fc2a376d9ba3c7bb9a59f88fdc3b1ac71f867ac84caa19d0f3959a3d8d0c51a1f931ba63485a2efc90ce0559032e40f129c153857f0c7b7b17352b9033be1a7c6247115aaed706f0dbba7327c2a6cdf3656b87313218a39ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha8e15a421bf7a32307a120ea8341cc49b4300b5490328917f5da6876bc28c0f2759e890ce9d508f228646e14ab1a64eef9914a44da024af65f8097d6466440e427dc5047e205664400b775c63fe7c7362aa1d8423bdf9b00c8045532c60dbe89c7b7cad27d9b6cd836f9ad74cd62b909bf079add132da06a18633c172916e2ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'habe46794cd1a8d304fc47d3a6b38084abf3b43b4bc9b3528790074a7139ee2144fa167d93a9cb100c8b979e0e35c43943783608d1ccfea55254055139ee16d7688f1b5d72ca2996b3c5d6abe8338b0ede059b32401350d334e22cbecea88ad999dec2ee223054974a3fd048e8000f8deb7cd4da91fb06d6fec81fb4a4414b484;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c7c43229dec8a4f848a41961d2886844da8e984a433301703ec3b40a1ba4840979296defa5c6285bb2b474fb63afcc87682ec210569e84d415c102f07b3fcf0b44c82d7f63337c2cda47c4599b842fb8f466bfe0e89dd1e4ec5485d68cb4e2905172b8fc43389f60342e91d96e3d45c15833e742025bb3e504c897a9fbe1c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2938f02ea8ca9067d80ea0776152a4f9b79a620e0f080065dc5f8e59f4b878623e09e7619d9ee28b00edf53dcb3b7919e1168ae9f62eb45d9445134b0a247fc7ba7dd284bbf9e4310dda805c936ca51b9b9a9a36392025f5a2efe3291002708079645c4fe6fadb3852d8e4292ebd1c18921aea6b5c2004380f8a53b0021bd5c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f068f9badde6d3f72b13015b1f48a445ee46e748e1810e897c974e58328d203fdcd6bb818fd5c806608018d34023e5f67110b802515c326f680e24f00f67211cf9c3bf7db87d8f35f08734cd1f16366e5ebf0a9be83a7ca9cd79bea98e35a8885c53f3233f9a4bf78e923224dfc4bcf235e342fbef828432cd0ab0f73163c3b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h149f5965e7ef12ef38a7958981f2720a239547ab9d21408a9cfbd9cae35980bcadef9c4bda4e7bbb4bc673e7804111e8020e7e2e02a6e50137a11692e8d4a4c676a8b198ffa762082c44094254ccaf9fbac6310c016e07511430b9fea7003e39096fd49a2013043068e139f813151411ef988dd195342cae8e17d482638b6c01;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf8334354f55d60bef4f97808e8eaa6bc41dadb42e1aff8137763d85942b756f64d1a280eb37ee4143a3a72bcdfadcebff5af01d276b840b9c75bb3013477b6df396e15476c75c0565b057c607f82d8dd9a8015c963cf17b98a06c451c936ef093d6aee9f385ae389287de1e7e8cc1aa867c0c86b0af408124160f67b5c9bd13b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6eec281e4ba5c54c3c1bca54e92dcd01ee70aa9f682e713d5648e685e0b012f4fd3d59fbd0a8c95fadb993326db06a9c54e63a9cc12c6dbf21dfe31683c3c43bb4f1eacc414547181d34823157ad46e16bd88ae6c17991dc9e389f2f806e939d36985bc7f330a44d7eb327c5cdc17c1800e79fbf44af45bffe8876ca474e468;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdcfa30deb754beee4eb60d131b6b8d46dd0f8fabcbc581fd9f4cc8840f2f8c1558130dbcf7af2d37ef5591796731cd0e31da8f029c1888365df7660cc5a7e42d1b6e83a9ae5c26e1f5c7b857714a35040562177c217a1f0ebb710f9ad69093001eac6a44529fd6d13d54a8003028639ffa162242dc9e1d26456906dd00f52d30;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5b8cc900874f554d4c422547e2a97c39467b41c47a2dda4464d246164bec3d84722026bacee8a37f51cdb51a9fa77f697ac9706eb5a118155f440140a6ed60b9e82e02f2f097ef75bdcf67f295bd9362f17a3c7070817620a71e34d05fcfdfe5e0f81bcfc1f8136c43fe3596fd0071d89d2ef31bac742bad957190572a752bf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8526fd97a50000d92dd17f7ea3ce1df622398efcee3b68a671f15cb4028f2737f969a382e95e7fc9b2cf97bc9dcf883af9a87bf595e3be29fd8559c8fed9ec797ce5a2a2c2f2cd8c7ca3464eff175504092fbb476b785995c182d5762eb231a991f702bc0373da15b8b5ccb26823c18f4a999f0e1ff67ca0ee066a4db2f3daec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc256e4d8dc4b451c2d5ba3e50bfae980b05dabe50cdffd95b203702120a89db0092abbdeecb1e8a205fd867ce6679824f6ec73f13117667d081bdb69a267b29b7869dd6e7689008c0816b02ae7c89753787dadfe4a05196d1a6f95a3bcaaff4a52f5e2e01748368b636d7ab5c4eb9b49c6aad75f84a25e00ab6f6655fdd279a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea59cd03a073ce5c1147372b65fcfd71059cac8c468d899bdb5d477905433bc257a0ce779922239f8c0a790869878a86b95d18fbbed206dfc5faa505caec42f1169e91705322364e0f09f355cd7af6a74347c8199448b99eb91c7f29c0f3d8af67b857a32667acf735ee5eac7743c2da85a6b9390d3b57a40eac1ada188c4ea0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e901adec9eaf14b50059528a55e1c9130e2bf1e35fb2c2f4f13750038e2a54af54bf63ecbc500e813cd3f4b61f878433b8a2dd2dcbe7fb0c973fa3e6e1c992169a59b1b5134ed705dd6673289f01ca2a1aec652c86b79c6c71cb5d11aea18223df2ae8f5f508f5b3d6dd3a0a6c068451189ba53cdbc4071f2ff0e4eca99db89;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h247f4377172d560f3e2c6bd01d536ca23c8e3351c6e21ab505801fe827f6cbb419d03e441f7800c6a5d3af5fd7394a720aedf84521a79dcefcbe7987d72668696cdcad389cb47ee39782710bb2320287695c34e299facae2b3efa18d7a03c4302f9f825ee68a32719fd17f257e848c13d36452ab8aa5189bdde0745cb7158bf5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8b8ca80bac0b7de8676cdd8c1578296809b8f9b31955b365df79d111c4799e80d4860d4a98b990fa755a2561ee8204f93957cadb344977887d38fe86128b65f2e338c352aaaae43816c3dcc7f0d3e6334ad052f9be860ef7b83f295eaaad52054d2718e9aa3a7a5cd01b412b76c52a002474cb2a5fae69c4af256384f5f1e67;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha8209642034b462ba5534892c3e947eaebf74fa10435525f0fa4083e2a480eb422e96296bdfc8564ce25284102301480e7e7a76e3b839c347d03a2993063fde804edc4a04fcd52c1cf1c74eefb5d9b70090134eb615b7c6dfd5c4b0819d19ad092e3f0819798566cfd0505be6c265df9e6b9ca0b9d57078c91bdfaa23ebede11;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c9a0968e5679e4e2c7b858a0e8edeaf2b3a4dc114e6441d0b0cd5352d1d7f63f6fb36866feb02645897fae593d8ae35ed5aeedf3a7799fbd8d1d314f3082d574c8822287ff3190c44fead2b843a2fbfe803f8567b7ec86a976e34379c5385faf758c70706bc386ddba10ba6c1cf429c53f8c4bda1d99f49d6be2b93d9ce0e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3d67a61b29b0dd7fe51fb2cf16bebc59615575000db5563312be89e9fa31a21f3c8cd01bb0c5b50c864bd8136a3c3477886d85bc9f6007c57adb7150476c2fb3a4b39f1ae74eeeafb4565c3df86411105b73ea531738dce225c2c9b17e43b9f0f9b255c04c103dc2cdc5409918736e5d14f0651bd772ad60b840ee92bb237c1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13fa33ddbd407a166a9f309ace8abf498bb6632a4bbcafcd9d2693c3c627b4c528fb9b7ba2434e7b04116bd72577c92c4afb03050ddac63b2ca87f411842f530654664eebd94a7d4bb0265897e5821da5af1fbb6d7cc3567e4c438cbbf6e18fc1f9e294d150868526888a78dd38ec71cce22b5767e38bc444d701644ff9e92c2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h163d7013a7925aa1e18285484901ec7d4de4c5c7a5baca7f6f0338d980a83729256d8a9cdbb748e5aded825dcdd72e19368f028ad7d64404a79af441769fca1c4dff4a1bc9d0e5d94f1d593de95433807d61a9e73161750a716826b404bf9bb93f4fa5faef30533c005a7b89060dd54266feaa0b3f9a23cd60af0bffa0195943;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd99f47bee4202755b2ebdd09963aaa3e2856ddcc54dcafd4e37f31fde55a6eebbec8063311f6f37050c717f7dfa2ca08c9a1ad25155003573cdea7f72276af6c8f6c6a0176e8a3b54cb06bd32fac57585e08655217ede05bb68df2f2d63970dbaa652c46a4e952df860fc92df61cf46f79ebd01c21b46ed21957a8c974795335;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he2bbe76b8b3c77a6e6b909dc4641bcb58144cef9fd9d16c86e1bf1eb5235e1ec1e87f61f97b32bd01727c2e7a3eb06da04393c65c411340bce4adf1c96a19bddcba0b8a597851db0b015f76c2d2885713088c3934232a0d6b08a0ec1cd49a73e19ad70182701d0075794c5316b5d8a3f620a2ae6a691c2f0b9d0a25e933d2bfc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h572c2211a205ad7231749260e627b60ddb0253aa2186ba2c44693bb4b022f4a9b5919e403cafa74e7c7487e3d38f361a11793d22e0a8913668d42c762d608a22f2c87fd440d893e8fc35e5c7e79156a964096424b230cdc1e39afca3191e3f4d620cf007f0ff95cbcdc89624c7f4dde4a26714aecc1fdef20120c5042e5a8492;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1b42ceb646a4ac7bd9d5c02b2ea664a039d3ab75fec0991c42184c974f65a40fd315ed231f778e076d52e2ba50a958ce221cc579f8b2b128e90435bb611b46591258358cc51cf19d181348d8bba93b3f041d9a1f5ada6dbffbae049e1f70706160222dfe2059e5fa1fae2515c76739f8fe891eac392042c902e730fa91f29e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55817c041a5c6ef563a261f254245514df33b9dec6c4028f185eacba880adbffdd0906fbdf3154f813b67b0d1f63f745fe8331035bc7e56f8469781f5f672e4978951ac03e837b6af2984628b2c04ff04e9e536e9e2ce1be70c4a5df5fc1064aa5885cf2f6a66df097aa16e90f0a5267615c17ede507508c71225d1b939e7b86;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43891ac92588897a55f12d9874551982922c8fb338e5073318bd875346890935fb46584b0eb23e0ae8d943cfccc6f04bf22dc8e2c40f768191cecd811ab629d20c8a473558a9499074d6c869bc5179717cc9804ec70656c3a684ee5a161fbb80356cd38e4a89094db9c5af128587bce374f9146bec3a59f441e370b5c395df1e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8454019ae0adec813dd9811bcd0c4d3197621e48274bb5905b5846b7d3d0c036d53dfc0fcf665e7e62e62034b3ceefbfc6be73fb0a55d4f905c76f0a789a372131ce4ab25fcb87aeafc02405509a8d2f1d3da758fa87a20421c13bb3b16991265160869a085d4713d62a378082af1f1200a2823839a61febfef1f8f526199894;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf141fcb4ff0dfb02ba6b12e654422c1db9e1ba1aba894c296b2ce35276ef1f146ac2d564848df5b66dcf1cdff46fc473d081c501cd2201d9fb9ca806a496662166e634e3fd1b00701376c93542820a6d6b700397f75dcc1fba556e04400ec886851024bc1aae9559a55b924cad2931d325d5aff83699b18773dbdba5451ceedb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h703401d2588621ad555196ef03a76fb5310bfcb3a044dfd4d7bab9b32c65f27dcd6294a87bb4b3bcc8206cf944a700471d393b6714c979150adb9907810787c74c70a6530ec08a43ced1b5468f9b7400f0d5aff76c78aef725644899668548a6ab5fd3797a8988f32f0459c8314fe3fe21d6fcf98e2dda079032d79129fee4a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h249aa75a67e1f892da063931140ff30397e8a19dbd7cf20e76196bfe1184ceb810558a2995ef5103366b50381710d70cf266b0e459dcc26946a1b27587af8e4ac8e5207cdaaf4d90c8c443ec62b17f4d133cef958c46314b22a39a4fc8b444c8ba48ebdf616dcc70c269b90f1ff1a0f2f9e6236637c65d52a7a4c0026de1af08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3d44dd44f8bb155ce86bd7067738c0c2847d4befbd4da50f86b5f2075a9d20afdb780d52c542f069965f534406dc5d819330de46a6450e89c7d9199f3f7f7d9955e24810bb085ef945114a339df9ccc8cd82646700cf41248e3dcbc7dbd2c8fbc6f6be1a5bec0510ec89fc0bea2e3a4c3d68fbb34879924289d69c6b0c0e15c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h922e5c250287919df022a9b8672e3353aac486aa9f580a0accef4a877503b1080802baad4947a05b3115003d690afde888717b0f28f45b6e0566e3beb06e9012e86cc4600f251c39a71572fcabe3f8bb5b1efa1112fdf9be610f4c7ff7bbbb34ecd3ddedbed0d8143f67ca89e4fc689f60609f81e62918641d41f996aed6ba19;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9eb184e5d7e5f3904a61e9d3c496920f8bbc53da593f106e99583962a82182dc6d2d804d9bb73896c85cd2b41e9a36f0cb7d4668f8927306c5c54c1b514cca2ffabce48f0902c4acbea953968f9f54b8741d58e96eca9138b6b5293405b439131090449a77d02c7a1cbc9100b076e7838beff31f9dbfb2a074da062ca1687852;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c64b10ace518304fcf7ae80c931ca87f905c101d0c27b3d27b06243171a0cab7f531b7f9e2dd0056e6d9cf1c7f5d90bf0450fed097831f6c34b0f137a1631ca96e1ffbdc9a81b75d4f9abab825ee79616f8983a431110d02c38e6e7e6493b09bed955a94cf4decd79b700d4a18192657fac7726d240914074a883dd3340ea9a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0b280798c04675875ac62950c520ad144a71da8d41e0a49ec4275abf9cee2c73c8d6c37e8ce73b03b31c508cfeb7b9520015da1e9756160ec4e4752cdc592cefed182eb169eb7781efc6907273c6f94178216969e73bf12ded7d446631c91fb227062b883ab2b6353ec113bfe54c0bcfefe1e150bb74ab95c3e783c3e6d4022;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcdc150efe1dbb405e8e970fcebad8a40e6fa85de0a0684210862bc972f69d7b232540c0f1d17e4386b4b731e0aabe403a231f1c8500fd91acfc5228f20c30a7576b370951b7070f0bcdc9364e3f0f1b611a41c7b05f216eb59da17f5631ce6406662d5ccc1a2df32e91872129b2023acce33acb46370d9b713bac03be6926ed1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8d505d2b3fd8ba60993fd122b1c135979a4c5aa62065c6adc04a76a63e9b4fa5a02d74d035c514b8dc1a6b85131ff417c408dcdbaf0116fdde43e9c5de77785cac1a9b3e66537b6f26619fdf5c2fc94f8351fcd10038be89b59d8c204869f2dbadfdf409699cd6fab4a41159704f98b2f094902119881485f637803523668b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6cc77eaa64923f20e68d7ccf8b2a49a1be729cd824900dad87b974664e8f85e44f56e030ddcf03ed68ddfdacd84475dded3506048f69800806856211eab44e1f63488754819dfbff3d77a20abf44046850a19505fabc972d0f0b26ee766568cfc4b601fff238c8ca3d38bf1f05ff40df7a9fcca9f7663edcede1d8ebe9e15d6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3ac31d0dd7d18e83810a0a05361c9a55c2835bd8ebfcff6e831bea10911ebf28046ad2a1cd1140608c08e8582cd5406aada7270ed5ec31db2329619830522fc031b9bb7bff77f786f32f804c39f353f22dce2090867eb45e073063d0aebb33b95f3325b7467db51b93af316896d930cff81c3523e0687ad60d62ca1c872a8d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc66d8bc10240a77886758f19d02ab72bd520d3b75758839efd848dd94e8ccacf19cd00c81b1ca6f4724cf573ab35139817d3b22ff788ad815934b161f6498307cdb8d2e66d8aff866c920e7b95bfa3cfe63fd69f186bfe4e6237cad48ab87c7bad2d18292bd5c13f2658b43e6cc6b97daa3750f1ce1e42d71668e1eeb5d9cd5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had6a924ab8175a74e5c4649afeaf89c828d53491620452a8a545906055a7a43f605b3fe2b71bd774363d251304567733e0f5f45704b6509b89655cf8f05059d3bf69f0c6fba39ac1fa92a31d95b84968817c7474f5a36e375f8de05acc55f752e76b69f5500b41a5dbf86b85c83dca90514c8eb2d6e959b12ebd39758079e0ac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d60c44f467576a915a5c2552babf9480e2921ba501336c3bd8923854135389fc92f4e0c370aff8e3d439bace35d87babc1f6e9503805db0e2d2f209b2e309a9e7a9b63787ce42493619b999a2fde34ec1063df69bc9db2552e2f000ead322b1957547768bc8e6933b4357da1c10bbac21bdcbfdf1f1c765e1da3050d25aa80c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13b9f478a03c39b50f65d303bb1b0fd12330678c39be1f273ad909134118ea7d9ab99cd15d15b25a5d8cab4a7ef29f5289f2c538fd16340156442f860042116d8873327f9f20f1907d091fa3f323eb9a3cf2d5279865ce7ca031202206179852df23d50948b4b36998e263dd86c8db88bf9a565efb2f1ef556b01c1613c0553;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9670ff6978c0e8a55ada1783dfb706ecfdf66f7482a9f2514cd553167cc2abe039607eafb20cf88a5ab2cf3ecd3e1cf54e48eccb2579c9641578d681836a3b0409b3d63c99af94bc112fa2601f7b8f44e7485e81ae982783892f3d6302b9fe575213c8bd17655732b4431058d350080d97d00907e5820a1bf9ea92d49148cccf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13d5c108a8e23f8d0d1213aa2ae6da33e761c18c1be6f1a18318a73eae346b9a5d64282988a2168d8f256ef5043118ba5d5c560c9aca07d089c1a4c7a0e0c42681fdccb58f8f4e8a53df39fefaae6e427b6c5b125d8899f4d82fe5b21ae3109361d9a841101712f99be8424a76ef6771ade0f72ed7f3dd0b1b29c4d406122d93;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43641ca3cf06dd574d714e5ea05f4394eb20b0a4ff10cdf26a0630be015fb5898d7d7bd9470817296cecc14e73f6889df34a8f6598798313f2e5ac5bb3916fc35f62e85b90f4e0ef959ca4b507bcf8618e17a896ee5bfc974bbae1b15bd4c15fea9b02dc9603230feeba85764074d5341166b6e9f6568a982387e96e393fa029;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h304a8c3347e5002b75ec8cf50246e814d70bf1e4e829972775d7a7b5a8e5a604f5f0f2c19922911cbe353c07ace3012bea26132a6b5ab927e3a42953a04c2a0a5c607cf2e661e30abc950c4caf2fa6d0c755386eb1c1a4d96747a1e61d75224b711b7fde106bf806638c5ac5e76cd38fc751975fb06df9275b03f967568d194b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f29e8a6e49a462a6509066bf4fc483248f35cdf7a5e41be2627c6b9a5b37100eb6c3e684124d6123dc20c14c20a10219525d78635d6b6beb7aeec31a3852308a0c4196012ce8e9c822cd12f9e57769fc7cdf1de3def8d87ccc0e776917d3470be6af294baddce7681bf6e3ac5300cba798292de65e600e3a06a96016927c293;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6119d71a5fdacc7c774e4aabf9ce8d344a62ecc9d7f97d7a402d969dc43d1238aafe4ebf781f82d9377b5fbe18b3d8ca16795d14b7b3861740d294676b905e9d2cab22535a21c91445e2dbb3fa13abf764764c1cb9f8aa9b40961b9a7f7fe00b330ddcb4c74257456670686ca99999a9adf33a7d23783adb284fb77abb89c9f8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcee5b8d798f4e86e1b92fe0feaeb06fa141ccc9c490043b8cea4d52c30a539daddf2ed81612a896ffe5162bac92b95683995a25700fbb842a1f4f79a7af0c7bee5413954d1960775b23a744a6bf0b856d14c23117d4d20279c25d80aa31eebd1f5a1cc8bc7cc5152421271c1f5e83ffcba70a036966eea85129e4ba9dd288831;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbab771ffa523382886cd60073a2630a55152a187fc485a5ae5176f80066f2109e3ae852cc2cbf0d0152ec59250454dd9aad14ecdb9a3864a92f87a03b0d673977c0a5a334f7f832c5c015657d786f50d6eba1e2cb92882931d0f3f4b1f352d3f63e8081bf059c6662708ea5a335a48dd1f5956fefb38bad089b759dc3057ba3c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17b835838003bbc48ebf0e61fb3da2ac4425cc8859253a57f776b4a95a8b83edb2489673c77afabb679913e1dd1e89fd86f5a8dd2c4105cd7966d5db67ae125a35d3b97bb86ec5ecf186daefd541aafdbc8904e19bd1232e2eae60fe0b33627684abe5791195a89107232329d4c038ee799aa6895216ca9cee1830e9f742652c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d62cd7bf298a99d5ef76c74b6daa1cf81e03ce92b45f704c114438200d84e646c61bf212cf322ec1759c5b125325b78b40817d9de6d8c73806e603ba39070c301ce31c2ce85e41b43be47edfbd7ff292d8c3952e4fbe160d9365ea757a2b811a1e8b37022c0aacf845dddfb322c02a741ab8c1ca9e5f8a9aaf8893b010e409;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98eca47cbb6c6a988f793061c91b4049f523cc1f1b6c6ac7a6505e1a1b29b80ae5ea9c3f9703d1ec117fa5a4fe33a4148e4131a8f6b9284b6ba35f21749bdc179e29623b55fba0247962ee446faa0a797c0571095bf41d08842b0686256401b31378db36feabb32f30e60082662a99296b6f0010b3296d7dbf0188c2c5938955;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8acd60926800ae9e688a5630f4d57d049f257ff44a85750c1418018f268de0c27b5128c605029288b5989c3be151930cf8afae542b46cf1e706c2a10ee26e1b337930ddcc5ffe75300577a8323942618931e08f4e48fce54734bc6e16728242a3a45ed4fc13bf980796d519c845b43eeef15ff13931f733d27bc039de7495426;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa485d4d775efe0f7fa90e4056fe67a3797232199d26402e9e60288ee00507163f3eb1a2eee52bf1aaa1a108a8e3b0ee38546af2b71ad68108e931286b22d7335a56de7f08d2ff7db07043f84c175e9977433c759871d7df2cb614c15e36aae5cab39e8beac5e9672617cdf0a737a5a182a6902730efcaaeba3c118823b558bf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e81bae7aca08a6cb6c6f6257b80b0c0a2bb0a414c2e5f1da13034632378d619b3a740d2666142ba6426c14bf7f0943985b250a62ca6dd0eb98d3ea43549fe6415781021cf04c3cc31c04a1ae220c1badec39e815a82949b06db7024dd33a8506c36627c720b8cec9c44e10d09a7dbf900c0188c9319c6bdc0376178c33e0519;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b605bdaddc80f429afb52df4518f6b4a4971777ac16b8bce4493dc1e0e797f68472fdb70f19efee67799a13753a238d43001ac60b12fc3bb98d6c9d2fe260d05b24e3aad8506c89cb2c840a5dba17c9d4cb49b0c95fccde8d7428933fab77243a7c16b72753e8b671f9ae5e3ced22379c29977f27287001b47f4b2668a1c3d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ca8d2320a9b1a93a2aebf7582c5f85a347a99dcb58ecc7e4e09295543357fe551d5cb37ffdec3b0ddc571f5ee2e418fe1b86249401b490277b305dd8775cdd5f5d925e28808dbeb66630654e2e2bf099fb455b67a0234109b34c6bf0f5114207a135e765f62f0bdd6cf060525eafe6930abffde7010c7f7e7ca6888cae9550c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4fbe48cd617c1377c3e3ed9012c56a1f697e716625b4cd367b2339a74ea002665608e90721b4b1ba9f231a94579483b90240b7d4286a5cb8d27d16e15783f4210ad8327f7f1ab57346185c8de2791c5452067bf91c7b47b20e705dff9afa5677690684efea5b344144edbb5d5ff5d23b3c58cb7e9b4b7f492092aeafc27570e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4bf137fcd1f5cf3301cd70accb210a138db634ed33a2968866a1d69486c4acadc2c6e2dd16c3e8b62241d1c9d5397bd6981336b12e0962114b979afc4a1eb303ce2e24230a148218b6be215caa75d4ed468dba2a1e4f04f3f5dce33ec8344840d7aba077c1e6b51e10309382bd1dc7c881058d52ad671a1c97d7d73b32f537d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hebcbc204f1ec71b7f9c372a2798772b75104e4b9bf52b2e65b7390a3963db02032b50c27c4c2c194a6640c02a787cc34dbe4265baeffeef7a6927099509ef15f9b74518c359375527fb6f8d02aef022bc3e072e617d712ab93887e803b9146a9a3387922cbd98e95bcf86a912d93dd7098249d5a7bd0c0b4bb7cb0666af1a36f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf8a63a8e6eaa90487390a76464f3b40a897d23aaf21703bb07cd52391645e507d1f7267b9ad0e95a6b9423ae38c5edee718be3eca2ac8ff02ee1dcf476465c5ed39126de2d043a6cf73a4beb2adf3ec578618576b6050a74b481556ebd02baae8db957465f514bf45448a4d02a5cbc17b89e978972c6fe9662e7996d8cb425e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4aa8daa577a20546b0aaae14810435338c7b24f62564f6c47238c0aaa848b4861b3ebe19b9a4fa8f5455e9f1b5606b1e111c95f6dc07825345dee0530e3fcd67e5942e0164792ae576eaf301931a62884f7a062bba26f33a2889d4e30c5817bab633fd951be11a1ab62ff8e04afc1ad41f6d351268a37b6f7745145b3cdba81;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa03e44451f1cb258f99aadc3e089f50dcb11ced338215295ba5dad7d51e1667d99d057ce515ce10936259f01626fb27924cfbf4378c47228bcf46db5c1328946cf3fc2dad17ae550a14d25f65fda12f27f0d7ad989cd7f6898bc72ee74851110f810ed55da60f7f494b6bbe7da5861ca02f74183c1213981978a6a57c28925d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39df3caebe7004d3b62dfac542daf8c80b04fc09eab20dabd012d21fe374b2eb7061a8c123afb4fcedae9ca96853f4ccde474f12ed8ae4d577f9e74c7ec03d8064c1893aab382eb4a1cc318309eeb4b01abef13a1499140b687a71724e72e18ac4ae1f75518af7b00238d0c2e10b77432ddbc6df239d95d137e569c22f82234c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55f7182a463903553f4b250908ea9702c8f6403474eaa63382bdff1119907022e0720128142e95972df172a436c896e9a013b999cd3fa6931f3af385b2ba10e19722417c36cc98b602f1117e7880e5d4015ffc242033527b8e6bb60426d27f2142971269cb00da2541dc8990f7bf052e2ea02adb9298c91bb016bef562dc3a61;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52ff1095832e3c9a76104a9e2c35468cfc6430ff58512672193183735765adc92b724489659bd1a5ff5ce01ef2d9671479978b9ecc77173e5707dbdff86713df54d51ad4c3ae5fddb4f2c66e133b1b54f227e8438e136f16c6ea10ead895558faf68a65e7f5d23644960d14240eb4e8dc1c1daa259918fc15b5bc9b3e600f379;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he633715e8cf05ee4089681c59299b1149b868a5756feabfeceddd730c903b0217254057cf795ca2bee397ebcb31da21443d3932cef5dc7eec41be9ee0234389cca5d4a1c09d3ab560997ad6cc5233081e632cc0d7429108b1c3ca115382d191c90dcd3afe4b90792fff42818ded9c476949789d402db29ef82a554e3186c401d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hedcb3ec2b997ef108fa29dc31da63c7accb73f787aa294bd633824a6dae22a731de183517247eb111aeebd420363a033b6f12644a6340f3096650019394809c13dd073240283e7dc4bb648073048d8262785e5e873b9e96942d122eb228c64b97fb730dc32262cecf09c3bf2a7ef2d174bd4751b1c9aee0684a2053fdd1a670e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a9f022d2cdd93d9812dfc55fc9bac9bcb801932cb3241564ad43348578ffde329238c87bdabc75c27ed7c2ea54472e89a4c393e9579483c8bae77fdd6b7af043933a609daf80dbc7640b6191bd40526121fddf96372a5b6df7806a939ea1bc5617324c3d60290fe7b76372f75ec55b058b545e39bd5683d1a0a6b7ed3becef1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h683d48d34dd6a23358e24869942315593d1a9aaa334096ccb279321b0a0af9a903dd08ee0aa33122dca4f60dc9256c25f6ccaad17b2033f417453c22e2b6a8c2040c30ffa3a5be85dc1c3bd3f4051691c27dc297cd3bf08ceb3fa5c7f85013eab693f2367bf77b61c858115abda702509278c33bdd429cddc08e62addc91965b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b31b8fe50236ac8d8eef50d28a8b067197cb1e0ff5eaca4ba154154467fe2751b88ab04da79e03cb43a8fb7e773beea115dd2cfbff34cf28349b6c6fdfeb3c0e528690f6147b4c68f982b8486981f1bb550f4eabac53e34a90f0e5a9d3b73894db02494070b353ce0cbcc13ee124634858a883eef24342a961f621e54652f1b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a1628dff271d232ff1f89e310c67ba5bc7ed5f6bd54348fff733c04f383295a8181c8fcdde90ecf8c6fc7b140ea49a2026ea5afff943b066387b74ea505134aefea629bca8cab2b7e02eaf42ad18b3f98642120fa71419ae7637db9997bf359857d87a9efd5b446d4bb1da4abbf58ae5a3d7ca3175d105d9f05d3e6d5762ab1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h634de7be52992ed48175f51c82a7bce038c15ff876bd80069bd53ebe96b11874ba5e0fe07ee690cb8de6092a0fab381cae72beed6ef771abc912d9e6bd76ca8559504f696ced08fff11c8f9f7af12e84a5288f2b8f31240ed64bf4e015d28079918492f521e1b89b35a493dbf09a4e28f277368f40f9ddb53cb2788a0cbeb20a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3dcbd9e2cfd69df9196fba48620588a8d074345ca2d956093844dd04815654615eba4f091dbb4f73ed20b63c8eeccdcf59f380b56f8fb1e144e66a4bc86b753c1ad4f9c452fabc1811a2b48ffbcd873c8b6989f2f86cf3c384e199e6700ed5f9a4dacb06ae14fb081a017419be01bfe64b7c06ab41071ffaab41c75675ab6ea1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h60402256c515dc79a595e4ad06cb7dc17a5c104b89a7d4a17c3be8ca3c369a25d34f3550792cf1819d3246e9cce05801a792212d082a0b02bdc792dc4931162b40a6babb4e2deeb412ce48eb0d815ddac1c2ad3c974ee8d6e2275c60cf9b1ecfa2efa87cfbbafd048eadad150244118b553bbea332541fa6a7401d7432065425;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2c99dfe493824a24000585fad51af004a312f4d3a8cba769e595bc36b06eaec978b0a5979955599846540e5908a1dac70686c198dd9e4c7ecb2d2d0d065cd02ebd8007583ae8f0f1d3b01c2ac5bb590eabced8a1243f2fe7203d8689d309bda38646db381152c1e75858215d036772fd0194b6d5f4f15d7d92f07792561a40;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d9937340aa9978ebfaba6eb701a474bf3d97145c99e73d7f709dc27a5c31218741a01df3a8fe2b8d5e3a9fcd771b38349ffae49a82f1bdc9bdd80d4f9af04b5e6af3f2f034492ba466aef8e3d7f264995d912cf44c2c644d4529aa914100ae3c961c73a68bc8b4367a51764bef4b76071ffd41aa8e5b8197597edad3c9167f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h980b771cc8e24d627ab9ebcca3471464db8b80dc23923d8393d680e4fe104741cea259e77858beceaf378f2f5bb8f140ca82e500b071f117c291ed90705a521f3e77ad2ba5fa98831597204881ce2de6ccd2a3b724becbcf5146bf284bfb7c86d99715e1530f40b0e8c768ec2bfd5e84e4155bf67efc9bab169f152da057818f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde4694a5eb2937e3bce657b1c7b3980cda08cab989d5a2091655a2b09d0c20cdaef7ef78ba72f6a1327eb6ca017a8d377142965d9c0101580e2132e0d678aed467eb3594bc9261b18f2a52ce307c79ec7d8b3d43ced53925a27bbf16df0333b9b3586b4d3bd7eccfec0046bfa09d5346db8491604dac0819bf49fe757bd7cff6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ad06cc033b37fef02f90d3cdd42966da726a66add85174c5213cd90451241b90d16638e73f3a90477c313402e371207705097a4804431011c413d3fa260bbc6ffbd722f55b0e5fbcdb42762a5b105ef92067e5893a5410f9878a0dccde1beee4d44eb6184651e9fccf6d2a226a187d400b6ec6bec3ad4cbad4454c67d3def0a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d932d08fd24c84fd02f0010a212e9d47f08811725fa804b4fce814d460968c289453fb1ab2f4992ea18d90b8220f0507f5e6200fc38ee9d3cd92544de34f646263e8072bf436115006af3ba8693c0af70506ce7fcedcfd854738bd735fbd59d1d81cb00e0ff4d144e809aab544c587be105681ef2b17d71bd684dfedff005ea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h14b708a4026e0102e42c9a1cbddefe9737dbd74e1edd8f26ec54c5e1e4cd193984cd19cd6bf47b5b1cee01d93da1c4912225b672b89e8171d91483a39b900f009e123e73e233e12577f90de6b4a49a49eb77f53b7398d71bc671c480c7c87084a5a2094448704c213cd5cc99bdcc7aea8e4e345241b150450961b70f76d4fee3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5648f5dcc72e5b6fd3184861db36e7ad446cb5d171bcd6afb5e0e1be8f6c94f5870479ca964083f25e8e219101e7b501656cefa5551ce6e3f53e644759d6deecfa541d7a817d70ca6c8afdc8a9a04b890bb8eba82ce704408f087fc64e93a53af446d8380b09eee1efebac051a6581ae1e266169f127570fffd02ce0de63494;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47c8e063bf381253a61030e4040b8cb6f65ccd1cbdb476b4177ce7b74d5244d0fd481b8d7b1ecd663a72c015a262c5fa000da9bd39e7cd7d1ccc49c6f75850c4d8cf8ac661a58ebac16a1c63fe47a23757dbad0f23d5be823b2f876a6c9f2f8111b898760ba22e50593de8b760533fab5c10fb9c91f8d3bc60840647810963a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ccf23b726f95848065836d20cfe396a12b9a1924df33679ea27188b96e7b19992049b4210969697ef14ee1b34b3bf825b2f86da69a12eded2e3f4fbab76596de9bebfb203fe1127dce46c2fdc139b002e6690e84b894aefd5a460d5f91c9fe32f90cca9a8028843e4c083541a2093632b0a5aa3917e72df4cc24fa371c843bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4c4e46aa3eb22630c2b1f27539d90c2ef80971180e9fd22fefa9049a2eb06b718e6591993eb1572bc5c7e478ba65fa3d9507cd34f36900ca38a89132c150fdcaa28e12e43879508fb19e084e62bce99cb3df182132d5d6c09bf1aa423d7259ea1255d16f7639b5a7d01d0bfeac199c39a0c6e20e75ba8a9e8144745fb5c3c1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h56e4eac9084ea40d3b58e7aaf899cb2d4944575745677a21db06a8fb7fc8e15df06b6879c985cba98701aebedd14f6784ae418e3031295be1d6955e7fdd17ded5a18aeda241a1a80bd220daf8daf7fb56da96f3c8b70cc54296720578945b5352a52f72059c94dc741369f8216c01c3eff24120ae0462355fb512a6275572e2c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcaf835b0e3c716a8d43a04841bf8378b02a320973c148f9051893ce176504c510b3d4ce1c03168046b453086f1c7ec0c9071f05f5b690e2352a6b91c9a49e1dbf67859cd2da3097d0c96bfe5af4257134d262d08ba8bb83130e7edca552c4bf1293ea6d15ff098893dcdc52d1ee48c3707ca3bb9b9fed287f051a3d8cca4ffcb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5baf5adade20a6770a226e354a6234957d530ea38177c23c2d67f519d9ebaa2befb9aaf37afa85bfbcaa8d025bb6c6a049529620ce176a8376beb4825f15da9212caca4e2b15d71a53b7ec52e2d20551e8916b524ce70ad85338c0d76688ab9779e2c9d5720f4cb831b8678fa58f3c50e5d8eddac6d9cca77b1909a7d524c86;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea45f0ace6cba2213daf51116683d3a12717c04e6256224e0d7c962a57fabcb136997e05c674a2a27c784b545443795b259eb2432da6fdb795c8cf140ab17f1c20714e94296465e3fe0389106f4eba6e3b5877d0ca19f3a9c62144017c53f09a74581baf6ec9cf86b22685801a7f0c07c07dd2d9e2d6d9467289cfa1079202f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91095f77f51d39d6ef5f8fbdc4325cc547f086ea704cf1b427934e9c476f17540eb98a4dcf9b2c769ef4e80c26a3af37fa443df9ed2cf77c1f61c4dd566c0c3fa1238072848fe0934754f7e9e450694b77ae33beb9f671ffdb1a4bf1c08ecc863e57ac59a7de29f283d56dde86bb1895c82138090ad55c0c58c74687dbd132bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4df96bf6233be35896a7610a938e2c87874634319ff5dd873534b52290df40dbc0a270f2d4451774502d2d0578599b2673cb38d5b55ed5087c2ef337c6a7ee499a77c5a11afba557613a3bac34745fd202594151ecc213848ddadaccfac43dc303014cac74acf550aba9fbc72e2d614640a478a971fa28dee50425326fcf081e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa087cfdf52ca86fb470b70c8ad8a83bfacc266e42dbe2d48140680278961c8162c4f9374e57aaa5f2e0d1236972941a94fc81cce5b360d6765439fbd25d5a3da0578dfd20fc6c0eccedde1701e998d29f988765a5125a48e90f356733352d3d58317490eb0951d39bf785dd54f47f29050a8076247b43239f6d52d0e432bba8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc59407fdee01a9856448c4dcc4b647b6f367b365ec01201ce8f66b723b130c0c4dc1b90ce7c2b74525ec2240f1179869e8fcac97ec238e1da5df8fd31338e8ef49c5511d14a15cb13a4161bba6b34d5c732374d0a4a3fad75f8e51b8ae134556ce4ad375f77f71b9a5c85b96b74f4e411cf31d3f0d9f3031042983f17d6cacbc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4cccbff319b3a99e6ad259f00ea76c2f01cf5b80f4a225e946dffe91eeaf2580b803bd07b815f2d4a4a539e09070979dc175ebc0c23bbd7cdb4c8d88f01e82e70ae10863116d74d2e0ba6defc5ff4b7d8f1f15cb037114da956b1654278558e0b1b21d5ee520619e39e1e4eb49731a3a4741957d54225aeff6c3a097b04933c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c4d7c47d3dba7aec68761502af5a3813bdeffca9a3566d2bdca2a8964a76e871cbd806c9cbb268eb993f7b75cda02cba71b12286b57137597b00251946d8ec344488ce03189374a13cdf07cf84a05602c0db9454fbf0b3246c0949718dc9cd40c82471290d5da7f5b6f8b680c35ce66484fb720c167efe038b4e93f64a46108;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6463c618c902eb6aa0e18fd00ab379f8ade02ab4e576f8e42cacc26b399ea0ff8caa044afe2865d4d49cdb5417acc37b0a3fd7c43d5871ee7433c8282266df8565940657323c90cbf40ffb516ee5c245925de94d6c0fae96f28f8606abccac7d2dbe8e34e12661867ce30560e1a828b05600cc3edd4367bcb2d324f74001f61;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha23c14b0b8d6901dfd3e456d9d1c5706a198de6fd5d269b60c3fad1a946ee14c099b922b7f52ee7a117a3c98be781e2f2eaa41af4ed795a8edbf9fc676789698900281d0158e85fc5168c44ca220af5c4bebfc523fc5e15590893244932ca706ee89653b738034a611c200569e7c1ababa35be2941dfca2c7c84774c4022677f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd86a3b3a8b53ab9e06488e488d843675560c9f4fedee9597baf63ea318cbd5973b9c7c290f37d589c80d9610a3c141fc6f0cb098e7adb7e08d39780ef8052d2a36d2b510cdf3eafde604655992e58612e4c9e320aec558a777faaa1fd6cc5ccf81facde6e0ba9bef69498eabc688be74f41771ad4f40c083cbc9d5d7be5fdf46;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33828ecf45fad647acb0489c47059d48a37805ad156b4d1d4664bbf06533e0be69b929f2f1d572aac90894813d2a10dddcad73878701d332c4a0311eb167c76f57934bcc5b0ccc805a124706e8f588f36e97128fdcd614760a6c12467fe358e6fa0b06fbfc3c2c151336cfe3e0246283dbc436555ba4462d5b76c7a800581a59;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h63ef057165da9d1e04c71e160b4255c566756caf00842e423595ddd6a2c7908b0b8386191d56ba2a93deef1548a85d0b5cb946c7826979466ab82a268eef49db4b96e333a90030fbb280265efda1239ecf13ffc3c3ecec992f9267cadcfc5d058a29e848ba8c2c14d035e77fa99521d8cb8506075eb87715c9a862d330ce4079;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5256162561a42e1f1fd2b426845d096755609bc4fa5de4b95eefbf8adf3f780176189392b393b0f9c00e8edf23bc5925bd1d12ed29adafdeb054674f957744e72b791e6ae358f5dc7a30e1e39d06817d3c5ba6b78ed8e9101b3689461531cd064d9c49ae79c514c569e907acea26429e50607ed955c1c279835546033414b01f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ab6d9c89e30f8b295a5e011e19423653a7a5a9000a9026fccbc723872f43fd0d01776e9aa2e44c57b4aaad3798700d25de26d206818ac139252f0625ab494383e548755989828b26aad46e340181fcd41384c31311e3e4f8bfffd9398e5d5cf02c331bcf2e78e559f97e12543cddb256f6fc377dd1170494da72a5a0d4d04e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f860c0ea4b8816928ee55c6dc8143ae3904a0e258d5392463a0a22464fa98689a64a2925fe0f0f27a017020164a1a7d8fecda0837dd9fe9dbac652dd007b7e9cd14ca221ca2e48d4af7de11a472240c8480415b07197630ee654bc7138ca594c41d6706ea8ab80aa27949fe86a1561b7c3c81d4417b0b029393061f96e7b3b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13d9cf76f6e965b217ba3054b2cd33a382ffdc059bf9aed4cb77177d448dd70a0d09d941cb3dfb224614a2d8f52e49cd27f4673e684e650acc9b7f8d74008262dd3c49551dc6572af80530e352eb922cbe5654f486926abf7af3fa361182e80846d047d60e603a8bcdfa7ea1ef7ad88e8d2e6c0270f37e3afb2826d048777b50;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd17e03215853260f00f43a3350c49bf38728b4d04e6b7bfe8eebe75f7e099118a2ed0a744a059eee9e15f761836933276fbb7284be8c4a992a6cfec38d84ea4eb26d062df144a792500654735ec9bb650893e2f03e6c6e89d44d68f316a14532b699b18fdafb40ca9cd9b5849836bad16b748547d35354b7cedf654f9d85f05;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62f96e92f60948afd3c784553b555a5340072722a82ed6b13c10b208643767e8eebb876da4c0bc2e7b5aecf425efa1bba45b98eaa0c6745aebe68ae39bdb27539102668fee18d0ad7addd90fdb64a6f6875858d8886fd7ca6cd079eb19f5d46cb9a8bd01722d4b18cb24ebf109dee002d2b4f32e9d3576acb9471a7040f0f600;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffd470f03b215d8412483eed9856da838226f09e92548f45541e39444ba57f1497563624951f649dfe724691db62e8391de0a4ec8b4c2f8427464a18a145751008076981ef307a28551b749ae82122c7113d5a15dfa388ffe84ec3c416d9663ae9c62799664d96d7c82442db235a24352569044588e9b0e7aa3a2945befec1ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51c92c373dc008922e9c5b2c54e2eb390939d030b6a91430a8f4e2b13dca76975fb5e010a704b186c060de2862741ad9326b672eb973f278f068438b7fbdd1bd88328b2ffda5e1660d9c80c88c8cca144c245b02dffca5c6f386e891dd56e1ba23d619e8ab99d26f3f95ac4b455fe189ad766326dcf65d083f5d73ed7b29ba6c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h989ae39b2f598e623d0309d474198cf48cff714ab662b20bc0e52f3832f4a4abc62034810ebed5932193a1ed12937597e61adf004812373ed4663f37f726c28bd2c53592ccd7a592a278413f9c80c265d9956ce305c9fc27aa00ed888a6738b8360fd2a887ffc2719f4a0e8055be20dbb4ce0aa06f7e9669d15bf1fc177a995d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9984f229b42bf78a4b1b15287a15e31b3f8012d5ec9aebdfa1d94593110774e5451c6b134bd8e302385e64d163e689417944a37ee1f679eae4c367596bce5a7026e42dbf3fea29e73386faae487445f6f479a61a890a696e160fbe3a1652754e0a3e7d03fcc9a88f74ca53c9e360f58781adc2c037548c62c6c5021c5986348d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h25c2f06b91e73bf4eba25541e3d3839df6795e10ca87e329be7efeea3ef8ce1ce508122e1a149b756e437130777206756e75f283456cbf13d9f22ce360c5b9fdd1b19eebcbab07dde77680d53e5007493c40ed672b8fd2839843549784c5128e5459d82b5f18d50fdc5e4fad673aeee1f7b15a477a61ea66f6578d58567396f3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e75c6f2b714594dba665056ffe8c068dadece29fd8342ba8a954e6418d4b28633235c4d9203c2fbe31c5d111093749db31199ea12feae9a151531f029909922c2e19cef0676e21cc7ebc79ff6c6ab249d83b6d9c6a8dbe6db331ab8fa65cba0e597f6153bfc474d636b7891e36e4fdaaf5f4671c04fc98676c1549d0f34776c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0cf6be76aa44381cf19084af743b4b0d6ad66190b257cf1fc613dc143828dbaffd386d858f67549198e2e7689a46d5ddc4eecc0d3af7ed6c3337925aca1aee22ea9a519500fc6c0cc6f7f440b8415a0cbfed1b380db3fc9d47e6c865eeecb38f9866e4fe7963d45964645b485843a21aad151831d498d659fc7552cca7272a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff6d55c8d1795555e3eb63b92e6752f23bb1a9b8ae1391e5ed30005168229d8190b71b29e9b5a8d0e9eee5285cbc04aaab5749c18fa77c49d365c32761f2b5da745297fd566e62d7c62c4c6b799497f021e8d3c3d5e7aefa575d79f6bfbfb93da07bba072b0e0fcd93798bfc35b007c481be0ab0427989a83f9b6408a0dcd579;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heda727e1a9a8ea7f02c26fef09a0ad8e7b1b3f0c09b0823634c22cca44eff259622ff43255134663279be4014faf8e4a811beedc04bf0dc9c64b2265bae112fcabcba48ed6fa3a9a17b7f81824d9e0983c18ab47c7a57d32ce753d372a85ec1564e096d0aaa1733d48d2b4e2bcfc68d7376b473dbda0d823869fb46877fa54ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54d065c7f2ce0b9d47bafa1c3fe5d98cd7031f0376c0d1c582595a040244901a27b477722cf980cbb702b6f6ae672316fbbfa16de1397d81743538b6d549aa9fb7d73b92147ff398c2225494988e091e3a39bce761788663397009625bcdce394bac0707f576bf339e241fc768d245e60e3d8cc9e34dd2947287956ac277ca7d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb42136ddd82426ae48bc30dcb6537ef87c3b6f769e12e0a1454bd1b346ceda0fd58dbf97d88e0ba818087ac2971e64f0a41e875e4fd122e4d5da91bf800e9c2480bdd423b63a2c9ed76338c30dd2ce95f49ae16e5f0b915eab0a5fce19a549c8f20c00d300c1dc4899e194e6955d9a2203c6260eaee3594d0e767192574c3929;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h996bd71aab1161db07251cd9ff482af24429a2989a74769522033040eaffe0528c90cdda7ccc8f239b26a794577e33e38d83afe4946bd650fbd0480057af86bab4bde86b1554bc82f94fad0d6a5a5be07fa2b89c6cc4cb7dee4570d8ccda9cdd181d2badd9dd31021f1e0034d203c39bb109247d4f85e3cc8f06fc2936c2d7f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e9bb101bfaa583a93a1f52d113a54429697ea455e4d3b994283aeffb7fda8d917fcb661cb2b3cfdd62c543e72c76c60340685ba58d59dd92aa9f229e0b2e1ca98354692f1bab7fa0a28d8253aac4e0d4066dbe1c11b2191cd9952e04840af4a52efe066e845c805634cb84bfd98fc27d680b1551b05438f3f494ffe60013658;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he63ad2320b48dc81911a5b76e5241913d3699a10bfc5f03147551800ddfda2433bdf6dc8a71461819f136d6e185c641830b3b8be99bb5af278a7527316d4a5e9854d8c04ce7d3b2acfb84784cb3863dd728004a35ad5cb56647d6f071772fb522023411f09a104f575df19ce7b95c231ac0640558699f9d75121803bfda76e16;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha442f0875e6d8bf06989b3fd7ead66c6708320b84d642ed9c56c8f4e2d4733dff850fc6b98bd61d8c24756ad5a17cdb68a40e884382d7edf04cae2395e67b036413d38fa01d8a80c6cf6b7f91e637090b8564158a53ab3ee5c7687efedc2a11845fceb3c8e3dbb7ddcec2f06d325a551e02cb9e08ab1ad57fc7ce09241b1e65e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf447cb1222940a0cd191b4e88f0920ba063fc531773460a2327689305d91e45f653a809df540490c26d64f11db85ac8597ac8c4ab1fc84dcf4bcd7e05cfc1dc50b724ddabaae0843b4322c64281249ed6a7bf5ab01df1dd40292c97da07ef80ea729ff1fc21b074096e1edaa03effa3c5c206afb12b989d8e3c38894ecafc644;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb56423ed065444c18108763669c598d57bbf0a9a282552a4d051c4737edb53a63beb4659b24e8cb9bd778e0e3a94900b4cea4fc469702ec14b9b47caa45bde2a91ba677a818c79a7e454a084f0b11d61fe42871a2454ee27e4b926640c658ef04ebcb1ef02dbff17b5bc471b4a52d69784688d995654ad45e14f15535eb6d2a1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f3c0d19b80a151ddd1ea6391bfcc4dd043cdb0435512e50df7bc4fa26fe94605dae052101c3df8cf5d817c270c36c016160e6b3e5350ff7d14be25dac1af61a2fd7489767f61f6468086c165145e5e3702cbb1f41a1178fb96ce385107eec4b56585959cb3ab61f7fbd8c81c255d108fe9ea2d59deb60747e3c52cbbaf8016a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5adf64e7a723713d3f15691280735ecad52e6d0c18f294964ca80480fc82122bf6ddcc25388827e0cdebdaaa60819763212cbecd51977523ea5f0649b447e4ac97e74f952f501c8485ebcac7968fa07b40308534a450416e27e17e6338a205df4cd04b28d7ec4fbcdc4d8456c6a6eaab85dc1d1f08eb093f345da3eee5b9985d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h242b300dbfc6c1bee718d571245aac50b77c133affb09b7a09bc2cce6a8081862038b8814a7d43c8ba5daad0bda4257c21d37290a78f03bab2441700ef5e1b767c767b5c650168fc75274e9f1557d2fe55f416f543d201ad2468c6a1de663138b3576380754136aa02a60de94a97c3c3295b192832233f32254fed8e4c692aaa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8308e44e4321e1c9d7117d9d7d605467e7bed49b6f369a3380fdf7e3e988da61f40f231d0d3da1c99383e905ff055326b4e9b485238214bba4165cb01058e36f949bd4033e00305883b75f1204e7ea8fe92d1b544deff8222d7731e478fdafa2629b26c1bcbf83856264380608cf2cdba1ef6a4dd88f8944842823887153e1ec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea20c442d569ccaa18e5418e1518451127fdc3043941081cdd5aca2565074f1047b77f585a983697f1ed9597b467c55dc66c1711c08d9180b5ee2f1ed2bbcd7e4b4d68beec7a95d48666362344e8a5a820002de78191b327662ae2dcf94f2dedcfe1809eb782e9e25165279332a84d278f98efdc3f24cceac28e390cf2b5773;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f135984847e4668e5394fd43fc7797dda82a80d6c5f407170e6514f744b7843e3bfffc8bcc24aa77dba8a17d129bf24aded685c238d986263557cdf4951842e0cd6ee48dc4d623b371a8e5010da44adb9784e89991a293ea170d8f223c5132341ac230d1354a66d8c3a64316ac4ab33bd03dbed52bd911621eef89b0b24c72b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67c42da9e251a8fd32049dd9ad82fbab73bc689df46ac7b4b6387cbc4174a022c73cc16706c704a4a2ca103003d3fcf12a80107b5b6660a7aa8b2520ae14bd47af0b1f61038dad600ee5020fabad2a92e97dd036e7f19b503e0d34822503dc92f31682b59a4f3f296568a7f46cdbb4e64e6ac31d0520942aeac6b1dfc7508ade;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had67d8df538a9e8c91f7be0183b85805130c2a70fb8ad5ee63c78af7308ab7b7c7464f40f2e703bf948780b657c9454e160dbaefbb1223c93cb52c3caab5fa26189a5edf020aa4b34f8fd130bc1ab0bd6c35725c835b0f055d5df7d7662adb1119866ebc2fad89b53657bb19f257fd414edf7f12b8ea930b4cc8264b384e5d7e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8748c5ebf7f8c6643b173b141a480a0c303a3cd3fc284be4c0d16521395e821716bda4ba8fd411e66802de4e3e80cadc05938da4283ff183be76d6406fe4688d1081e310da61757ed0dd266eb2c41963fa11ef4a68434b66ccffd137f7ff36ce72ded38a1db2cb1e165ace270e200f04322279ba32c10e09fb1c47cbb4e438f6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5984cd71f511a25142e42cc422bd14504ce568724aad5660d32d0617779aae9cfe751b7c1a48f67db6f8cfcb938c293c56fa8e669be1bd54ae93d58acac43886aff208d10221c82acad847f9b234f5a94cf0b212cec72e243b653f640eec6dedfa4fcdeb581d7c2f0497857289866c879daf8ca5c81c60468dc490590dd5cb72;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89d787708beb0a4659291299880767ba5207fb1861338131354aa805010a0d35ccf95dda7abba377331d832aea4fcaf8f4f800f683eddf89e6000b5098addb5563cbcbf00bda2819ad19952a75836716cf69617a70fd4f81bb7c77dd10147dc80970a7a6c1fc54c2ef4de537f290a53e6a975aff31242ad9e966647eb9ff6d0c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2bb608ef4105f5e20b3fb465c063118da0876d7d65a19a190fae9ad500be05e20f5fc3de70bf6bdd4b05be233df9bf8b490b1bc6429a6ed214a3fa86e36a17ad0631adbab3b3656957af615fdd57f3618964e67226f6781ee6b470570a8986e6d135517bf6e6189a4d5dd14d3a8d306f1ff9bacf7dffa356c111e5e1ff4663;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d9ed5f962efb95db395b8c01660455235213fea558702f27860a0ae9bbdea2bee77d579796215428989ec083ad0ea35ab21b28748ca2ec85454176b6998e0d41965a13eb3d0b04a82230432ee31b1b68c99988328412a582f13a6d911a253b7575651f6982a146a876c2795ecf823696a8abb7e74d423120043ec3ebe974b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7d7726a6bf10ca9696934718e8aaee930e545b84fdebe7ca44780f53b93a2ef543db738227f14de7f6c7d5b7fbc45f06f522513d403609c1f1cc6c8fbf0efc6709c64d590132e962710c7330273866ad2b52c21d989ab3cc0be8c39df3101946b4307902e539d89fa84a6750506435c2f62009e9bbfe23e8d0bdbe9d5801a2d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h96a4b21325e7a9803c0f0a1a78e811c1f782e49d016d6005e88b187499dd156ccdd78d2a5aba0a83358fcd6d3deafaa5e38b8a4c50614d9ceccf07cd28ed2d7164350c099fadd1ad4cd193809facb725dda8d34eb40f8c7dca774e34241d9e88b8195fd091e660b222c39be2af17150c2054f76a4a8743f9f718674aae10a49;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h979be6e3701ba70369c05985915530af3b339cd39adf23efda385931d06a1a1df9b6c0d0cf9b73ad292b938aa49a841811bd207d21ad2852e9453d3163af26e1ceae885256691491f78cf11e358128451d87534450cfd58e2ed555834a7c31d86e8c9cb62c85dabfedd2e076fc23e761e5c51b28baa95ae573fd414cfd633f98;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7bb96272c2bfa26d19206cac340527e0defb4230dc6ea780b3df5ceff5b7ab1841ca1ca4c678162958a25575eba54682934dfb39b5cbd64cb3917a1d5de2bef416a83ae84debedf62da34f47b23425cfdade6927a7cd4a47b93e42988259c5272fd3e259ed5b54114b4956dad9c7fef2387317634729e51b25f43f0bbce526fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h180e81e8438be3b962e4e6d972f16cbcd52fba132bff161a489ce87afebe4c4d2ce863d7481b5cf4895014c0a0a0ab7b7514d20e0754caf8e94913f7110615e9881a6b117707848714791ef8e835a7b96730747c13dfb86d5daaa3b06f882dc570998e5a5a9ee71978e1964452650504dca36892e6499eb95997aece4b289646;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf72c51fbf9c150487c714ee7e19c0e29ff573e1654d4cf64c54ed1d0f946459c3b554a7acc3c483ae0225e263d9ef54c8cc1e184b8c10fb8969434829dc942d33001c4a7ed9ff23df1b8d4cf118064a984e0e652874af333156a76c17a6df6043a6b5a3879e2a35496e6bde22ccf01fa8f14e112c3eb0917823791c1d22551d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h882aec8598073a74f573365496d1e777f53c543a085e33b94e4e6ef550139e8b46acae8a0f0d56f498073659c54b7ca192df3e51e62cbd11fb7be190d2bafb712ff65f2287a70a38392156d43363ac38284ab2b35af4f7366367d0f9194202b4adb85ba3ebecbad271309689681bd3ca0d13c33868e857944710d5c21adf863;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa6ff7487f84f5e47ca973bf7ac6be73ca85104b4e815e16aec798f06dda596354efc03dd681d1a7e9ff10152737d39ea6d782c9db5dc2badf9b6111ba7323b2fb9937e7e366a1d4e5ae3e27f1e05eda580d6e47a95a89beb1f6d3e1d904e41992f28812454475de69451c00eeeea7983af95e6d2cbfb73a91a0badb1d20773b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e1809562b13ef280fded74c7c0274c998ab2df7b057d32f50e1d5782aeead591d80036c56844bfd0260d7eaf0a85bb4c2f2b34501cd362f703a7f64c8f76a90b5c6d80284855a9fa003796f448b762681cb9656b04f07840b1d7457170f2264091bdb94f35150c3d72ab3a3b8e0c038318fd5ea1b216bd30bccfacc484ce37d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbcb806fbbfda6012934502a580f6d532d8dc4436178ae34014805a2ed9c96488ac096826c88b7062c1538784d1785c1ca5655518df782776539142169893088515b4fa0fb6a03d4834bacd1dac2d9b8abd33a2b7162587deeb300240b3de4cc432dbf1b63a8e2c6f2495dff8ed45981330a6d8f2bbf6b2dcd73f2976dd08b359;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he51d4bcd1a63ed082e8ef269acee36dab0bd92473bf81af84fd2d56cc917db5bcaa64f583e4baec98acb63b1d2f4e98dbf5d8f0acf6477323b5eb319fbf03fd7450feffd72c816d8c444dc717c5eb92e926d99c2864c030e1c41e44704191936bb12b9481de99932ad418fbe5f2d6a52c2f7b9ca8d6e2dc33116f2c7679e36d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f715a97749c73bebd2075a8e47c5edc7ff76d08fd1350f7c693d9c2813e9ae92e1ffec152a66e1192822e0dc4bc984ccb2d691ec246c74220581134a6158c88481cf4605057a58dc7869de3b5fa88c07ea8e3b76b0a9df21b87bad307109fc546571957da04601565d93a684c27a79ba7d0436ccfd335bfe0cde6f51604f0a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h77b57f49a75d6d56485be29bb60e7a4b4c6a74721e0bca93acc6793560787e49e91697e07d30d63ee3085cfaac5c13eeebb319535c8b6213c9a79c7f50e4dd676b696868fef0c73201fbf4fa791f9495782023ee9d35116b91c6311251678c9a6bfb7e27426be66f83d2c85df13498d497e6896e45516bfe6e2f26371a30ac4d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdeade0403397a888f2c3e1da050dc2a43344574f660d2a1c1f5820b36368d6d11f9c5b249b82a0a5ff0b77026ab74c517aad1e6aa03d90628f9cdd9f559c5aa8da35b3635f571a1b23344a216411cfbbaab221baa5c2bea2b4e14859ad60281cbd4bff75967fb95235cfda8410c162e3d0fc186d9659cb33ef9b2abb1da86a21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hecd519ed89ee350b2abfeecd52fb289dac548ff4ee3c6eac16816fbcfa695763fe0f1c89d8bf55860d62f34d70bc16447654a2036584ef40ee50210dfdb7ba881884b03c79d0ad59b4399e92a66969014c9ec7a499ee12297f19bc79ca63a79f0e34d3d721e0cee4971c19673ec8d73d60b18eabec983acca6095fcc7689af5f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he97dd41301243257d9f74c0786014affadd7b23833b3b1847cc5d5c9b464d03bbfb3c2ddfd20943b46dc600c36275d0620846ed901979da6a1f8baf58fca016745fbc8c88f191f34de71bf4a893bcbae7a143bc2fabb96e78c285818013710caab81a93682079492de1e6f464fafe54eee63f0e3df7dfab402244c6987006ed7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86493766ab0d3752d0d367c211561c2d55c36557bca6dff472350a53d0ec9b5e6bc8a58a7e9443369a9a42cb19003d3e6a01177ce16db30fc5d90e53fa1e2f4437970124663e0812c4c4184fae320e746256ef530736a0bb476537faf272c47a4ddde9fe10a04e5e1e9ee45cbf0fe3a4735627cc67cabbb1aa7e242f6dcd1a1b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc59c83295b3bfea03e674560e63b308705b239d687613ea94910ee5a358ac422df906912fad6810b18b084812c70a9b16ad038a9059bd7f914cb7765ef9a38cfa8c8e6a9d5657df01b184ca45ddf7761fbf183c86ef97314ac6dc0ae69e1ece3f925db2302683331ff37f2e8c909c08932965e53122d8fd09dd55d26c90cc1b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79d936969b4e5e74f683e4d6ae0f723f40e3afc890f0377cda59138a7fae96ae94ede4d4ff5e44fcb2b68a765966d9952b11d7a09c25b06592382c3100f2a3fe2ef69b23bb0eff5169b199b48913667aee62ec14c2537b4ab0ac16f9ff00052259451fd8b386a878845544138e3646e82dde1077a27f8947bc44c9bc3c1fd583;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb79edbae25774a49b37b29a914782870b73945452616aad5f20d83db880733a8a27e157cee4d7aa223e7a2dfe249306af16d8014d1883b011eedd1ddbcc55953526dcb370013f5d84a2b42373ce0788a612dec4073b06bc678e8d701a7a24ef565f522daef484c4fdfeda2fc02550600653fa500c399ccce06df6faa3d1c00c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53dc18133a11428e565e0b2d62143c244359e70286566e583c754a026ad636c0a82c68382e9dd183795b08a71c876862f9ef1c1c433a9f18e0474b1b5ce4527e72df06cf5d8b162501513c992bbc717f33ca0e9f1680d73edb83b70bbea693c034a31dd5b3d26884a925fd073d9e4922e8054ae49bec6c7731a8dda8bc880c1b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6fecd09abe24146ca6e12c492cdb873f09878fed5caaed7c36243e4ee23702a96f563b5c2e398fd671995c3db4a44cd0c12220a27bb19c53fcaac4bb6862e82146f323dacd582223613e19fcc5a0091890161f9c3ed7eef17627f7d6f1cc098989fd9f7227f799c3f06d9ad6a8c0bb91822355acb47befc9d5e9662cc10138a2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e2d38800fd5f55e173958cd8088b3203e2d3ab078bf1ea81b3838b0883bebc221528691e6ea7fa44c6456a52989ff367992da6de99bb986d1488a705f47692555a934c4ddd0f9162b30283634483964de675f9f0299f12a3727a7db27f36fd4279094998641ad4d54d92ca5a0d34579a2e741c5b6ae445f3b3f8ad565753f4b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a653b00e6c1c7796266d8db45135a2cf17b781d79e86a8e54dbb2b03793cd81df7ef0d604676865fe15d45c3536c0d1088352e8c2be0d9de20266677b21fcd4939232cd862a40d3a8efd5daf426c4d3b6ed554e2403a4536f18cff3b21937d4b515bcb207099ac077a22499ed9dadcabe49955aa319e8eae41561991c4aa8f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3be1e5e207b0b2b992318c5dbe9dac0b89d209210bf8cc112f8fb49b9355315a364b1b71c081ee771b0a6ef83992bb706e7384bc9f197cfdc9c230f8c8c6fed8ff8d186ec68543445fc540d7f324b79e27ecccf3387d1e9152c0a4d5c3de45cb495b6a5b7fbaa58fc0805e99fe9206de27120de65e73c17f8792eb488911c7f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb98dae61e5085bc1f400c88f344bcc5aaae44f6c5f6b761fedcd530cfb3cf6529373a2f64a65c784033d0746bfa2d3e8f046bbd5b61b1de0459bbe57ce232883107deff034bd68ef8476f9f00ad5c6e72710498b677069926a78bb09687a5888f9faeca5f2c60ee30ec638a4d46a7a143d392c63409fd1694a95a0fcb52d28e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h981f4a93210ade655bf96b675f575de878fefbb0f09fc340790775558645e93553cdfff30d6cdf9b8a89c372ba6be15cdd2734dd505a3f8e73b5bac7a3fd945252c7fd58b7056652511f0ccfcf6df028c6589633975f4a3e8106725e1c14d510758d5673741bb7fce368358028999f17a80994531adab7895efb1f4275a03c3c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1cd0fb7e1523bbb25a2d402f8d116c3ec6f03a6815605bce3fdc833bfc5caca754030f13f0106ad61b4306cd7abdd543a4ec1df9437cf2e23a7fdb4e1689ca191118abbbf3be6c42b52496d4b170938e6c2e7d649fa02e17f87a2278bc4a4b6059640b6a555b8d2bac625777ecb82bc4d62bb263edc5b3fb902cca2919c315f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52894508d6741a25882ea22bb4a47358b11ce48b97316e1702f4a34d38c2a1fb733ee47ed777e29dde93596f02529c7606487778f32ae9711d9c93837222c2827d3e8b507a608ee186a5e0e431e503951e9f4785b484d505b793237d1062f90e71b4ad1d4826175312ca12f0040c9fc4e917c68405fe45a0ffb4c27549adadf4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5df79b83ff60befacd6bdb1c43587e4592696a951057f6c52eee035f0c80405c9fbe1022a6e9948c10059249fe570935ab1a674156bd2a41088c15a496eee3f25b897471ee10dfba241078f291b5a69a8105482e2d5a97e7c690c7943b6e757fa4a03b474b5a2432bedec1eff99e2cc459c27c6923d6b3d16992a16954ebc690;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22a9d47df688c076fee2a1e8c7ea255508e1cdd94dfc9dcdd07d456f1bfc6f1b567ad3687f89b27026c99a52af2138d29f2c019179a889335724fdc63fb8a47331330e51b587ec6abe229487604d39095fc8954373d1f87afca39e5671fd325b10f90e02a0f69b9e1d0c073340b089f58420c91d9f5dad88c23baed40485ceb2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4c788fa24f04cdfe061f263f5715d33d9766cb5858ed09a1e00bcd429320a074d9480996c03ddb0b9394238d76810dfcff5f2a90c5790eaf2c1d3f35e729546976133b0786fd255286b285c99b312309e63d496b3fe7f78aa53a480f251641bae50b557cca81b5a454484a39f12609130e27673dc211b0e3b5a470d9d605937;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7da6124de8dbf0f15d4e248618417703cbed85c3d5d4e815f431ba6a4f35bbf4019590be32eec775ecef306519b231898ef2dae7752e073fe58eaad43b82fbd82baea8123d925465fff5a83ceb6609bd658337b2c47a98c597046aa8a905dc8fc0b5f2ddafde9327106f50ad5b8687b9f55ad0bf49288b56a361ebddb8fbfd33;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h839ecab2eecff471851eb8b1cbbfc4ef5012a66706b2c17c9f8f254332a9e95f88f9cef209942d2e2b02b53f7ac25afa8f95468398cc7b92c87cb02949cadeb6cceafcf9586baf89a98a157f7b30712d17818fc1ceace392e7f8dc08b733441a2d3aa65ce3069d423bc71e1003f39331baa081e8b0f96bbba911bcd721aaf212;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h304e8320bfdce3b110a23505f5a42f918c4de60e84395d50237bf074ce95ec49f1b60a29b6f3a2cefecbca2204a99886c4c3138247fb820145fdc31eb97ee4c4038d5435da691f873c3c5a542bce0977cd031c3c082f5fd25f6e94c9c52a418c98da432717316a1aad2ef3f1a4d9020223c50cdffc1e247494dcd42868118239;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3f987822477e0cb298d6838c5eb8df2601d3b95db94217a3c08d97420934abeba05ca37087b121691624b05b068f89d7ee3c5c5d8fd6eea2ecddbc9eb21be7d02134b95ad03d74394a1fc9cfa5598c9ca1e25f7d3ef1065f5073ab23af1e163b24a8fb7d751de17aa7012edb0865b74a52b0e04c8c2a8928ab61537b4a1bde1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82328bdd5e1edcf0e610a9dc466db9802abb621a4b1bf3e1f56a59906d0b419b9d7eea7cd8bb8a610f91ee84443afc32778e092ca5dbe3245fb8390e10e79e507e96aa2964a8dc1b7d8f6e4d5ec6d89f149f6324275293fc0bb05b17e97495b915a7c629e01c33d48d82220a144f38332533adf8290e1e9614007795b5dbe939;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa55779c56c9e5d7d8111b917428c41197e1628c6a9013afd43becd95357fb61354dd7bd72dbd97920a73b40f80fc92f864fc9951abf5b99adb0605db6e15c08a1d867752a1ff1eb8e2ee2825fe23eed734fe0be3b2c0158a700c064386db488fc268a81d803bbe9a90d2c9090b3f9b6c1eac72639d131485565418f404cf0c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4266f23676146ee5cf062eb88d3655cae581acf32e04a16af44453e381a3b796b9bf94979c72d52ecb030b90745a6e79c4d221280612a01603e09a025cdae36ccbb89b00a8c1b008c58a144cfccc2abee3c36e35ecf1c1768c2966e770134b290415e2ec576a889f389f91b55a25730ea28c60e489c2495678617e97f15eb33;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdbe5c990716c5dc0366501501d9126205037c245005df0702a3d7ad6c87ca27589ed0eca15bf6bf51e995e92500fc69c540346e7e4ed4f03e6120cf0e4ac8a9cab2d9d9622cf98102cc0b0d5066385e3989cf2e3d141a422456bb4c02f089134bf2f92b6dba6b52e27d07da8395177ce0d6af9777d80dd6b7c7dc86c5661bb75;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4cdfe30374b6959a667610dc34917426f43eaa80ce9762d683c549de0849de30e8ad733b78f04b4f557b3ccca8b480593445fcbfd39d98fb66a294094bdeff04b64b3a5b24c39e654ff9c58b5c0d1c303fbcb4fc78a342c54e3d15f3612e4909ab37e3b32a2f988293c06010e22a2cbaf7e0c8afad1c5bc23a27147c8982153;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f136fa613759915b18958c0598c54c4b83f2edaa2d150b2903728e7908986a175a147b0914c87c43360744e49b13127e6fcdd9e99272b7d5736b3f7f43bb0ffcd5c0e63307bf876c63294b3d83959e1d92f26ef1fd8f1f1ad39f58afa2ecfa387d73d686b920e1cbcc085182926b072380caba64ab83755cda6276d591a3242;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdfe5384650164da2b29f1901003792a5344d2f95efa38611548f569dcef6a4608e1d4027d112640c5e7bab7871bbe921501e71bca2cd0e638b66fb207f7b3f69b41deb6c27bd36db5f6e25d282f721e70f2ef09e32bd7c55473f9bbcc654ce4f7e5a0d28d2de4d695fd2fab9b6723d89e12669d3475a561d8846549b23c506a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe0c5d4a75f70d29fe4839f7b34ad3179f81bd351977280ae47a557325ea3930438d96644b90e5c2f4cb65e696957c4b257abd196bbe4d9f1d25612b130cd4ec2da92225d63c0a3d328feaf54b2dd83bfddb5e830b8ee99bc56805b681d3e8eb32666a10c90cee11243e36d872ae6da1bc11d628f7a3569630f1fffa4fc3016f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdad8d94e4f5501799fddda1d7a6b1a3bb14661b0df94d2d686c07e6678d3fa0d0f2bfba33ff596b1795d8dc6acb0c7c845db98f34cf0a6e46c2fbe75c26141ea9fcc506ea2097576e0dba1c3726643f4e28a56ed261c814c4d9f936c4d9f8edba06c6fbcfb1dbb79959373c2575b35ba013a2080b21c860e55627bf11b37da0b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1920ab50b932aea8c1ed4e4c5d05d29c4d4acc542fe4f6afcdb847293fb461b841e60dc592561436e058bc216c8497c86e8f67287619c3e01b2aa3b39717bbeed15eb57a5a5a667f5161228439f655e049a9bf8ee49cd991ba8392faea96a85182cb09f36cf7f969ded5f831120f1fb47aa31a784ca92b5e26b9f9bb519cfbd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f92dff7ead89f6935dc1d015fbbc4644db456e7c29db5144ba53a671d53607766c5803ec12a0456bd622157d625fb6fa563a8987dea530abd052c2e6f8cd67f85dadef04634ed1029d8833cdb659b153619de3d4a9c3d5ec22464a190a965d2363f5ba358d3a527fc0844b216180f1574b4b010d965a6c111c9f66f5d8b7bc9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2eabcdbc5f817eac0d93ead870cad0f233d56499bdc6b63b9e0e46446b11b73bb2774a49c1b1ae4a855ec3361732e2d54acec9701a14e242eac99e227c1abf47841006ffc79cee545436f8e0f66a5c63e02193bd0d9599b3467d3a409d5aac12bb4a3a27261afe7d10c18db8e47a08ca22041deba6d54bb3f18fbefc8b71da6b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c5901bf37d24fb0520d37de0debd0389e54204d74aa1c117c1814a0afc7eec6c94a1c6f2c1265296615667fa78de6152a59e095a78d1b4b973a31504414305a4749c14b7b2ea853afe2f02289baca59f7071635af2a956019fcfa5e3d557c5c117df4494e283baef6301662d92d4965d18f602fa486e5ab4ac512a31b9e76d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8108ba05a46c0632afe149f2fe8ed463ab80c7c136495eb049efbc84d407a5e86df5aa591482f7d61af4963aa7001e3c28f43c37d0bab60b3c445c2c6da71919ce69d48f027b440dd07bffd05d43663956ff0e47e87ec2609e4bee0ccba568c16b9a8bc1a5488e033c32ba444ac4efa5c816bec60e52afa97febbeea7b4a89b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79b16b7e7f507effc52ebf76fde0e22926b9fcbcc589e52087805405399592ac8148f640ac1d0031af885f3c01b819eb844162f5e0f3b29dd552427a140c2eb9bf52fe2bacfad26192510cec3deff7edf73aaaae21f1659cf5a01715847cbfe6f327113cf0210095776e90e6c5e9a61dcb39482fc451e8b81650dd1d6b9e5623;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f8d245db49dcbd2e70e43f14c6c6ef5f908c9ea0ef19e89824eb0a6466db8903779fe87ff626bd743c7f1723cf4ab6582afa8376621b1f849f824fee8b65fcc6a097f8d5ce5dee28c131966f949db4c0d91d2809b042548f02a882408c29d9b07123ca7be0184707d23e0cf4a2e3ad9c146458f84178a20be6cd685704c52b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd348d8d26f10dc08d304f6b154ba9b5290a4a993ad0e7096341166516f57392380ec01dfbee082d52c9ad0191c2c5cea0a64bfb184b47ef6f71a9482098b6ed93850a0d642b31e996ba93617aeabee18fac8b6aaee8404866d6f1ed27a45f3a4c29ee4543969746f2804095deec844af3842dda3cedcf0766493d2dc0bebdca4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h700491035808eeabcd36bd8249d486131e36b4ee7d8d78294cd44b4d96b0e0ce43d0f0b656ba312e05c675b1a9ad676edb7a4579893be2abc1a9ecce8129c2c1eab0674518f1f3a1e186c0edc8dfa4d93eee0dc9151b328cdcc91a57f6d395a5a0380b0564901daefbc6d4199d939cc31486724ba12720f8225522bf0b4b87c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0daf6c93be5fe7c105c0b1eb4c43b005ecf67884d65fc7f7a9cccc500c2ac7a9805ca0b75da253ae54fae540f766fa159957534038edd4ed1195105dcf0eba381ee49d1e37dbe0cb9b26508f43527b3e5bc9b7a189cf17af8a8727d8eeaffc0b7fb8df99bd9006a62523ea7900bef42afcfd077a888c291da65c0a2f9875998;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha6720611e3522f62934b91507fe8e6be7a4cb5a545b6a21c8bd02f37aa3e12fa606168abe527fae69a17c9c1651d54082f0b47940b10329878e9e906a62e28d5185e5634c1e87b61bb98e7612d3ea9ab120b809773abc871d6cfc2d02b3e02524fabad3edac484ee4c6f93c8e156f5aa25cffef33693d7977a10737d4ac298d6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h80fe6dda0f48561b757ffed502eb05872c7e0f7ea1a343d1fe0280e24a599e5e93af3e182ebd59cd9dbdb16a0967404c2a523b9a026d02c6e11bb38ded42e1096d8acee1dae1d45c91a36a5a84a3686f37aad6e85bb257bb996aded7d016237c4aca5c5fa587cc60b66736d001f920977f60ea55ad376b3a5a4c82d7c7ae39e0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbfedfa40ca894ea5aa4968cecd10620f33be7f0a7ed877ff0fa731ebe63236230ee8f6fbc38a16ce1e2d4254f4c252328ef6c76771887c8c8bcc5c1f409acb2539a697e4b74bba04afba9d2cca639ea1c9ffbe5639d12477e82f9fc13ff2043953674523876d122faedbe3365250b0652f03ddd7b68000021a4aec6d5e5716;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h92379b741212adf210257ff4079e69014c9cab491537f1ed55f0508409d7471b617b7e77e74ac21c001a7efc25611da68545c7b96734a80248f0137ed00dd40d0610d14573d15ca88a61acb894b5ddfba2a919a94790fc6bcd27f858b5d94cf4647429b715ee93e7c482ed6ae2b6dac7e17ce7f11d523eb38cdb6f8e3dca571e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe7dae2637970ea15e6f895c9e4b0d0ca5dae070461636dcbd05031de29842cb64bd1f2fa0b78779672e752bd56e53586af7ec647a03cef55918b0722fb7842776b66cda834b732d41991112e0048c76eb3225d23cefb270c88f015bdf202cd92183c1a6e93e163fd49e026b1a381ab1a03c54a8281d9f659a8ad7fcf5de9d62;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81833088877ed99ffcca205b13d5cd31cc03ba1ba6337c5935dbfdeb8b4713d1923bc23726704bc98c6e0eeabccc4d14be1964cd2ed39a3a71837ab7e8d9a56eea23d5114d26e1331dd98cded8fa30b9a526b408012b471b3aab6fb2d80ab86db5bd3d513510f29c3d667a6afae3b0c88e0339650ce81e5ecf02ff0fbe98721d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c4f14a3549113a3733ecf96bf4329610072b3f0dfa83a76d457bcc12fa2c174055ebb3f1b1797dd5df3cbac370e8a66ebe09acb6c634428f38b7041460fcb5d28d416c0b19ee32ad8fc1aaadc3294087769282f14ec3bf94c85d52f3e0c4a46a297e01742f74a5327a5d91a1b26428cb9617e467b2fb58d04f0e4e2597484c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a0cb98b6a4108d35fa16004af4b50b515a75d6addecb95d9e48d71e1cb782dae74343e427c221ddfaa5427e2dc1007eef50d2ff0900d5185b40e41eb0d0b4fa9da5e943828c1499ff0131a20d46e2169223da22f2f80000b6858bf9c9b2c20ab5e789ab1e3ef6b0fcf6c1ef5f131a9c19ee21cacc59166ad236e4a5eaaef031;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88fee30fc8428f35b2074a045afd82a7dc6c9f028533cd73ba179378681e7f23dd8fa2999a2c9e9eb594ff0a8742178aa3260798127d467b57b9e1be6f013c5c8dfaffd1e17c6d6d4a1ecb647da17cfb21a38119c2c56bd205c5b67b1b4197733de3e88e61c951b768592b92d398471ade99b06d10d98b5753509ce69a0ea27;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc9a0f5e7c284ae52dc0337a5526f7c144299a820140b34f97bd3d6d931350a394f24bd0cbfaef2c2cd596ef059460671245d3f347670bade4a51a43e65e266c59fe651ce39245893ec13ae89ee66d48b91875999d8c56178be0e5330708c1a1e954e388fcfd358f2f48ba9ff3fe8a1d75e83a483504f549989e0177f12a20c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca92d0473716d8b6a888c35845f8ebef5ae5276c8d2bd5fce751f25605efb45c06980f7bfab8e76b9d68d51711db96df14a737c19e80b04c1be9c821ae56225a2818cb6cc81e5287c625d734c89fd56092daf767c5071192f69167f9d61025edca2d9206fc6b19a5202c7030075bc99740b416e09b64196c9927f952d9859e79;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f84f3b24d1d05486f5e6e1df9864106fefa8a4adf28df64e86b339ecc25bf57f77a74e0ce37f2a413850303466469a75c4c5ba64034e077a1998cff165f812ebb15774dd033e9ede340f0256eded62f65cfc71542096ff9b232ea3c5cbe80ac41ada10d680cca8a7a86906acacf948398f33d18d9a22e5880d0d05a4bf980fe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7008f22244338f45a66d81cac1b026bcca860d268161deef8ff649cbe1e5282bc9aa8ad7ff503e4641aeb8b0899e5d28fa33e0bf9469d21aa9ae475f688ec53720e4375601c302475d2249e4454bf334f87559ef4c654efc6f680e45a5357657d11c2febff61d364f1f509dd82e342bf294346b995ff857502e3b4848e90481e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9d7cc84969181d90d4bcd2aac26b575667ba30d352b4ee72cdffea85f8ee182526fc3ac0eb7b3a74ce782b9e2da34cf4c6a9c1f15e59ddcbb021a9122b906a1c96ffd805a50c1c528f60cbfad0cf4e2a1d50676ba06fcbbab9bbab09db7b44da7afe967c3cb18858a1db229e0d45c0785a170cd8ed415bace68b6f67688b0d7b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba4fc7569b696d4c39d6cb0ccc0270f90f811c99c86041ef75f2756cc29f7c2a9ba0f9fe48c7b8c051cc855eca2d06c55364bbfbae597beaf7520eda793280021fda2f29a6d9155894802cc5f46b6e8556b4f3da8b0e33a7ad58c0868c795a5046b31ea3a330fafd6cc4be2d75b71a1a7bad8f9c242f02576ef1a65d8b357227;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf414cc6537debea4e6763feaa7f16c59486a8f740e1879a9d13ee33836f832723e051a38a4843e25578c34204c9992b131fbba5cd70ae0817714509f954b45bff902a790f48c641e1ba504dbdc1d2812de0508cc205cb04b7321aca07add04e559e6f6ffc48f4cf9d6fb0782fc48d6669f361334d28aefc74bf9ca6c6e10668c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a076b97c23de87f0c01d042456bac7bd79b2e1e7e1a034c1bc16604a4226589af2634b81a8a9bdb31dd02e230bb5c321caffaa2d27fb981cc4e94e9a7985c3b17b7a707c1c624e9ab0e3c2fc44636ea7aa932ffa6a73d78797353fa07f3f318997b535f78feb972595be14e510238f88099f353fd6e9259697bdb476c6ebf37;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf24951ab091442773195826bf5400219e0ed6fc7392207fc94cd84f119bfbf3ffea49b88d2eab2afb233ff2b6767a43466d9252cede4e39d3f21a02fd88e8bb936428fba61acf58242278bae54239bc19c9e81d931653260d05a6f1475f476ebd9f366b0d8a9d2d8fddacafe3e1d980a88b133469331af7fbe4c540011422817;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a513108b7fcf479fe80b69cb9f327616ffa887569526a603c695e8b76d723ee60a5a1ebb1b331eaea0febaeb4815d91b9a053ee5eb689e404b5b8001b6ff3db17596074108909f65b248f4076d7f994c572f584c131a21a67cf9edf65aa751011ddb72602514eaed8ad9cac8c773708e64bd1787df01efe668583e5226870b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9fcde8c59825bdf60a2cd67bfc4b67d8c8ff98cb50a44831d3eaf1f40ef413ffe454ee064c522ed1e47afca34c71b56f8453d7fb255564ee1f757dbe3a608277630ef0ac8b1fbdd9e946afd1d6adf2f21e94b653d0c6db642b77492dbc8947b1313960d0d992b69a48c70c1daa50906c7bbdfe3759733d4ace393a58dd10f49e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10c59b37fbd9042ab2597e8bc3ac225c797d5c8726e3f25c3af6aa9090d0a4b7c8a935bbd271263ed30b2e313e80bb96a473a349c13aec368bc867ac190e1cda907e1ec08cffee4938a5b56510b68279c1e74a38284293ba244801d0cddad262ec24492dc92e62f2aa0205356df9e77ab0e29d09b8aff6c32551a8ae99ce5b27;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbee65635f34cbe484063d6879502ba732a0de06ae6999317b22ab933e177b54d7bf428b2908f6858a7c5d4a1d1085ca346e87347911ff6e1aba494e08b1b2276676d0225e382369310af7433c5a69754986602ca51c35e528bdfa09b611ac55fc9165bfb3aeaf956e5f8583e44d9f0f4dc60bde78086120afe30bced32507b70;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54330a13a08f000abd559d527c47704eb854889286d5797ad2891d26c5a910a87a37ac9a646b4690ef97aee3f3fa9fef81a8301ea68afc8c6be797223983bc4ee42fbbd9299380600ad78b7b80a0f9e04a72c2c6da2f6c9c42417b0ebf9cbf94d7f26ceb21a963960c30d892a406a4af0e26be11d2d5ff9d01970e9418c0bde1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1bf2e2eff75c50d8cac4fd57860c20fd0b6c3784977ae066cbce55cf81dfd8e1dc4afe80390c073cf1d2a0c203f9c99d0e64805f4fad6500d88db9348f8cd9b20a844b2dd9a984db9b1fcd4a6561fc020fc88a13dcc3569dd69f88bdc87d89b10cb9b616724372884e0e8107d081eb7073990a14900e7aad3fc0d295e44155d7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d4b7b43927366863820a0b0b0e7bbe9123ac5d7f047613f820c5832a1d4427fea6541a501dce24aa619489fcd32390feffbcb3f28b2c4519552e4e97520db1ccac03db5a7c909e001374f9391d44046bed85621032779a54e68f5d9753cba1540331202f1ef45888da28babcf8036d927c85d2c72447b69157bdab5feda1f41;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4537dbbeed1621db048ce8aac2342939d15dad1ad09a5861c061df37a24b928775586976ced0582c4abcf1e3b3a81cd4143238383aa0c30226dd1f9c739f11966ce9b18722145e32a773c2e1213515170071162f48af1e4764b76006dd25efd70481ac046388ec431066e029711b185a72c596003bd0525633cf401ad91a022;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h700d27abf42b9be8d937e4101e58591bf1242d511a44bbe6f2bc4a6865947b821c17c3a67085e77c960bcfc46ceb10e52147b23b9cf71cbeed1325f84c397763973ecdc4537de13b987686773b759b22ed184e76b9feb2822ebe071d91394b60b78b0769123cfb0aa75a8ed61b057d1d2c8464d9f88d72ddf788c5a3e4bedc23;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0922d5188d61964f62f61e5c921b217323044f47e11d201cade8695cb8c1d3c4a3a8af509d327eff42366ba055490e9e0207f1c334d4a2479a0e964942e4935c0883e4142e7465b862da322e18a4109c5bac25fe93f81d779b01baa79e0784b101142c3c4bd892717e88d23a3e3508ea280dae7307d418219e5e52a0ec1b4a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4283f198111da1c6602742217f25ef20b2ab2ab001d15f74522501d456e3d1763948dbfd0a200fad77817cf59b8678c20155331442d88e0899681b263acc0c01c299725ed15e732112f664243568380bd399f78aa9dbca363e4857c9a026e345758aeb6b9e0ec9b8aa7c6dcdd718d4f4e1bb6ea97525ff2bb632573202b3b466;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86b3d441bf904c46fed84a6f01c01c42cf781ebf25a6b32d44ef5288fdf3f38d58d566268065abd5f3564f559391f567a3f558966e151bdfca3f8880617add8c636259a8aa60f4a648afb3e4b347a386b245cc851d4a57359fd771961718a03380bc2dfe6d4eefdcf597c8f3509319aa3b8db3baa2e1d71b4c92f3c0ee8ea0e4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf9964ac11b9258669920ad1c14f50118ac68256f7309bc07ccb77ad27a3f620547006fbf973c5ae87640521318e7dbe8295bf8ce309cc8cdc2e0bea248305e035ca9a0bb22b0b1aaea78b51f8fcec276ee72b7ed3c6fe8074f43459d1a7382aa16e1232ae537dd6321ab68e8034a39e8ec6d8952f68f0fd8d1f8de63d94681e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0cf81edf4f293689cc3829bec9edb72038f4b5fa6a490f69791b2b0e462e478c1d317638228e3d37f3300396b3339912b4e47a8ba027264b58ac042175ddd538a4b55e556ebf0f87199492141c63527e0e1739d323f8f759eaec4cd8ad928b96b54f554027897d9438e5a61081a052bbb61fe83770216c41fe93228cc022597;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h728ada261af00456fe104808e6c66ad021e39fb53e2d98922d25219b29d56f137867ef73309199d55b134d9d56bbf18f19c067c2f39b9551f9444b39c6ecd330cf9ef213b4c0f2a3c7a91c9762b98ae7d0a3e22950ae86ebebea81de8930b608914cc07251320dee71a410d264b09ef2dc9ae16a63bb234d115b0110b4cdaedf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb900cc235f36ab21a2ab7f294b7052fad33e717171e56aee56862d110eb41f9ee010ecb43cd2369ed23481e7d4adb878974a3034625e74908a18190c6a68f09ad4ee0bf027c15a315a99198b3a83896c8326242207fae2cfeb8fb3785f871ab24356b1c9f74309a250ceece492117c58fe166bec1182098de33cd66d327229a8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7f3c17be48a1c3c53796b619e8c1fbabd4217a577fee8491ebebba6092d831de192d3544bccb30181feab59766fbbc5ea97ce3ce8518e5adc97fd6f5476e6d8ecac12eb61e3ca1c55d09e94946515bf024b942f974a5792a4c6864fb56b676ee3cb65c90262123d08c061df2093dbbcb577b240ccbe6b0e8cb25339e1b96da0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa51f69f7bc2f7b638a02839329bcd88e550c60d496e8128a328d825464f1c4a7f7351f632e184ec5d2afd8b04148787e5e02c25701e2dd888e97544722cccd3a3a84868ca725a8493d31f5c4d09cd8744079d771d5f51f8a99d58b55a4370c2e156bbff7d3daea2d0cdaaa8b2161d2306430d62dfdfb7f852c8222dc414c8c8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b90f1f10f45f140ec352a4e9058b3c343d60dd2e3f1c42cb24ed5c73f74c9a84b113fbeaf7fc5a836736b65b9fd3691b0aaaa4e2b6b64c619322d8be97466f847b9583222da2b276281084f4aeab9b8f225993779fe3bcae7d0919d480ae07c3ed1b922409502cca01e4c6c61a096513e19cf1bba9ac005c66fd13b13a27e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h683b1dc7ac7f327c8695774a651f1a8f8beb717c4a3f73bbf64c40047ed450e02035c7028b12d7159cdedb9782bcfb7e6ba9fcda1e10350f430013f11fc2a0e4a33edf663a7b0d9bcb4f32f76e7537e5998d0c3cc6f5d88de0729c8b0dc34b755468deb7e0af4b95d01e3ba53a16692798060b70012a6a14a41a65d545ab9398;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h206c6c0b7dc5760a1d9d83e98dfdfc3fab7d8ab6906b8e14b97bbb199de75154f18a2efc3a0170e4563e5ebbfe301063890746eb8826a942a4e077f1930504b7f8a2b7c984270831cd2b87276e99c786d36238f71831745124ae14a4c62c32aa1c709c0ae593c6493e560a5811d181588c14b49cc0a6d111cd128cb147b2dba5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h944424a98be120f48c3db3080272d36a9af7b74c93ffb4f98c5b27ab1c2548d9908c05bbde3fdfc69ad4a0e1d729a4dba0b8818e79ce9a5a9c39c8fca049547372a53b315a39139cd1232bc15df5596140278d02a70b3bd6292a28707f1ca442b6b3d3dcc01d987407dc176ab964941572bd128e74ab4c4d6f832450a501feae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3db1bd9a4b9e88b7ad6818455babc0e4658fb69235a8588da2f36c5323e9e9729ec9359e69e2fbc0e7384ef9687980a116983b71a77ba2ce80dd0bafe4a39a74e3ed4b2c0c525939cf005e381d7b39d04ab64dde76e1e65104c5f38dcf0ea97360e954ddd656daf653a3c010aef75236a5271840acd69395133fca7824389913;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4abf24b4eaf587bb37c02c99c241a24e6e1c8353182a0c5f890b1b5d004e07c3279db3d4503e51806b59d562bca03eb5610f77b1898885f1b1f9036769924d090595f4ada8b94976ba43fa272510c0607d8c4a6f12da7b95d6e7f90ca019442a91b7a9dd1bb414e64cc18235503ab04c87f801a47153888b741ed3b48db8b89c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdfb200e439936b4a41fe8303308485415f9ec506c6bb47ff7f715ee94e56b430e6d3139c72730c8c0539c652a65375d58c4b13aa2dcdb23bb0bc31e0954357388752813c49b4df24d564fb341f585d42dadc8d6b3f72a5157640acff1ed26b44909adc83dc3c1b2932e2c7276b0f957a49a3a0f36480e6ce8249d3835a50f544;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha94422d858e4b9136ba4ef0c5cd2e2c21e1a886ce1e2f98f960148042db6ede28085cdb6e870d4697e0240b4cdcb882de4148c999a53c6a4a3fafdab677618dc528c1229d15b78dd64f3d0bec5130a5636b1c860a53995630fae52381597fa1f5161af5b18cc115c074f77ab809039c2bc9a0366a35a454d3f6ff165a3ff4c1a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c89e154b1d48ffe7ebdf422834be7177c91c7a8ca4bc9690283f473767722e937e42a1d77995868c2e38f58eb5f9f1d60e0fcf8d80227b6ed6c70ec233920f0febdb2e59782193ddc5b2a6149171feaa85debc3bdcaad38607b4d36863193448397947c30f34b084f5bc3fd5513f78a818a35797172b8acfcab98878421983d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha97711d5ee5d65770e52b41e9b9e43feb68c8fad84d6af213efa245c91dcf51876c637f93918072ba347143c3b42bb38f1a28139c989bb84dcdfe8a37cb1263c350a2417c48021a474d50e00a8304004d51fbb2e897e45d283b5be43843e0831acaf9663e76f3a3cef098a098695959ab05c5586d0f432806a4d460c65d6447e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8431b7b7eb73f7392dcba21bee36b5be9d77998ba2da0c0a3ea9f6f13336211c298718cea79364bbdd18da0ed30a60be30b210aaaf3467556dd33b64d930b50add7a97fef3a1a4e0d7721a66837f4c0f506eae44b50d6634c7fea49c622c927b0cedcf837d13fd611ccb731a1b529df9dabde93916aa383514a0b7502f508f3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1f3a4fb78e5d6e03fc72cf5f78e331db29eea77a640f1ea725660d6c2de769a87e746d6438d6c6b4516cb003c6ad82244fdf5586b4d3bce199176a044e2ba201666b47af7d9a1941935c60c0199bb31860d942f7f403295311a6f9474cab1dec9fd819eebb5a930be6bf51566a6f2976d5960312b13dfc43086dd18b1fcea6b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c756e0cbb9582258173495f6327fa72cfec92eb28fd8ecc1d76a9bb9ca2e4066ff3ccc7df9747358de7bb8f89621bf245c9de3db27affa93e5619cdf1ca22f6118337cbb515c684d7d4ad112e2bf82b734821a9038f48b27f8820ab23ebedf3f9ea757f1982d56a1cb9df09aaa81da41439d2eec2d746ef1bea482ba7a06e8c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c0a88befe869690a53646999d7775940b9a1bc0f0124b5fc671850c4a5a113e07bd69baf19a4023c967ec15e078adda8c6b8badc12ec77cbe9d23901a4daacb43bef3cb1a98cfa01778929c2c460530bcbe6b2b66111c54f427523e50a9b5a96e710620e4460b0c4ca698666f01ccbcb845bb67059b4bd9cea095719869fc85;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1721468263c36d37115b47e5fb82f47e63c8be47a9e7a7814e48c826558fd3757ef076eff67744f49c2ff2e6b35068594e8a42de7e8a41da6395030a98b5f3666e212bdf2212c2364555bf9c3a11d3c3ae842b9e1eb10caf9965e2e60c1f7a9abad9b32288c3d2f93fe3b2739a1e938523c56f62fbafecf7044cb665e6dc80a1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f9630adb5f668e9f74695f3bd5d7093d1aa77d96bada9c90456fc7624e8ed6c2df38061f942f17df903dabf7559b607b0b8c2082bcdb3266ecbfd12bb1c5ad56ab5e3becab442c02a1921345ac7858bf6b4e30d3a8daa29b9aa4889bf9f62c78291e2174ea6f1c6ede20dcef16d7a079d590137ad4c4da89db5be062815e7b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6cbfa762c4e9c7ab8c377f593bb67b556d93103266250c72e4b854e4d9cd150fe7c416a06e2094896961ed0ddde6bbd3c6f26efd4e8928b1971cf1baf2ee897ad11717b1d5c5e986718b1c7077386120253fb493b5e1b010ccfb52de34a1660cbbc8d4b244d8c2f337eeb294e2933b1ac63143098e9ec51364ac8a9f9d599ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5798592e65a8227b0345dfa6acfda44b36c6783a7ae32667dd16fbcd715c5c06788b9a9eef5cfb3a61e40968c777429dbec4aee2ce98b41de43bafb4ac08e35240d8bbfad7779fb671f33857790fe297ecd50bb36a45160375d2c0b2c4665fb8e793638c2acbcabbd02b58ca21675df7b2911d4ba97f679f497a6e97f39a29f8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha06467a68617d9d7f7b64c710dccbbc946a956e4f4d357e6819040656326d52cd017adc51f5c625da86b266c8f859770aa7a258f79f7f8276e2679b719dd3fdcfe02847bc580464958cd1236de96822eaf88ed39584d7a243c71f0dd0bc9d3f5a24a6e024216ecd0b54695c7cbb53d04138cf17fbaf4ac03064fce6d2725c9b8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee294c4cb305fdf0f769ab4750c3fd873d26b7c71ce61b4e56365844cbe81c9a14ebf861c7dd4c6ce024a6a53a5a20d816802c963777cd0c6a63ab3fbcff6ab6dfa4c4f88b4cfc29a9528ef1ddf265a8b41798cc32675697a96cf664414b699f79700184c226c272fb4b5fbadb333ed0b075a7c27f0a9c96655d63776c518f18;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1fa058d801e057fe3bf16258271c2e786b4f066cdefad65e18a962c20d482a11893c96e657dfd2fda1c6d2651e91cac9a10bf9ef78f82c047010f1f13efc093b5fd3072059bd7fa4db4fc4c5bac70f48fd85d2af365f3b65dc3ea1939cd2f1ec38ccf6ccf2997b94598396808507003e54a0d136221422f0f6f12929bc949a9b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf8ee1742140c24fedc7e555baac90c56fb8241e22f43e77dbb830695252202cd0c878e3d9e5954cb9afb47b6a6e94dce83ed4b0ffe1ebcf40d0e8dee7a730b146f7ccb61a3f9837c077051a243b945642f4e08d0f4745a15ca299a3c692189af04cc2a30404356c2b27c7a3cc9e8362a1d4dd852e3cf474b7f219b32101382b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12b65389d5b63c296fe091b05b4de1b2bca49e160f08f0f684d4a6bb98830dfbab9aca4d8b66dd15840e4f546971b506540f0db0f450a1be02b81fd8296d3a57d957e18fd595ca4d2f350eba76396da62d95b2c07d4237cc203110820b4b4519d1dc3c50e92d9091fb0b25f2a5237fef68b60b616d00eceabaa91a60797647c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61463b8869a0d8d8cf40483e93dfb565b2d15e94910e11d6b1234e98939364289b79527706c8ba5d6149d0f94ccc17af9dbb0c6641ce25f4abbde56129b12cedafaf690b977f315bc74eb93336825dd6e26e97264096f2af1d7240828f07eca56392ecb0a3a32ccf84f0d935349a90835736f918163a9566e6597bdd1adba60c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4345dd995d407441aef5c4e8fef6e5aaaada5bfcd29e7bff5cc34e2d99f83910fdcb11dd95de72ddaeff2c61a0521e2bed4cc38cd29083f8c0aefe485d5c0897fbdb13e8cd2b464817237732ea66bf2c75a376e463643476931bca2f4e0d6fab16e09bcc9d924769c57f8c6c1295d8349ddd9f2324d26dd8d94c7600ab51d3e0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a810b91a188090eab4b1de07bca4f9171815431b1eb1a54f1190ea0214bfcd7c57a02b2fe790b08106491127d2d48a8cadaf993fa32b90c05e59fb45dd9ef3dbcc306bca87d6c12c78813bdd740363532f8e95fea68ab59706c2abaeba345f6b7b94252bdbfcfe3f21320194de0ed4c38f3ccdc6bd5b984b66fb7be1d0d5d03;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h217d8927cc3a56bd0a8d5ded26bf428c60b9b2f64bc1ed2a8d07d20cda6e8de674d6bc303938fe2a8390c4bafeb0542038b648a0156c9c7de07530534e94548a3cd7734b2928cc6a8d71ec695bd46060a2f393cee0a741f0f1dc3eb9114fd41b7e41d05372d3f293b19b0982919a06c70562aeafaa5c1b6165a3c0f55c169f94;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7270b9f2eca1492a30c0e31e4ad1b488fa5ff85215b691743f0a95fad4381c223141ee5a9a52e5c0f3c508c65714b07b544c331efd6ad263708fc9219e69922d10912ee6998ac9586218be6366f3daeec3fba3a9f430bf3f37197d99642273ad642350356a7f6bd8535b9dab75aa0455c9f0a6f1689c89a8c2aa709520db4433;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c6867a7b44c50fa7adea1e155a606be845b69107defba0877e43cf2c11f5baae9d11b6e50f2163f6353849e11687ce04881185ed3ac5e91508f718483af123e457004c0e5e47e869076f932fc8621e6e7daed506e0975d7973c4fec28c8346bccbd5480d418c89eca9e82d6d08d1f3af8c2683109230d7ab0f3e4fbabb09203;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd693523b15e52d63c257940000423cdf7f773d873dc8ace6b8c59b0eb2a117309e9039cebb750d6e406cbfe1cf60bddfe2fdf4f506421441becb9e86a2af035a3456f09c73794c7452c9898faa7927b33fd58d4b2b77ac66a421ad31c59ec475945ba8261779d95d3322bfd769cb162063356c1364097673b5844250afebe1ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1b3e66050144a065bf625a9694a885ef9e09d681299c90d2a9d43825869ece330033e0b8e3ab3c279a56daf60a5b81c940bb302ef4874dd02214c5163de2bbeae0dddba2472f76df44c14aa9db9bc5c6bb666ba2a41716d5c6785a8e66324c6ce37b0f544aaf50240abb25840da227859e9e00c7fa42aca91a69e1548e88fb4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2cc0b2ae7389460f24df420978332a75be03d8fadba686e22f0b3e692e719b1a50985225caeacea4dc6fd205cc5e4ca0368b74959e5a001260925b4ba9338305b83de28831db97ed085635662e5fb366d0b6859d7977e5b5876315dc2fed336d216d907b7d633d6f117dd60906319f65f52fdf51feee9da2c1ef0a697e9ac12f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9e0fc062b20a896f5d2c8c558747cda9280249c7b765d5e6522ab475a3de6f8e35262d73b120a1a8c78736625d421f78bab112144df91a7657cb22b7e0d1dcee7d143fb75b2032f0c1c28623f1c14e8a0bdb35246ae35d35a8ec7754f2810e672bfb077b14b1fac43c85b0cf1c553ee48236e260fa3b98e45fe6ab232a0dd68;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e7eba1e2c67c800b3fe4111b016321952f96c365ac398328e40f9d053cc555536bd04bf5516bcece266e638ee10a62ee784f51039557b7c3ac729d3bb513c824d78ce0e83e9cabcc22781bbf42f33f725c2ec7cd95808d5be76dee990959f191b56d61e6dbe004903ad9c551383720dc19d5c6fa0c1d3c4f2ace57d8a8e2bd9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc58b486c80dbf85140ff0cf4932aae3cc02a01fcb38dd23e0acd248f0e9105d678e003ae49df3fa8880800d71ba0810179b62269115c5332213e9cf1a333fc290faa71c37dda1494ce5e81efd7b4746b399adefa9cb86018d939bb2d33b9bd87e70fd622687a21f6fc5e168ac80774de4e1726a180ca7ef3db94734da6c2cc2d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hddbb1a9ad2343e5360602b73ee4968ddfed52b8721e04f2ddb413e0d3b5ef2658f907cedff4c161022e952397b7695dc0c607f1465e2e844594c55a2d0488675bc0c91b46ebc2d871dfeb082896dbcc5208c03b35d48020197e3f63cbe7114c970a02cb67b24d0f1a0da13810a1bf5082c64ebad53b5999985ce45bbaa0b28cb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9dde4ad2044ab25a7440620aad2677117c5ff00b63df9e5b6f7d95f07ad3bd1939cc3035ffa807b003fe0e07d379cec0c912f49e5c141b09dc0f7683a68b1ae900402721f50d131ba671034e831a74d07c3dc6d44ac6355af23a0f5f06665dfffda6715fab931ab6f24bfa153c0c0dd8e115a76da3ceb74527bb3b9a8ee3ca56;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23ef05467c3edf5f52f607505cc8bc32c7b6d43bd6b91dfdfdc9a22bce5670ee179f226aa53be3e00a0e1aff7ed036d666bfb8f23c234a39de8774cf61724d7f48607502773c6173ada006f642a736cdab96973fc9cf7292625022256b771a1fcdb5acbd0feca8e7dd506a71cb2e05162bcd19c0677b32926b9a99d95ff8bcb3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc115933b6e25c6ea840fa886753e7c2c7b52154baba44b2bd901f369a6357cbe06ea96b8a42e354a3a04eb0b08c93c553a7d27173c5157c5042a0ae6f66d76b5e05f615b4a88cd943d99598def92785ebe990166af189b5e1cb275b996239ffe3dc4b7f965860754208b09c35f46dfd2d351738aff97bcfbe0eb4a76e427e3f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd33b5a9650829734531ef478365a9f5330933d34093c39a81902bb79faf3c2e9082407353237c431a96a412d5445fd2af20352e1aef44330c7c9b6e9f20fb405d3c9e1cd37860ef5a6349bd689ebcfea8ee9e492fc14a2cc374988ab29d022f9b58c72fc1f042049286cc6b5bff592409d32b3f78b21e716faf06e13300442;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82ce3b58dfc45115926a521ea60ff9b5e72b6720ba0a920b16a1e35132bdcdb8c4141ed8f45ec0e70e30407146f1532d548247ea751c7c3b22d21b66d081e62d83b72d37736c83d929be2c8ae7fc6350b1f509595a05aee8b7715f92523f14c91929d47a69d9dd23e1121bc44d90942df211ef0ed47e7f5954f21e02f737e2f8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd302ac704c49e71219d253053ad65dc1bb8ce664fb487e7ec788ef46dbca7abd7052a5fd673cfe1a8ad8128fb370f996ed24785d96307b264fd3a5f6f3527f4d5229aa43756cbd849d266860bb36a99312f260e87482a78b69b1e5befdd86ec6e5f7294e0bc4b2e1cad9d1594eaf7e97e77e75be34c9daf7c656a9d78076a144;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c70118845f715acc66203ee2a715cdeb7c784f1173609fa151aa911269c5cb579dc393f4e80192a3f627601154be4fb183141063512d4f8d4f9d55bdd7323f6d1ec70f479ef1635f5f624c88df68511ef547187c0f8af329a0994439ab7fedad20b1633c39d5a6e729fa5b51333285a52a80e15c63bab5bf1a9a7792ad8e3ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf2e3e3405be98191affcb98647655bcec12ee4b6408bab77507760ca5f47fe2c55a6b9c9b160190f871455e2fde5c430163c2af72f5dfc81c7b03dead9bf4833ffff71b886ffbaf9751e003854053ae17ef584663caeac5adca683b5c9be0a065cfbdeff9fa32a9d88105fa448423b58860f6c612610061cbe49d480379a973;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h147f026c4bfccc84247fad0f9270dca920eed6192f5be8fe40e9fc80851c2e36a8ea3dddac26a5089ab3bd756a3292c8c5d30b68dbc002ddeb911e0941a374ac95c1d8cbc1b683c576ee10112bfb91114e3d24fd71e367d92741bb2c425cf046b43aeee5bfc38818f568bfe74bcd5762f0c543edc35a66d97593dd3b41e83505;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8bd92a2d2b83c926cb826df9c787926af811eafd85588b6db97b09673c4649a0232ad94da3f6bd4d639add6543cf3b704cd55af32e5a94cbb648874f4936acda72b7f9647c14758702521c6ae63fac97bcf2f0f24097c48d8e0369658f8e2c3ae67381ec9e3366c8c2904d6ee0c0fb13006deb85cc5c3b6ef5a89732b8506e3a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42cf00a8835ddf7890b6bb46a6b3207ef64fd2fb1a6ccf29d2c84307115ffefdddbbb8e338c09d56f91a2ebd3ed2fc3ff651caf4f7bc2f76a5bf9e98fcefdd1325fbf61d7c24ff51fd2720d47991bbe0d052d856f16b82c2ec4c66a5b85fba7f70cc5960ea5f41600efceb149143b7c273fd4baa9b02d1eab618dea02b74df5d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4498d0302fa66eb3c0d32fb505f51d3b7d7a6d330cac46b0c881840a91ec87bf7f8a7823157e4cbc695d4a84cd8b2822cdff67169c13ddb5c8afa75c4815bd3e94b1657fe36b29e02b431b996599faaf87cba6cec978bd8fbd889e15d21069f1b8381ed75ade7afca273267d1773c5e93554561be8f7ba430de2076846ee3682;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66493305d342e04a6b0fd7c7d15a2a7e8cc66197239a3cdeaccb17ff5310adc558be0530d49577e970f12c4009b7e6043b385764e69bfbc94e3709f5e9c9a19d0be14ffe6b993cc81fed29561e7f2edca04b228109c553fabe367c367c5dd8ff29facedfbd158f8f0d82104e609fdc6321e2c94cf3dd3c9f324938246c8d6ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h557a99287edbc881ff0a5b18450088812627c564ac5781461f3226238336cd78de6f3b9b815163953aac8db4cef361b0dd84f200fa787c48eca46487a618edf3ecae71900bca2d4e3e0bd35811d222e1e03267f3330fac355e49697709291397ee202697322b1a52d94795b53a1f5eb72efe73bcc11a8720405400331cf70c02;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he6a2bf211bfcd75e405ab5cf717a9d580f3e872b64fb4c8945911eb6b6471322675f8d218b7d1dcc98445eb5a68f7c026e281445b973858cec4f399cae6773a00446695a29442d248ce6f512175357542b0b12ad56b8887ed7e69ab24e8d1eaff48c458d7698600bc8e744d6fde72552091413382a6769872e75aee7751e4fec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h307811979a152a94942ac888bae0e59d6a3c99a6e3722f6a5379c28f5e45f13364c61e1587e5e3c1f1910bef098cb694d42718c6f9a095ae6db083496b710afaab24459dd4d8eba786461d48e4f57163df3733f3b656679879249119f439dc55dc0975f6ef9be53c383c06a3f9e22664d6a9c90a7151e153eff36786608bd29d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c1397d9175449da4fdab61528006eeeac43b8656fe40333bacd2ed08acc2916562a62c26dd9bdf87bb59895a2d02ba007940708d0c6623b9f37c73d08faafd1d29796bbbe2572633d42ec1948e18c5a06c089e0a6dd9127aa66631e2484ab609a1a64e2bba78c3eb8a0670b881b9e93419f27402f62d5e490b76a274f77c5d9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57d79a18caedc151b84fdde370a7be9a6e158fa6976d4af3d14f3190870fd81e8405c49977b4d33b86cd78a54348e3149430d52ae548a70043703cb1c2505b9592c9bc771080932ff132d4524de3a14c6e9ca999eabf2494aa3531f64114d71b5aa79f4e614073f55bfeda6670ced0e5e490ece50617fb24d4d59f5d22142e1d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78fdee647e76c01feecb4eab58bf18067873eced49b7046dc0d5b21d717c004e49cefe935eb4a1b84e0bde1c6888ef1c8928d3cfdfca45740b770186ccc4a21bc634c09d4113bbb797757eb2aa1617fe57372f70a2d51231fce782075291e81f3f777d170c88d2e67a7dd8cd6d0d9be553b8207d9d80c82d1a7266d00056ea86;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he0a1525bbe3b8898143936dbf2cdc6d8aca783ea883cb0cf0b3176e7d085dbcf287f1a7b2bb77481caeb5e83965d752d532616d2384714c7f3432cd8ab2d12b7d768d910c57d9b510612ca798126daa5c45eaf924e70a14ed4b2a29d3996c39ad6f71c7b06e792ef0ee265d39d31fbbb8325c57f62fb055e65d122dbaf818200;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c2b16508abf733c950bdfe7e5c600eb37e9c43fc19d9a8c617474f296fd9d6808a6c16f0b4562b569f5d644aeb02dbfafcf772539aaedd0b540735347d9538f01f8939fd100f5f1e47f59349f80d9edbcfe346cd60d795d9e35f2129f41f57df3c52a725eb7a36a5144039fa637db3eb70a8a22daa3417e10fdb48b37f22278;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h627b7d0e327a82804590ee99bf8299a12ac7cfc8769c8c84a3363ee6ece530eec773830d26a8bb7a760dd3276028904bd80067b629a1f41c25dfb2882cbd55a464e988ba3d653571dcf2522d9af2c8fa00633e5c7c85d110804cc9b28afcfeacb062fa9ea3826d7e0050d075c17d79c76071159f0c0998844459db4527368b64;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2273f8fa4b6eb81535bd448816789e36aae01996ac30db693adde77d24f5ad1a41091b9b5d2c421ef9223f3a61738fa116d7ae4a33c31407f9b2964d1e3beed4d7e4947b1059b78b73d1ea2b77f12f831dbb809c0901d39a58512bca7fb66575514f384ec89de7665d2bac4d8cc4d0ed33c666406caa0ead9e7c3e2f5ca4ef03;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a2f04f3da17c2ac21b01e213d3c651c263479191ce272660d4bf3e3882704a97890ed9657e7160c91e22e2f2f9f89c2840e43e1651db0d10d851692016573f4aa5e42bf51b9b96aa1918f3f98b71b07627f3247365c7e05d120674ab2d50ab62cce7e342ff4e056fe88c0a74bb964d1ad6a9b889d31e71d18d853f8da8bc9b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h968a0b5700a40b95c93b916e40b0452bb4a360e9497e4a52170d5701b0c80f243be6d261cbbc9c4c435467543cd7b649d063f925963c3ce65f10b309092d392b1e56815dca23ac57f5fc34f56a37fd12ea9aff6b3ed40dd3be9f8cc2d0e8c556be6e226eadb7898409237ea1cba45ef95ab171d9d74506ead09bfcf2683e2905;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h813514fd0da6d241b414d31eb27fff5bd71af37800ce1132719018c49e6a2d98723a1bf989d36da464f7cec5f977d12f0ab641063129b75c6f8a63660873beeab2a1584a95b532b714519327a7753dfc5ce8a9c8e953f47673b9c8d43f6893bda985d245c6c4ad666c6c1ab88186eae303dd7f58c33f43a2d0ce2ecd714c6ded;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b55d4b7572c94df5fb0d5ed39f208181bd662ce06eec791d47ef7d998a01bf11ddc12ccb05e7313de373fe85cce9995a9f76235e6061a8b65eb37020a7aee893c45dfeac99cf503bdadb110822ae28fd49865851cf0ac59a1ee9f51a31a1fbaaab1e54a335bb18013f926343eb65fc360e0ec8082fb92b09001dd1e25f10982;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa793fbea096fb66877289be83df891eab7d731cc5974317214ecdba9a298530802b7ae162a85954b13395ca1fbccf9c812d55f9d1e81366165efec631e8f310af7386870044bd6c1abc550b36d3f42ae160aca48474238e745260a2e464c77002068d2f42995b86693fef7f496ce9f6ff8121a817ca847cb5b27a9b472ac3ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e1966b729b47004e03b36d250885a805df317be2b08c0f1600c1c084127640051eedab601f6a887e232f530d2713829b11ddf716a858e358d6a9eb5308b08f28f626555ad63cf341747bf80cda74643d0c014332d78f88512cf0413d70ea26b80a9c66963319c1646aa5e5f4577b065fc3fdb4b57619a9e80d7838e47d11b36;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa284d304b3258be0ccdf89d0f72d1772e946bd44fb8ba1aacec9e5ac474bd819b1a979a1e3239da709d918d84aad9ed449b5265f2edaa4d80f48cb92d5cf590f50ce2101bb73be7a8f3eba3924b4b28474c20f87359e90133790f78d31a62f685cc6b215aebc5d3d6bc502b650fb90be4d07df210bc7d2b840670bee7d25cea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6beb7c4e38bba87bbc04837b7818f654d844f3fdac5fd2dc76f13d62b1b14e2b61b5c5a010b3831d0d49f21f17e0c05ec1d911e2260a2b001697f1efed465e98c34b2b37240661f74d353430298cefbdcbd672f3a7b1083c882c786e5c12232392078e5c5ec875e3067ec4ed059e9e9090b624dc97bb1a7e2e82940ed37d65a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc109bece23635fcbf045eb6c5b55200502d6eb955aaaaca8dc1ad655d0af7987caf6828f1d92bd1bb8b19f7f9b46b68416296d2652bbc8f6f27377c16e726ef8c6f83f93d2f9a03ea7c67e4674d19f2f41023e4c30715ea8a135f8f670afd47f141b8ef770a9563488f7eab95d15cb9a3bb05073aacafa07c03649f42c419fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa5de2b0ca142d07287172b14188c9e07f1aa6b2991ac1ff34ce6262af875114a7bc74dc4ab8022c725bb3fcd457666e6b8b8d1a6166ba87fd68d4a2b390089b70c2022ff63613aa7815fecc5bc52d4256712f3532b0558520c4dc943a821165d728a57d13852769c368ba473347fa245d105ee66790154d0672bfa39c85ba3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc7ca0bb37f88b4648055eb8feba4555a283a6c5c9d098cfb4d946c5a565f1d8ea5cda21a05291037d88f29f3aaa96faf5a03fff4b886e262ce92a9412d162a5ac689d9f9d3e0b51a7f1afe15bafdf1a4ae57b0a843b6b24eecaa0f427c941dbe84ff9e1352bd87eda351a31d61598f5885bc9c7ca3efa7d42230c0a92c8460;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd087940b090e22bb10669719e750a56d29e188e9ff780c15f3fa7243a4387b169f22fec8e26b673dd3d447d42210ed7314267030ae0799510081f70dd4dd469a02b92288b06e1788b6022e947fa030d04a96b35a6bfe29b762f16d2d6e3d712d52232eb8a9287d733e4ac412d7bc37e1368f1d09a21dd10b370951d62636d89c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7844665f0def3fc3faac1e2dde517566bf830634ad02212c5e5289cc8f6d415fb0859e90409915e0ad67841dbc3ea1ccd03c831c89183c12163ad739955d4d49781a4434abf23e729681df2c14fb03b7d0d2a8c28447f692a357078ab84b2d6f3a066444234570b3d0d3203e23305f884eefcc479ba2935ccae840f0d7df0fac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4eb1cbab1d14a6f37ee4cd2cf517dbbd954456ddeb3125be6f3e246de562df821924fbb7af9f5f3b0d1cb0c3916a224181637007788b4f42ef19643208ffc494f12101858b5f1b944e79d056d4d78a474e90b0b12d872480b758fea23ee64af484a36a785c4760ca89b649bc64452ca1da97e20d617d9761c36ea732dd382897;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd1322df13e2612676d38cedb315a5a882a6219ef306b8b0ec6ba642676a9093c9d85928efb3bf4e48652f764ce448a6c8aa8832094962e9cab4e6c6166b549d876cc278b645bb560d389ca5704aa2c8c36a64d0ccffe02d81882719982fd4fc19be65fe63e5c7836ae6ab82b2e7bf5f000a4e586139ddd7a3d3b2941c8c3b3c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h196b6e0a9de21efd99b4cbf4ef1c6a67ce5661869bcc6bb5395e9ddc1de1555ce99590d8bffa1976ca782fcc3ad85e6bf30ccc931fdeacc980003dd12c73b5eda3717cab8ca884b15de7ea864e0abb8a31c12ad497d117fbd742865e99839706936ef79b1ce952b9ca950982c7f753a8ce13497d1a9ae089b35ec18d9062d18c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7970c499e1845768bfdcf75c3e6fa1eb5916e1ba06462b36bebe626ad614628f23343e4cbc67e29f1521b2a442de961b26effb181cc2412c436154fad79102cc3d43e7c6cbb850a5f2a0150599dea5a828521c810e7da61993bfc8b8e7be5fb5a0b2ffbd66c0014145afa946a071677f8caef26410e084f77e7a1b375d22b21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b4b8951b387168a88257c7c605f6aeae5b1a60a3abce2222d8d50f614ff6947530fb59cac2c4032b9b1b6194bb2bb2a53088d44f3ae4c24be386bc40023f07d555edd973d9da01922095cafb6eed5332a8c41c47310f7f5b0353bc32357bed6831a34a39ef5e11f77720fc2ae2ac51e80eb922ffdcc199773f17cdff6ff8c72;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8cd5d9aa69545af3f77c772e0ea80ba83dd6f47aeebdcd1e7a35a20bb0aa2492d44024fb8bfe90c19a0ca7bd35617387ab3ff59a6099f70a2899b68998ea170ff178a7e81f1d044b1cbc0f34786713e926039812affd2b5d87e1cd1a7cae19a10c0c0fd874eb8d9cf553e4f200cdfdfe5c023537337596d0e897b01bf63e792b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e8cd624dc5d58de60a4809bad4e44a28ee1e302fce0e16174d0cd370aa4b3419efa4ee42f9936b986c81ebb1fed14db175862d6f6c71295342b50cba6f5419cf9b0acc34d8c6344ff653246e88915f9498df7f7ab3ab4f5a69dc46aed781c5dfa490329f8387f041d0fd97adcb11e93d2cc759479c80d9d1649417c5864735;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h684c9a7b7fbaaafdf7eeb7f90a22370bb1e1804ef7ec98baf1408ea97e800de1b6db380e4ec07015b2725cfbfe91bef0b5e2d41285e51c2ebc7a1834ba87f0c6861e0ff9650e47faf1695f925301330fc6119c0b09875da28338dadaba2b6c8c561141353636bb241f0090503ecd3a5f43d94db3166cfddfba2bb3803e61f7e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha440b6b658e6147da40bb599582174bcdbbaba98d935e60caf8d02752eedbb0ffa0189c301c4bbb6516d87ce36fb50ed7bcf49fb3b2784d164fafd898bfe7e6076c141812e91da13995cd93abd713c3112f20d31369a44e64408f41368a4b8e7076a8b60c049070a13295b62a9d581f66797873807155833cfd297c5e804947;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha8dc8e42f2ec2069bdcabf7d0281368908318bfefc45c3e61110978cabd33246a456f2d02e71b9f0e63226c54f163143d9f355267b6371803324d436388c577cd153b8ef6bfdbb6c65b4ef21d0dd1a802adb16a995da7a31ebf1e8188b8af8008d9b825b9ea9e9cf5bf2c35ab0d0a069e6f05934dfb7f9cfd32da410060cbdd9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb53addca28e8593f6289099a107b018e692bdf362c8b278a8b70b7027afd73c140eeea3a96b35955d342e385ce7bbf79490137e7785aeb5beee78e325dd1b2b8f197288a1dced2cd5665bfe23b2a9170283f90a49a349c4892da4d81001136b866229d14ff88e4e06d67b6872e3f1414664d5e78ae5d52792933cf0defb2dad7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h252ab4e9b7c0f877063767f968f882152adaa6904b266c17b5ffb5672b637f0cecf66792cc270b810f3689c66a021e105f88592f832264f4acda65eede16f2e4ecac811df06b22e4e34a02ddbb7c899c91763a250e7df1f09bd8e1ec0ed9c8585457f1ee27ba34d574a091fe1e1df0d492bc314313bf38b953f590b45e47ac1b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc04c2784b1f02bc0727066c02ba9a6293d97563f64d556776ea09a6e1b31b5fa8771c54fb2be767d466728b6b50ee20d3caf494a26ffcad78371d26a395f49f1f2275de25edd971ad9ef731da582b89f44ffef8a32de9c091b0b377273c992efcb6967f84a7c9964889dffcdcc9b9c52f06ec97b7032bf84860da1d1496f257;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h786c813be86e248ff73ebcb083063942a16f081b5ae0fe29aebd46682013a81ed70e943c1059d674b7b043590efe64a5a581318f9c8d7fc2ec08114c025769a61f58929471ed3933bbcb9639ef38269159e3affdda167f316c4ddbe48431878ed4c022ed1936e1494340d283d60bf6b7cc898b7a32ad854a56117647debb8628;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb99a8bbd422b53058fc67ea8e92733e3d3d481965b901586bf4a95e29d858cbbc5cdbd6cf401484bd62ff85d850c795f4ba27e2d6f0bf8b4128eeb7f089cad7e4bd78de87b6fb102d13b9b12ad547cd8dd3cdef30e510b7d8466be7c6a41c6eb2c4ad89fc9dbb185c0e5598ec666bcb64c8c34200b05a6a6327f1d68750ebf7a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a7b5117aee3299071aef2403f03b9d62cb51386a075893038d6e1b8a2e74347ca6358343309f924ea0c9af66c680d71dc3e973fc37891839452cd39df21294646811bdb1a3da53c9a5f012fa530aa7051cf0e188388cf8623a8d20a575ec5422c5880a66679abad7e0745b797b3d3a11dd78f70881838ff9833f8b0ddc0290;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f6236b6e3309fb235043bb27b87d0cb1230f4571a6b1c4894c850fbb7e03076ff461cc8e80e3104243a682b0a7299b9ee07130203e47c0f4de45abd35f2b89d6c0d0f02dd7768fd45cbd88d043ba7683b486274b47b0c4e932c9a943285cffb59f3c76233784bc54d0a72ad2c6564d0dfc8a37263d4ce742478a5cee0efad83;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h438cfc6ebae3741f6a550e4792b1ad347e072c3f1da1b153271cf5ce8bbe7c89a1271a89f8486707212c2ede054d3865c20045c171b9d77f8ce9016765f0a0a60c30bd7e09f7755cdaca57b6f0f4327f8172aa38e8e19267a40334d216805fcd9b3273f6dea483049ca2ddd817db4297da8eb461992fc430d92b918bc03494e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he00ec4c4e95e3566bc4b5950b601e6aad3360dc81158c3746a07b1e2b8014f6027549bc426c1694282b6de2081e99aec8677edebe0f61ab89350ff2073ab1026a7c0e3c634058536a6278d57d85ad50dda37e1dc7c0d1f6d8239231166b2efb824c0bad8189e82b9c206086c2ab16f264bf1345fe1f4e84a16e3be9ac42cf199;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40990adbe575c73baa3178f6b1690e1756238683b17d212de61b1df6e385f5c4e67d3f22069d097f69172420a980aa2e010dbfe2853c9003a8ac748c75edfc5df9f8ec8364c31def6a2a5fe831f359b8f82799f3ecabb9396b0eb0ec18b329dfdfc3431c092e99b42eb29251d5aab76df96894d5970bef8166864b8a2983acdd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79f48313c08894496ffeac32f40321559876ffb1dfeed6f2f7670ee7622125a97f6024bd896d30517db608f40b31718e3a1ef56d9511db6c8e096002fbfb1ba6023bd06b00445250cbf3cec845cbeda25f480a19ac54e3dd718659c17731afc8598ac1d5d96b986f313409ee20f9a7583cc218cc3b0c524fc755a1c45b507788;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1b46821358bbfb821427694f794d182d20e5f41c16a1afaaafb39e5a110705e555eb47be4e8b4b095464f95f3ba3aa468089ca575c31f994cd65fb7659baf6ddcdab14df72e63d8170365fcec3f09ad230064a0355588c41fc29759ee8c1f51fb72c789367c3dc4a079192f6dbcd23e6818bf09c51027253ec81ea197c281b9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2595ce18905b1a434e247bfa11f8f32a514dc8aa4966466560d1b315027594f2a50b660fe2e6eda4cd33f223766d843130c542b27835c8d184cd931b35698b220f1755df46e31143b2b47b4cd707b3cf402656608f56609e9b79c1d80ba2caa2b04a6ffd8a2cf2d8e9d180f606edff764bb60a70170cd570933e670a043bf6c3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70c1fa108d1238942233d4fb89c0caab4144191de891a193b3d609e99aa40c1312af64566897613dc28705b3da32724d4eff405f267e80b136b627f9837ac9acf7aa06997531370b113adaebeb8fde10efa08b6446231623ff3949395d68a93e8edde0350fc6c32791a42396ac8ac71034f4766b1aa7eae6088fd362a391b371;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h936aace73d40f3d7a8864b6c8c89c8dc06506551e89b7494bec1f0b42aed63b58863c7b03751afc5fa61c01cb6b3144c2ba2b03d7a4f72336756581ec5e91186cee25ce34e9aacea50bffac99b78811e16c8bbfda36921039b29642191f84e354c3e59915814bbb5403bb3ba3f6881a7cbaafcff30c183bfde052ca1b094fec1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha83841e817f88372f7c8a0d11d41e448abf7c05bc9253e02c5203164e079ac25510e0243d729e132fd0a8168cb08826893c8e89627ec08882519c8cdc28e1b6b27c474edb286eb0384eea80a06fd00d2ca4ddc73295bbd9eec52698e6df63c920928248bc7122de22bb35e4a85687ba2c802eaa1107986c3aa46cbdfaf1be59b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3660b7954f8698ac0474ab5248ace64f99d5b90544bc1b3dc2f16f1ef3454c73c8f530699112baaac1846be23c0a23b655f18a699a3e1a97783a81ee18c94d90d5ed50a0426f7f465516d735dc2fb4f44239e049e3ceaefb6a66fc85cb1f9262bda589bdf992657dad0ac82bd23fef727cd213ca6bae717c9dbf45ff9cf67c56;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd2942cf4835f597549ac16102999c83d3783170ab2f929a82dbf9460f3fb81af051649ba884f67a54a43bbaee27022199c480551b08c0ac63585a63908d7a101b45ad089373751cadf6d4cdbda115ea242b68ce78b30777e3e61aabf1ae26395eb49fcd61386d8822e9602dd0c2a5b5e6e8c06904de395391b47cdcf225d04;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h64ae43454319df7a7dd0138e4e461762109832b4d13d2d28988394f79c0fb5fb0b4f79785c43f2d356dfe534fdd8350e03b9eb1d883a092d68d91a367756b8abd864bc7112d05044e042187caa9c7afc0a9fa54d41ac9230fe13dfeb9a5aabbd24ebddc48c1bd261dcbaad0946ff09812a582a335165e8e4016d523be3be0be9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ffb9de4404bd1243ee26fd71c6937efd196f92f0b8118d422cadc4207244a51f02624c04e6387134f4842eeed0cdd9fc7e78f06ad2939374a714a6a6b1272836bb9e2e298f84338cbe480e8e8f97698d594fb490989ffc8dd72a38b7920626aa090ec5fab5f138e675d27eb56d8618d327ec5779fd34f32537a739dedd30083;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9fa80c0db492c5750b3ed4858cb412a73f1b1c6102530f8ed954ec5ff3270c21efa485145eb0bacbd1071b0ef4fbda138c1bddf7f7bddfc8ffb37f1cfc2f6656f3481adf61323c1678192896e2743ce5a618271094d74ee7f502ebe13d3982a05ffaf9d167912bb8b925b61baae560c35b58da2b007580b42f0b9c4f7286804;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6424151715b27afa3bc5e1dd9462b403d1e665c9af0746cddf994d0a17f67278f0bde1b543fe708652e93d62a52fb4d412d2c6200e027868056f23a7ff313e24d4c6ae966d3cb00030d6ece3b70205665b3258bf865c3c6c015d4466ea5bb6b24b19e4a90ed8d644acbfdf324ec55789decc6828ee2cf2e280cc220de1a0925;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf71bdcf5e2125c7a9da6168f541be81f976152c4e3bf569ab7eb382331bdbca02361f8b4f4c580360cf03ea22d82ac3170bf819312b9f8211e6f99d126d1a13511127c723ea6f74c72c69f14aa5bc50a94220e0aa667f205540d96a17c51896e2d2df7dcdafd4baaee7883c4bc6c6be36340bce818235fcf83377ba91fbab136;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8eb423b673b50b2403f3307617f16309d30da81633ff172586e6689169f6d56e5c77189b217cd7aeb8ef26a6d58eeb3193102a7e24b9606f27cd1741de4e1c451876613a588e66fa3374945e2517085ba598bf5a68ac5e5d053b728a3e505e59a81a355641365c664c4be7802b22aa7aae6377d6ef76cfa49ff48668c29fdd08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h678d4143cc729c165090709235665c922708f43b07d20471391448cc9fcecc59422bfa775ec6800e0743268be75f684428fcc737163e7eb82714365e4cb2008031f602e0366002db2a55d02c55147fd45c35fb2f22402a092e374d85bea625351e5108e030c9f4dc4e02b67d6ec11486d5500ca8c1232b7853b09006f2d70265;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h130326dda4c02262cfde853054d7c6bdfa2c45f5f70dc12e4a0da0000d1f65cb50265965804b3ee90071b764d443923ca11c5b905ccfaa4c48f99826d3e861d18cf086370304816523bd762546293211ece8f3e24a9c17d3513c20ff027a35260c36374078078dd7e88223cd2c9b592cbf378f59716f95f53089ac68f120113c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b8e501eb01b9268b8fad24e311d349294b4d525822f1b01f6d766577f6b4883965a9de542007ce0257ecf63204d48f9515f8010a10ae1eb66f844aaba87b7f74c4ab92b8a647114a661a57edf4530a8a58aae8a8baa183211da7597dfe501d3d391c2323b404a0d6ea50d7be9f675ed582c215a04ef59b2ba9d0cc9bf5cae4d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haad02e2759225c9673d9637499d13eb071ab301856936e0aa450c04e00d78a84735c265e521186a1a5a69eca44dc1eae03735d949c5d7f885c947a89e710648252aa984d04e78c6fbc3f0298567cb561bac7d0d615e3cf18b0a7e019f2797937c3168431725c9874336512e1e8e1ff58198edee08bf7e9e95efad07777bdf75a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15593d67d528dc0f939302725280ffbbf48dca63a464293cc91d08b9d6084a93ebba2539161854228a02468b8b4bbd4d1ad4c4d478555200af08d76edd8d8aff64c8ae4e4efdcb98961a87d5371ce26f3b0d408a3b08341af973b6ab7ac287b852d29f6333f97e0da1b93c9c62bc37d681133b195005ffbdef30f8660ea643bf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32c364c935a4e1578fee2096df637e99220295fdfc66d841dbc444b6f98cf33014ea9c2949bec499b4c825f9753ec46a115f9af7f324b65435eca7dbaf5e402db134c9970aeb53771d8288d53af60a1ac3e8c4200b69bb1ee163e16524387f5f370ed87a188862954b509f5ac0bc5cc4979ad9fa462b3404ba41b40c6eb7b32e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35a5937f75152c8902af9960e5286d8059503d867b4ca7c54de9e9ab53a378c2fa5b1f9f58eb845402a47cebdb34266259b86c853d0f5fceea3cc60563aefe9d47a51915bc619ea33ac0b22361fc7bfa520497378894220a3f706e9ad8bd91d6b4ea3a4aa40c96eed77b49c591b2071a1ce149947b623817302bf93835b96b00;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb5a03ceca57226e2b232675d0e21c159a808d34281075d612df2a77d7b7b2b933f5acb8537b323c7572fee9044aadf78dd6e4e3cf615232bcf17c47fe678696bed30da78c0794f76232054f93b13e35ad1d046a6f888c357cec059b3410e8f1f827eb1bc2cfa1445a2770c08778225ceda85f8f7cde2fcc52f550c68d55a76d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc32c73d625c466c6c766a11f89fcd9ff6346e6bd3962a9a9553d859b3223b161e872b762b1e028245f144f22ff80a7e2398fd2b2de1922014661c414d61c44f925ed27496e33dca6158c110b915eff89f9306a73e60c0756855bb779a35113eb0c1c5db9aa53cc6e711921e8bc134e28939559f4ed8cca29649bc97d49ddc0c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd83ab77933a61d50ef84ca4463592b808361d8adb3dc6d85dd4e7550ea782b092016dd0db6c90f296e53ae4b32c04435fff779d886156a130391ce3a394a9beabcff065f0d1d643086db7c37bba13028954c8a60b2468be71dd1c54b6028059a9a1676552404ac7c098a54a755870233acb43cedc3008d16e7f175d6bd0cef56;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5bd2f227e5c13271d542db959cd7511442184f4525194c06a33e460f593a2d6b8c21e8b26a671f2a214540faf9b5f1ce6e1b05f47740dfa7ec0e9353b219410257a641965412dc13363801ce520401cd0f0eab4562902ee8f6dab2e99aa8dbc35da956d17ce534a8cccac524aebcde16d18bd3abf78dcb5bdd5df1107f2f7df;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6642e2574a0eedad57c9e0b735bd7132bd6f8e66a4172357f9c807625f5caba0125149e4cddde3b76f0e487f18d16593d4428e4a8a6f5a0a3789caf6aeb22a979bdc436e727dc32d6393cb6fec25fc0b9b89497651681c6a394123639ced48e33276f7a6fba5a1e78a9464ce5d2cf47b07aca0dd6d72682296bb514efa27877a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a8929c28d979720592f314b01b5d9b64664c5f6d1a3321b71efae4b0e45070d05e40c0f1261ce2eadad3caada78f5d50df3d1e05d3418413a57b967d472c36ce3027f661257a6c38d205e2e93c7270af1028120f8fd64c8e1ecf66680d0c0ed95c352be356358e1ae8cae25771144fa31fdfe27104095e7e119c59b6ca87f62;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e7eeba6e2546227ffa3199191c638305ec18d702720a7cfcf785971ad56decc4fb907a5a61d11aa418ef0f269e5e1017b46f95e811e633a228509e837c6218923b9df9fab68247d43d316ece40e7a6d20d45fe9fe711cb5372f51a572550e9a0b6ce86a9b2371423274c2bf3464141d4863170c04ecf7173ce1c9acdab17c19;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a0b2b63d137f78ae8aa36de0a94016cadd47eb8a89d0574c6ad3bc2867f3984037ac6feea0bfba12ba409f86c91835fa385d6731d42383f5c665614322388b16850a4d7d0d310a790823e869bce77c259331bd6d3fd7bd3efc11d9e903d32c217adbbc431587f98abb84582dd31d91b750879a342003cb4cd2b249af52aa23d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h456e934b1b7c0879eb87480bd6fc6e7e605abd51eee3afef854fc53d982552ef5ade693a2600cf96fc80f01005fd8a429b32e21e2c6dca53b5399e468d614aa389b7310bd59024e38208ef5f67b79b0198e419c5aa298dfe5716c1ba1ed1031ffe8a3cf7a28f29200ad3690241f4f1b49fc472db4912a82f0d8e5045788feef8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72d96eb0b722edb4bde87c62b69a111161e113d1d4b46ecc4f01b438768f5296bdb64380ba3c7f6fec25c1a2c7223cec5ae690423707a860abd95eaaddf3c8863325e5b0866ba09332eee46714951fa933152567b64378d62774e2b54de7c84cb83595557d7c5331e6ce157c44b6223675697296b180a20034e75ba279f56ef0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b406094d520004dfb0b35808ecc8ac66aa30e0abfbba704df2d59a744d60742b7254d8692623be044054a1947d97eb64759ec649f62e890043aed27e78bfb3ed9c21410470ab7c8020be9b5b650b55f99efd8a39dbcc46ddd0610aee29f9e9713c2408284718775649263531a8269c50da5f656eaf1bcfaf560f75a1b0513c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4614ec45e815b328dd3bb36c3adb34e2d46463ac455bf17bbc6178400c83bb6737d6f8071e140e5266f266eda63caaf5314cbb50f7eb058a901f4d64552b28491d40e4e768ab176492c3612a69d8726e040f26062c282d3e0c8c4332ab9c1c8b29695dc99ad10870a0952c045219049b46379dfb4de684a733e84035944654b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5c8c4255ab778ab6e40ee5b0c77777e791bf4c26a5a339b4619236f300d70ecb65b7cae4e1534de02d4200e0b1730337ae5c1d226b9a78e8e6f2f329b7216918d351753e84bc9bcd82f2feda47c39cc01f8727d46c04a6d7dbf1dfbbfa93b27680370268605befb892b1e243cbfedcf730c0e1318dadf3653cf20142a37304;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h31742bf8e81fba5c480fb2aa3d73cb5f5889010b34a532448aee889c05bb01a1c2735982592e4dc97a9b7f283f98e38a94a48810f8a16725f24dd8fdaf9c757702dd1b7f7e7948a5b43ff6185875108b78cc65608270ead4d853fce36d85bd0e33f0bf53775e9a232acd38e174e5e6678ab1247018b0b817e605fff735b27053;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3d3d91009d6923d35dd06a1d636477fe216aa8fc6d8838ec46bdb8b4248b5e06c5460de21890466ef32ab1300916578aec6c728c11df779fac4e0e5c27f1b1e4640a0f2cba5d69d64d39892e8be67a611c8a98f7d3b68a69652a4505d09cbb9b4a09b9a63944c4858a1e58a9494f9436cefdb64af5b0e52d0f054808b5735d9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h444a6f5b4a01aa11d4f66a26319e7156c827447b6b8df558eaaebc1f52a24eadc3a21287140cb6e61db42b8e3dbc26e220406729808c61888ff7b16cf04d0b09dd5ac961eff98718c397e45a5b1095a280031781ec90a5d9b743cb953d1887e04db6041795f0626343d3a1a7f57ecc0abc7cbd0a7f0a8fd8cb9f6697dcb8221b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h100e3fd063e0ffdfb8f4df1191fad1181b38578a73b3ca3c536922b9b1fc2b624c985135bf78f18793275d4357fd723be78bc4f95615e8400d9d97534676c6bc025347018fa94332624ba94396a057a0f8c17679d8c0ed370fc6a82ebb13c04ce2a5e9199e2222912b30c35671bab9d900751a78c2991252bc90a4c055ef4051;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7429e1b4f87b23893a1d56b06079a5b431e3c8b0f4d3ae990ac54c6241adb090770185adce537328723d6269ebd347dd42c029515bccfcd0041f6c666db16456c4675cbe2e82adf5d8f6e7ae540d15f1af0bf4f1c0c7bcbbaf2c373507b7c004051328e394232dd563c6f38270f2723cfeb6fa5c99de206e3ee5359d4174d19;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f0dd1a9323c94751ca660351031d60655062072b4d167c5d2890f1f1b107b88dca0953f58bf19a91ada1a30f04ed6eda4b76d47708a4619ff47d8faea8740584655d7cf7c6662e4b15874134539382e0e39ad49efa8595cd8ce41afae5a6992efc85430c0d9f52be613435a6cdcf789fefad44eace65d0b02fdb63ca13cf5ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ef5e9ae1a337b452d17ce68b19c6415649701f32fdc0699e5269765b2faa5d965f2fe3c5c14096cb0dd4326c9c92c373ed414c9b5df87d99d8ce8544488b0f76e9df126f4a73bc8686fbd8a5161da74ff475423be3b8e0787aa51e8dbbf8607ee9c2621add77b4a52d4c1f7eb189d01d1154dc9e46b0c3d306f8a0aee47c0df;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8b5247a94380c399121f1ea0df9a236812f510f3220bef9f7570c6e1c742c20c31cd820c5d238f1f01a53e1a399be10824b8c03768c0bea0fbbd5ae43f7c131c773ff0151dd40801749d9f0ba9df71f56a04388f25aaba02b8f60d4801fd4d98c8d4e84cc79b2e9ebaa6a1f4ab2e03649a8f35ce80a5a9bb73a1de8956f7be2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3ee5932127789c715ba5c8cff5b67208dc84b15aa16c6741eabc3d47b3958b621fd4be4f64bc66f14745ef11a392886797cfd83946881b216a2eed370c915feb8fe7c80768c0647033cc1c5dcf4934c22b2ac8c24e47fa1056e819dbf17311e088fa8d86e99c6a30e0199b9cc7a160277cf026190d551aa9a3ad88a4efc92;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha72577c7786491188c1dbbdd1ad0c263db7fd67c1a28633a7930892d4dae26e2c372a50dc356f922c3d507d6cb15d3c30ef15ea1e008cdc943664f605bd13b285c33643f6145df84ba2f8f63c2ae8e420623562e99f16e9ab75f4c834378eb072766a205cf05f566a1a449146019aaa04bb6fc894b54596da1fd1db244cdcece;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4ec25e9f04eb95231a29dff86fe7e08ec65688152e0012f54a057168251222e62e5640ff406f7a52922c0fdb6c78b8d99f0e94ef1e761b4b4866c08831b2d966c422d766671edb84e1a8e87a112873d2f8a18c0c881a0e7e1e8c96cae43b93d20d2ad4d0c02770b7f7e59a1b21f49779553e8067522fb43589c28e1c07a7e5a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95da61805c2fcd5af672ba47714d2a4330d3aaa4047ff12b4892460b8ff4e697679c63d046571407f85aec929abc2acff3003db5b0e1fb3631256cd75ce0cb8829927c4f4f935e871f62765ab59c04b68238637092387f34e84456a6c3abe583b602946c3a4e78556ac42e35a7ec00e33ba0129f30d115c060142fdd73c18f8c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8cca9c578013131f4035bcc1d3cede8536a2863503410ede23b1f876d4e7136ecaee4ba79e8b2bf64590879a6249ac8e7d63eb6a08fb842b16bb021ba59aff298988fb244a8bcebed5531a3ec9afed8012624a22109f60ea7ec6580286f7a93f7ef7ffa870c0aeaaa57757e2bc6f42f4cef2b1fcc7a1570846d968895699e8f7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86ba132540a61916b67dc53e411ed5b96580ef6eb73f608162b6ff91fa529af10ec7d43ea9fd7aeb30093e5b2aa7fed5b429ea26df54ba8098f5d4546a440c7f85874c50857c9b7a63c3420cfe2309ccdd11bbed2a6b7360a9049642651e67da5ff015f88c08d35825a857152ca851cc637939683c2c016fa2aed30935acc742;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbc3d8d88ea015f43baede8ab1da5cca753ebbae3f5adafc2c94cb74a43203deef2a2bd51ea7beb02d43425214d5b144bed57aa2c534cc6a1acc30d13c22714c7daf6a69386abc104859982dd4a195e953065bc5d2281b81711fdcd52e69354c8de24bcec6daaf7577b74a5927308010fa7f9a4d91f4365567a74aea609843f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26d18f62a58c939edc5e307caa31d3e1d19b7529647eaa65b473df6459a8ddac9c685059adc87f8c65c6ac7ad92a67d9e334648f3cd2b7b91405490a308a76b3323265113ae267f2b134dbe3af1aba335cc27a8a92f79530d48affcba2dcde5938af59e16778a0625dc365062d1f0c3172827135e46eb070db67ad9e9eb6bf47;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19e4559582813a464706631005c9a0531f114b684e192fc2629594b2a1465476d3aa4df279568c560c2be688709c69feb1afca1198879bae6361f3e291bd0dba1cccb3025e95f2e83bee1ea538f393f837ff63e7eb2b8e9888e27117555b0dfaa5bf85ee385019928d5d55a8e375a2332a9d47304f2dce27d7dc9dbe7560d9c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46d0726db553dc73db9aa7f0267c103ae37f9e24fa7f6900ff70c8228a012bf34b824ad2b2eea3da12111c042038abe6235aaf115640be94567641759a4d890aa99bd73774829a39f24cf61af90aa45094c0f1dbd313cbc581d0278ec2bec7794e3ea42c021d605b5f832811c54e2f48dee9febb262b110968fc0bd2f11df3d9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9946747f0d2936ada1d0b2a15132ff580e3c6086955c92e0e3bd2c22e91b695dee39627cf9a9e079e9d6ebd92d94b0bc14b2c43ae0a994bb9957e79528f4960197977ad1426fdb5f06d6c8eb7d19123016da0a5425eee515401ae7a089fb7d1bb8546096dbbb5c471364644de21d018a51ab41b2e2c2952c7c81844d3f5acd49;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10c53a4eded724c0c52bb790fa1709d05adc2a8a44c7d297ca1162f7657ab5dee09590c801cd03381fa3f4c4501272554322df71ae823adc42af1edaaa2458a86b9f94adf51b6be6cb6885f1ebf0d98b0f149876b5e626c1fde22e47135a15ff678a574825a06bb71b8a54d0da81dae8ec054691559ee4a9e4a37e64ff1db035;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee44cabbfd62bd537a8fceba12b625ffe71010247bb6d983b8804c183c9046d280cc6ee248f32e1a8d82d114b36c25449d9bb57564d5fe1db5640fa4716716834952cdc531f58ac94f52b18859b4bcf6bddd7053b34784f6d1ce8090315b935d8fbd3b174ceab7ee40b7d7681a59705fb2e7979d7b689ee0092cfa68f6d72122;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34c29d9ed8a8f15dea63aeb13d3fc6353a4ea799719fa6784527b79adb54e8fbb4c217715b0dd8718c65386ba99826a599117f8c401682a60535d1c9adde703f41b1613dca2017a32b5ac1be3e577e122e25761694092f94e51230e9ca0cf15f800fe7579eef0f08660029a54f12ddffc9b688d919e5593f4324b97d289b2c7b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6327b1c0eac88576995d666aba0062172885eac3a736059bff068d302ec49daac1df27cd88dfce3106abe8304ecd2ffe52e112c1321247a3ee5adb8141e57aff1626efce2abee13c10ba70504a7fe3a89b6bd7e3f41b91c3f8903c3735c0b087917637251c6a02c300bc267e12c2ece48fa5c0317a3e94a6391624db804eda96;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c376926b21a7d74a54b7b12c0abece692640c15b34dc00ee70fb5f240f17d793a96dc83cc02bc8ffc6fc4568c05f9fa20242988ba5f41dd4ffe230f3c1976e8f5e7377cc7fca8c9bc2850ba0c27c9218bf65cdad114d62195564b7ff87f3500c60916ae4a94270ce6af7b23e14256f7b7b9c0d5b90483d6e8766931579b7b6c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71541d312f00caad949e637ccfbb8fcd33476f838986c89898361c5e644a9f0581d7246b8dbfaf61aa7002af2a8f060a3e98b8fe5db058c285d4ed494a8bc35e956161a30c103345ef5ee050de3f55a73c9c3257240b556fa7c59a75e99286f901fe966a79dd1461446479be883e72fb15a5c35dd4cd201108ce090b1dc7e2b6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc087ad023f92ce56b70073e0767d7d769af67cf93b7659c40782c1eaed9d0aa3c0c102989d696629bd7f758250da3b3fd4f6757e5fb604cd8ae4bb30b60a221f9970a756bba0a95e90473091296e185fb713e5938c2ca160940fb3e6a22eb978fd8a767015991d2457915ff8402e66983e336f7143db27293ba242bac1015d7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h247d56139d28b116e69d1380b3f66c3a1602325807517be5ae4a71d4131d107444743cd7a61a20515ce00d614fa3424a1e1b8b9f17b41a0cd28461e961211136b9ef24371c4083239eb0aa438fcb44fd847c0c97e634eb8abe69e5bccbc8a5854449549f39ccea0445d89b31fce9a8adc607a81fd90eae649c8c2890a7475b66;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf575b7bef6da5b3f0a1776bc15185f8869fc16a10a10df03a2ae71af54c46ba48ca722cb997bf3ff2a1768f44638f289ddd6e701af5ae95a70287be0d3fde947b22d393a4e07e53f2d4f869f20353d89bb55697ca436df203edd3b1ff622a1b5ad1b4317b0d49492fab8e433b6805859dcbad8ae527476fc5185b8cf485a097;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h271f1f74928fbe51435504d7ffc3e6cc766b0d814e465cd60b38fe7c7601b42685e14e936f6b71683398abf0887f822843aa2b2abf308ce398b9c711bb4ce1086b1a52383e26a7ec9857b4319c5d07c4a6b0da6a65e468f9676e809364bda4914be7e6c65163c94aad5920b148ee37e9659ad1b07afb17ff059a5ff52ae628e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5a631ed52c82f2cf0ee7bd3b927a9e22a8f014bff73ebad595cebcecfe2a0434724f76edb8e606b98ddcdd843ba536c46c969c4f4824564ed072dfdb6b1de564cae9f178a84aaa9d4297831fcf9bbe1194ada452a30696073377da48586907c15c0d4456b73be6fb5f0d734c872645905467ed6abc51c6c8a25626df3f188fe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3013baf1229c037ce269f8e9aa236be7868230a5a6d42161b923f5665e182e9cec2773d5d33bd76ba353dde9f743a39f75aa1b1dc4a4b981139841fb1bb042cee255c6fcc6db880afab0dc0ccc5507298f4e8d50e7368bb032071d9caef51941fac64e6307fa2db61e9e9bc739ba098442eb9d409860a55f301efd7ab5d2720;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53a5c77621b1b2acb3c74fb3676774ade9871881e4c96c8ee467fc35f78dff3d7d7ba1b19b6abca2036f2f1213e821d3f19c26dffbbee09ac6e397386d3d3f84a236859f83296d873f2debb803f5328ff08b1b4e8727cc3b0f322130fd347747f2e00ec65f3b8b766009bc643dae54bb910cde07c657025912d437fba14f0cd4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c5af0741817614c45a940118d3118cabb4a4ea615632e98d216af2a73683fbe5170247b9d17618545e63472a49ed908b3547b92c7f0496b028d4d4e6bc3d5e02d03f40345a8587866c92889de44b39d7b7a16247830bc3015eae4eacbbb9fb2ad10104276529f36299ed8ce33eb89b3598bfd1f85ff8567aba6a84bc6a2f189;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'habdca6c22b9ac366805fee38b844fd2300267ca44f7212425657833418930ff7bc99b092a5e09c2c21c2286e93a0584f5dc763c5433e72de82485c0723678d607369ca44b23647639cc2a56a15eb2cf1a3c1ee647bc092444df9d4cc1ce18d74879ef261d49cf7c23ebf7348919faeb1a989069344c27c8599a72405cdc3a5cb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d8a7bfef7032cd648138fe268decfeb4b8c75b84f5152bf796cf047438f8b5540122f5c0b0a819c8860a20cb09b81353d6856e855fe788468f4a5b91b0259c6c1f095b81574977b7d2bec012f3b6e8f3dc6e680403fb902e6a5fa65cf2f94e2909297949036db94cfb9e192c09b7b17fe408d1bc63d2ed21bd450b2b7701726;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha64e9ad31847cd2f8307968a7e6d54d18399902ac7a9d71051f1e60c08e14ab25ebd63ca5ee0c8bf5196f0671b405be7c1a7b96e109a50006bb11cfaef41fc49449c4a5724900e5b9ae1f9cdb5fa5818941c9ccb87a0f251510d52cea9eca652259dc8192086be4eba71251b5332e34cb3a8a47e8a7fef2e59a3ea02cc5ea0b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a066ea8198ef9da2759302c0f223b71e008a9f287eea2a3e2c45fac246301b6a6db8900b4e175495ae2feee99662a9f537d829de060f05b3d8a40a69e4801dbc8b108ec938065920c152fe6c76dcb71544f6c3f886d211114b259f5b6caa55d025f0583eefe821c41939ac3f07bf8811b3d480e5a226e0185d87fb81017b6a1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d8eff7874bfa31c27b422f7a5555d734a41473f70b1ed1e9b32a0e8d94f6cb1e4fbe517f2b5410ea8c7586855f65a98aff3f2443bdda494e89846d29e1a9ed0516bc0b74e49b7d19d9741d9b5b07ab19df996e2a81d92f6a5b64e5c1dc14c513f0f67b9b695c9304104ccb61ff4cb64b17a6cdd1ef0829d3e6dfcf219b1b777;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b889435b0a8d8bf1ce25ed8c4aba1bb60252cd04dd629b24b72fb5fa333c218af7037dd76de78675d2bb7e34cbae6f7aa37b1dd8c24b09ee43fcb06048aa1ced5c0d1979ae49f81261747858bb1d658fbfe7c70f930544139f4c4534027348f1b9a62008a72a9e55b184cefe6ed06cd0a8b140329c1161601bed7db16b99447;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha023717a8d17892ee27852be6b916b71f0666372a00a7abd638e7aed2571baf08cf54f3932fb599e717c41ce9ec9ff480e18d9a3e711bfb8e7df7d9660c480ff714e2baa33253ce16723251b98c3504dd3de9060ed7feb60944fc3ad0ec3fbfc2192efca00c39e85a13e692b622378e0ea923a6aa91c98345d59f0d55ec3c94d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c8546c416e8e99aa15de5102af0d6fe5e16647bf30d81e5c763db6ebb41ffb92ddccdc4929d930f5bebddfaa6d43b47a6f397624f2da5e2d49849b15eacc902e257994ea75d809d654782dabb960940edbf51e0fccbf88c4c08b99b8fee8a3b49fb055e0999db0ad1b93e8c6b460fdf041be75c746f9d1921a1657a8542d363;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7c61b6be71d672944fdc2dcdc43fa2164be6b00a5b695ad9116ad90e0e9577f62e15ccd4f041563075970c5d2d5ea4610fb677bfb96b4f55a530518313dd5f29e1ded5f060bc7a4b40b4d182ae5f1ad703f523bab452cf55899e5f63521ce32dcde39ca4faec3e3db5e35ea93229238645e2491090a7f545096e31780612c0e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h375068098ee3b9dc5c702747a83f72bbc495ac293b344af298b9d5c5fe9416c2f05473c42d0aacd01730df0b15cc85962b1c9a4fe01954a46ad8a337b6aca94be2db232bd1b1a1d62305f2dda087844d0690048e66d71bc97987c259f925af9612a243c15c07f52326bf0130b4b53ff0e540934f67bc773de9eaf49b56c0ce37;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h796bae9b81718c24b33de4cf0c14f3e535c50c620833ebeef7cb276670dcddbe2af2b13f051fa36bb97bc2be5214e165a41e14b71b98fa0a96849047046124c0c8693e1baa48e2375dba45e712dda1af952aff51f88f7a014f7c016beb5631203bcd568a6455562d00f7a67ee6d1325e6e78f9674c11cd53f5e269b8d2c826f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1dc3389d4b1fc974983b7b22cdb1308a0a21105be4f4e25242a8bae1f5d023fb53fa9b4f250bd0f737237808ae0045a9536bcaea118d05dde01f4c98b01f0dee50243dd25b324c1484b876a4a492bf52be74159ed7b9bbe7e942bf2ae8afb95e3902af636939094aa50db866ad2fd09c619e2c7619c02d4363b20cdb7fc8950a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a17f3e4f62f20f9e29c739472628af7dbe83b257e7d3ded179366a43055cce2922372ea107f67751dc9d87ed7ff1da737065bcccaffeb915b6684a8ab1cb3970e9b69903ad07e03dba5e83a495b8c4c6b32a19d497039398332c5071e64b14076aee04547ca445cbc30840970b9c19bc36e391fff3d3c2235184244bedb882a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h456b2c9408557502af6ecdc71542a838cb4cdaecd8a2d3465134a5af18ee928720a31b081f344f5184dae6dc2c82e22d4e61a740e7c9d888a42d2bd81405ab48ec3ee766534674787ef8aa321bef3e2460f5bd5a23ed8ddd1a038ed5d1cd9a0c5301e424864c37a9a20e982cbe58d8c3a511b0979f1729529d312a873784dd07;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70a0bb765197b473d496e9f4df485af6ffa149f59d01419f4cb5ad9bf3408fa381f36dc75d51b6900cddcdb2158b59f0619ad44ea39846c5d99906c88ce005ebb076788094f6564eaa67df8ebe5e3bd10633be75b9f815908e050bbc7b13761b1b2f4be388c63a16cc7064e60541d7533963a430d8713831f828bae057a42810;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6830bae57b1aa0c71967447d278e79e279356ab7c2a08eeefbc82ded326c5c573b4213de0f3ba05040be44c7b52a719536ae056c3b67aca03cf567865073ca74e5dea9e03d0e49ce9aec9029624b3b30ca46db6a49f69c4a386e1660a0345cc3de73daefeaafd8a5bf9061fa6a4cdf42f2cd112cef8b98a2f8efe42ace7e71;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf74e33352edd16dd244aaf78c464a7b97777ec06c0b442cde27aa5843a68895d52b89536f9040de479b3a34b7400a32ab903579b41b811e5754d64a6c50feb1a7b3d98ce87a7e8241620defe6dc3de63b256d18087a11786b0621cd3ee5777a01113e3b92cb89fabb388008f83ff7c066ccf67a604d788826ca499f55ae3976c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9db48702ab97991644d3af46f5ed2b45db8bd926a59a7da9b46570bbad8f39bb2a7521570c2defb37a7cc09e09cd118d1ac5eccac6ff83b71596e7feec36632c54326f3bedc5585d103f3c416fc151d2c5f5f5e02cb163457a64b768cb744fbd7acdb04bd5e6b1051f3edf43fd19a394ef4b01f42ac4ef821f9c4e6b3ed01a2c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f5f849d8b9f9a8d76f5457c31ebaddfe2227b52a9721cbd3327b4602a5838236da0a8eb99482eed802e5a5e5ea8b7727c86cde093347b91a1353a8166bfb6840b6e0e116262e2fa5309ccaacffe61fb7276996c870ab82229be4bf5c71b9d0a5224d42381c444c47ada6e2a18ffd3ddbae779affba94ec953422ff464db7d04;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3bb85db248fd8a831550486808d112164fe5ab01d87075cea69414b6aa5dcf607322be2c88bce65b6a56fe5a00206fc3df976342bfca66e7606a331fae30f3b614bae96a6ac89cf6fb6d81242f253b119be0f81d26374023a37e39fd9f16c13e6021cad1b28e5e56a8b69b14ff63a249f3f9539be20bf3cbdb8b650c667601b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51698da290367baa8413b0184158fc659a33d33de7a213cc3b028d08bb67040b13a8543cc4b771a3b7fc64b75faf4ba5de91af88e9c652683c874552a6df9b1145ed96a4076b1fd0303cfd8dae4d4163304faf902090e466515eee8cf602def227c2de73d7ee61595378bf65658fc8741d098ab4271b4ea94c9ca48b42cd4905;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9e2140991fdcadbd0015ed146b39cc03af60907a6d196aeb5f53ce5552bc61863b9081bbf9741f448764b1411b01e2bfc693f288f30170feef9ef6d24d929c28b132f0a15b0ff27973a427a27806b2a69637b409be83c4ac81ac48efdbda6e62651a58daa3e0ad4c9ff51c032ba3a070ab0c571d5c01292c9f17622bb238df9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49f77ffe3af4982cc871672667af9fa620d9ebe479f3a582aa999fb2b12c30c5863c2f5ee009e4f91f20889fa57d5e6ba956bcfecc3765abba5267479ec10815b703e7d924ce9e64e56eaf4c31f57cfec38a50d31cd90818ea3fc0a1f09948eee42499649f2e3cc3fe063c9ac11354ee83d4343292c5531c141c1f5d5976a9ec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'habe1dc8a501e01c61296712cb1c569b98d2006f4a373a781a0fcc4b481c55689c311f7ed739d5ec32e7f7a332d75b9a5b7fd030296891cee3944c8d65fb3ca7c44378fde3bf00e957b26c552d0c09bcfea774ce1e36650ed097605ff63a3f503cdbd6a836dce1d093a4b41ee0cbae335e844e46c44ef3928514a4bd77826f180;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3dbdf4b20bf1a692887f8d721bbaa38355cc629c8024a7d7d1f572781d9a5598bbb9fe69e1f41ec6f9247096f9069cd6f9058954fb385b3a185dfbefe88c5ea1ee9bd8277528c9d42ee38da64039fab59696499e351a36e09ea35354ef00f2bc75f7956608b6557989145737d1dcd93bd8698714eaaf3c445b4679fd7a3bfb7f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4cbb87e8abf8b342b2dbebe025157ec4dd2685a41be5f4e7ae79450690966f6927dae1d0150d3fff8ebafe6499bd71c44ec8e4d9b35822906cabd957540a44941d50c2f154f1ab8f541cc6b3d9f9c3ef2be4b770a2a16aae336678ecbd49fd6379e91714e1ae9f4dcee906f17f64965177d8fe444ca5e0e242752efe3342361f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h361d4ccfdaacded7177350a58e4383aef07fa26c928b06f3d432c79de750d2acc6b64a15840939c250e1bdad9bb926587c7ab38dcdbf82b9bf98053e3f256ed1c0ef964716493ec82207211e0352bf9ef0e0f4f1cae044508124bf2e01e85795119f55ee3d6de9def9eba7a71eed8bbea55abf97d9f8140a2dbfe2de5df691f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc394a6d744d4e0b1281ad8bf34b64edd67d130b3de3a0e0692cc8dc8b9c7b287de4e1a77c59ec6b96de4a90f67c36e39e38824a5faa7440c0377ed4715d0c88476f7fa3f2f474abfd52d7ab069a4805a537d0eb93d2dc6480fb6a3dadf52ecbd00d322a999d64c9a91594b265494fdc7cf88fc1d535e28d275f9066445713619;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd3e8a07078756ee6afa853ba1f8aa92a0c0c96c94d86ea98e7ba682506c221651b4a8c2cdfee3540df05fc5626a96df2c25af0674e4073e1616ba4ae9218e4adc042b71174c656c643c8ae730652a1a9c681a364174cdd325dfee7bd19ef658e5ec64822b88a364f28f546bce707522c4f4b70315be0fc7d6e740da8d283e8c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78f5e71a97a9e1f7cce56b36331c869cd1f694705799e455b78ef606b397e6c2cc78ece4daced7d1e6db5dbdc5e9914a9af1b987c41f1922652be96c63abc82adc1e0cc312f38f481bebd3af1ae349090e2d1ddf53a3b381d1ff8c714908dbb3e4072df5a3f45943183df9ab681d584090398e546eb3bdcd6844ef0e658a3fca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h189aa37a2b99f13f351365e89017d47216c198cdd0c34d30a837655fab1c421c14f6ea59de9c8cdf59396a47a8f6c0d14b8bf119d963f5ae607ebce7a7268f457798e50edac8fed9f9a71f137808b5db1297574354eb36b6823b395fd81a35edb0b0f50fc0251ec476f9829cd713b062f0e62ddf4985a3cf009d91bf8dca2741;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he01b66a8b02c76d84ee477d136bd3ee8c40f9af70a222cb2c111277b4650f8baf2b2e915c9c9d2a9a6db5ff65b5387cce08be625b95d63ab9c6231ecfa350e8d295d4f9376e69a422deab36e5930a5bcb9e9fe4d6d7bd804f0779d8f609cbbf782f23e889815d28e0335ef8595c451dffda07e742148fae9d4c306e2f16f96e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha05e66d95bb40a090239a2d7443c029e9e6983f326853adffc70fb94fc364f5da3b8f7f1fc5dc6162ca9b9f36f2e1c85041ea629dce4f10b12677a46b8c6b8518be069cd0428967fe83cdf9fcc03eaf008cb54a8d15d0efd5cb4fc1cdf8665565a09f18117c0fb00cac031779ea14c8f901896adf91abbaebbee393bc9e6ec9c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd95aa9e38f67f96caf60db766b9c9f98fc25e009bc7542ea45bcf5464d0fc406130b06dd94c1d385291c6d3949ce5c9bbd5517f499259bf1506c9ae34fc6639f8bb546dac0ec6b13b957de8bc2ea3ee79e335c8cac91778f58976653bba08c66cf0caadc51b20c19e65fb15c2bb2a2a112fa8effad749bfc33a551db0fca64a1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a83264a7352f3d817557cea36021277727b0ad270ebd1386f97ed071084a65ef5e46dceac98d595e3da7c3064b4971bdb166f4f688ee02b0b3ab155a9b51fa4cb57e6bc95700af39c6217c2ac51505ad1efe3c30d1c7a7f978bfd8c1b91893c1de9ec000861c5441f8fdc252e616daf5ed16034176383672e89daa0a215167c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce8dded8c80d85261f5fc9c13dfbe3111349d6da9cef0487762c6bbb78ae62e5ee3bc7e62c773934225d6dfaad664d553ad69eae59ef90c74c722672ddf0bf1fa124652203fbeb2bf5d0c8d04a25d3db15a9ab4ec27b69668bf6d57887746fd45a7240aa0414793c016930cda20305f5cef8fbb4a0d39bdd5a337a081f85af81;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h33a04b2d41a7a541a03f4057800fd44f97f97cae923d6edf42fbde2cfa7693507e3046bf009760922b4a366861a349bd40d8c464b6d339bf7b75d4450f284f20a1d78b1ae76cd074754194b3607bb7b6ed2113eecbd6ef50e9dfea96c6cb292759893d75ce22c87daa70a432b55bcd2b5c2ea0c9b955948ff77207c38861f8e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1af9e860e05f80d4eababe48ed96ad47409d0e920df6a03a5aaec6fc12f6413af4c5a9bc760e128c14beb9e093cb38c627129cd94833430521a0f10eeec44aa6b837abd45a3762b898f735d83eb37e588ba819a42e69091a4b896d468164fbcb42fc90fd992844e3f57163d717d65f238c49452b34e74bc39c9d51bd58f074fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c7de8d898a8f5dd438781cb9b009d0bedf0cd664353e888d5761c91f38e9d08f6c4daf1466868261831138001cc1b9b0535f9e496fc52c720cf5ececda60ce878409aa8a8179b4c5037f80756a8b9b72e5ca368b6af6c719dd011cca40f076a1a4b616870b3b9a07d60ad12afcfa8036999b1b4f55abb65817e5f7ed46b2539;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0e456e7e3899d62ea19367cccd741342d0ffb92e00b4cb52139c40be17cf2e473b37544e5989086ce93c65a24953c549490266688ad5e87d116e628f786b347261f68b27176b50d2eb3aa884565ea67132325605cf36e5b03a4a886fe5b9ecfd7bcaa5e2277cf71f2fbd5c1c2ed28d06042e51b2c7cb6a14c354eac3d2dfbb7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb88da7c5bf1629cba38172643c5fe84cb49106012b94fa091f4fc2b21062ba63de5fdd24546ee534bc01e4139b17375d59266879b6aca2e14a55c4d06b4006d7128fffb4e05cb99414e9aad00a42e76784f2e6379ca2c493f50631301224798afa5cab0175ea843fa353f3e70a7ff053a5493a608e518483a9fcc056566e2eb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2da47671bc9efc74b97516392b6b0c11fe621d5c83e7977ef5b769195c2f14e71d4d86c46393d84a6ef236022e540dfd175eaa4b5798417e76367ab6e6da059615017016e639f870f9721da2744c9e9c38ab03fd6b0fde200deb3db4fda22fce24ad67e028050ddb32b079440f564f7d8095dda74de081cbd0ee4b969335790c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27a914d55408b2cf192f1cc5a8e52cb8a1a3cb9c1019b9dc90a0a1852785034b8b19d3b97afbe22c93057bd51fc58c352c7d7bb095501aa8dcd0577a506398ee3fe891a846a2f57fa028c8f3346927f57e21e9638f350cf1af4332c3cd302359fd5a638469a2e76b124d0f47cbd415e8623ec4ccafab0ac2f127cc723ac4ac98;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9fa847b98203157ba842deb29b5399d9196e6012b706b54121cdcea68755f28a9bd9acbe21f98da468bef16f285d14e7e720edffca61fc7e22aa7a72db2b1216303c912f0674e3de94214a16b4aeb4eb1aaf36f8632d0aa7481cc1f3e4b7e7c3a0dedd9c1c1c5558acb7f3a3faef89cab95bcd159504725034027e5e262cf970;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6315d382cfd8b195dcff6671f5a83691ce1f5cd861c6909470eeac3bd03dc389ec64a45fa1a5c845ad49a38a1c087f9504d70fc05bdae84be3ff32c29041cfc6c1a967a04195c7c02b12aa35969720ab323e8b0059e00cb9662309aa309ab61046b4b1e6cce7d1314e8535727f36a05653e94f78040ff5850e0a9aac90a9bd9c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd70f8e4b2bb093ba13297b83aa3826bc489be28df075857cd4f657b0318a0bd20ee0d03657715fe67b42703781477169ca7e6d86b0bbd0fe38f24d60f9879769534eaef5fb1758305609968ab0a8fa0df985de0d442044ce2d2c78c620c851b3f4980377357726cadc1eaf2db2019923b8a4a89b61dbafcd03dd0364ed92452d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9393ec080abf3b7520b20d3d2cf55c2a0a6bca9db87193431786a7a261700cd7dcb6e9bebfdf3dd9447b54a2fdb1ec59860f05c4cf1be552103888e74ab6e79c166e2fb6d2973a8c2a138ff3834895fc7cb97887ff3043d500b8bba9aaab4e82c55a445f5232172db8af7babbf0a81e5cc1d54ecb2180c86f59696cc150ccbf5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2856914a9aa03d1f684423765a63a2f3fc0c48f632e6f5e37b5144ccec70c780979814fc800498e269e8540d054064455d2d834c3d25ecd449b563c3343f90e52f832550e36febb079969cc7810c59d416a30e24ca7592cd4b6c783eb7c5a482c1a79954b6299ea6c6fb34982edc0959a05f585419b86d25447d6614d37c4e0c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he42d68a67f622f92099e6e19f2fbadea7d707a382fd9bdaed9dce72cf4f5eeaa8b04e75a80d041ffc17130f3d93ac9fd4ca17a87442175b32cf7bd6acd4beb78b5c002d88a2f6ec3d1ba5d2472af7db43c9536b34db9b966e06cbb2675fc6b3f625fd6a794c43ed4e3ff1f81230f1d81fc7d5029f7b8b969d9c28c4f474513b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7cde0140376970f7351273f382557a738551ef163cf593c66e21b9d4dc34b3f5d8511c8f6030e914d6fab410ab0e7ecf2b9df182788a6027966c9d363ae7d1385210a7b750fdc7ca2afcbea67b85d7c333622d227791f103605043929c7320bd8704b09753f1655c2c12df8c7aa502ced8289a1fb596e16fe7c8033337f57773;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d031a0477f554b03d616acd20d0d72dea84b4e028fe8ffcc25fa7b624994abd9298bba34a56a300991554cbebea82378cf46ffc401a02627e50046da5d78925c534d99082d09d7bf81988c366616d0196a3c4bb590835f2af0381dcb66f3f0e1e76b34a8d5dbfbb976044eceddaa9d41e80b8bde5ec5ea3ad6aa29d40c73641;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb0877aaac81c64e9a0bf361c16ae79eccc8c3b161663c87aad9d0183c29fb506b55832d4c508f10934d27806fffd1db9071933f9ab68c406c135d24691a4262241cc9348c7110231f354f572d954f8198566ebc26fc9da3890af650128def48314d60c9f1f2952c197c39498b27b292893584de91749d3d81214806ff65146af;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h573ef1362b884557dce143f66c11c42c59d9d9a1c58c8a733dfb23184fd8229fcb6efffd31ecfcc09d4da66cb3f3346b0f9ffc5899986113ae885ae5c989005f74f774ca7c6e6aa43e0a6f0abc5082b256b37546d6a7a7bda424ba56d940c392837e788508067ed053c48ec467e3c8ae572463c3392db64d798a072df6668606;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff351202707d749448a534e99ae60690f1d4a03622b3b8f0eef9ac924d9ba31a2631ea652179888158440712caa561ff93f3bb6a8d532f2a1546d8e8d52bf0ae6b6df31974ea71c562b72a0b4bd78ab35b82ff0ec067f8f16728c00eef4391e432c64f75e0b0b1282b6723d0f18859da32f13053efbda09c7744296ed46d9d4b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8045e61b2dca4745ba901f44908e88272e1eaca4a36dd12baad52c7f64c852d1036cc848854040f2cf89bfff951547a7c93c6833e27ff5f6a9cd67c0869514a1f906f866c6dfa5914ed61d3b8283d32e9565d4c10eca3a143503fcd1e640023007d00f89d875df41f804744fff5a9a82292eb2a2f47defc01c96a089fe3bcbec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65adb3bff2aa8f1e5ca2dc7c3143eaa1c47538c2af28f12da607ed75d0d009e902e2a9d5bd01bc7dc44db4799f7898b02fe69ad29b33478f5c615995df5678889ae7e78c291ff9bc9ca45270ac44af59fa80ec0f6339fc042b86d6f1ec363ae9ad51af789a2ea5fed5a98a078043b8e2ca1ad3027c3bf349faefbad438f4e79c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ecb06b5215f9ba1fca7cad26b9f1de29ffae430e5edd7ea51a0560af6047d75ddb78178b62b8f4c21fd607c27a8e0edbb29487c9717bb0331a531bdf91ac9c59d757a7761e0012cdd894be8e3f183bf49fdd296d1a974e46674c2dbeddae896190d26cd62a427185712e96428557e31ef81f0dc955d42d5236437585bc758cb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41d37167aa5080180435bce12b47c4f4708bf817e48de21087f842d425c75765571ccac6e80070e7305a5b19755b262e355b829d7bfb251afa16f9c382e30a15a2438a233a49e021a4ef15d57f79bee38b1f63d7cd3f9456a4dbfb597cfbc3495cab9271a8eb68ffc3f9f3ee2ea942c1985ffa46ada456fdf8c44bbcbe703ddf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1def44235501cf719189323536ad89244d03ae2fdc015b00e3f7fa73211d62a0c98a4e8b771908d7025461f685009a0da54b550877b2148f4cb5b103e6575f0a18481529fd5dd84856bc9ec4c679cf945bf68e845a1e0ce227cf42f46f76b0a9330155dfe8502dfe29bbd69f223b5b53c22030b5cf127c4eb056ab513aa4f85c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23c739b7070ca9e79ca72d818d3423545f68dd4c7aa0739a50bc0a1a30dbcdf0d0daf959aae1bab3050dce1bb108f8c6165d609e6b7bd595ba78dac1e373564e851dcf1a00d7acf6387bcdd478fed03ef0d9b3d82fec21f2af1e3a3a5ae0c1a31a7a260345932618185c3c6d4a8c49c70bad3eac28a857e3432786241569a36a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he468f2aa518996e1e4dbcc8c68cc02ff9671fdf138ed1274915e1344da544bd1dd3b38dcf49f4adccb62fa1023a6656877c4cefba6dbf52c87e06fe73a2fdb8299244c6e6c3511c2f8ad8efc1af7cf78d34ad40d1d427b03f96d8ab5d7a4f1641edd187ddac636a7c4b7270eec732fccabc56016cbabe8db5748a7066d5b7064;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he98bbcfb921d167b4b4cd1a5398ba7f36774c2493a57545286c2bc9355c588a47188271cae1c8c9a11e42426a83c02d44f2bb8e7d6e01798b388abe6a1a963f8247e541e70b5c2d8008a834f86211c3462efc2c8414fc8e81b3c4de146ff55e48b7a8a60679704af62625b611ea7ba5db2dd8efa679f6146b78eea3e9f9c9433;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h221d8a8ac463bd8c95684798cb5c2315632a6d5e7ab41a0e866e82754ede15734d6b402d872e187afeed4ed06e0b0c545c620b784bd15fb4e5a7bb443675ea68a65db0ba15b847b0ee2573be4e14ae9849b59ecc334cfd16ceb34b499266979d2d400fe5481fa878d1dac3f94bf319111269b2b26755af9176752082d3acb5d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a6d07eb6cd0f660c166f0f6a4bd24d1b4a935a0c6eb53dd9ab8f1cfa2cc18e1ef8084d80ea5245463fa188c3cb01cf4808c4b0fd3b7c7137e9e095a1e7b8ce3c7836e240baa9d5b1c30ceb10efced45197bb5ccb0695fbad87694d8f7d8926898447133f7af5b3a38206ce115a5d94ca9d54fa15be0c6940d833c721c24a20e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbeb0642e398bfc55ecf7efd94561f8401fc3b5d559bfdfbba0489ba0368800fb4af752cbae49db200642b4365edd27cc0f295569908e1c1940658f57457d792fe1d50efd2e6a2a8058819fc8f8479bacf8595208c91b5ea012b983dd42f05f0e7c51d7fec3c29c2d37afd97d2491e2bacbd736b22569f2c65ab1481ede1d3b73;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b2a1df099d5ac04b716435ddc2c567b5322be10471474bb28cc41a2439b1cb1c2a339e001f4dec39635b4b315aecdb908e5598f508a1c3ce990137dcc66e124a6bb898848b4387a2559095e51d72e72f9e9bcd97d9309a61dfa4a5b22220c9e70922e5ea544773e178ea0aed7ebf6159844e05f8c66188168435d12254c6c42;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43d82ab2d16914f7325072787706a500cf2f99589f03be0a0967f4f77e61259d75141f4972311c183ca646c84012553168a3fda6e58b0af6ec3fde0a87a9ae5e70cc9ce00b48c64e7badfc62e9428fbcb0b9fb9951e603c01a922ef070fe5cb17653925a4448942704476a67d856f1a26ffb89f1080934c6e218c0621ccd4033;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2a1820f08c7cf8a2fce735c30b548f4a1fd00c8a48f4b651d084e01fbbdbfe110bc300ac9c99e6b7d1bfa16b11e4c66a7862517a51e7ebd77dc769f94fbc4ed14ea72a47a8e27077f24586199d0e13733113e482add205516f9d2bab7dd39d22046a225553f79afe06d9e305ac720972cec61dbcc6eaa2dc798053b23c33f23;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2390589567a3956cf01a3aa30d859f2ef871ff699f03c6ea4ab3952a5c57ae4518d92de42705577862205defa8b7cce9bc627729b10832a756e8eb9cbaba0e82a532ad715c278e7cf011c1f54f6fbeca04d476b85b1aa52c4678317a29fb318ee4889cc962af3e7122f484ff2d0e49c53727266a235e78ad9905cdc07e85d5d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2a095278983eba6747f6f0a472bfb60a20d7f6bc8b14840351674f5fb7026c1dbaf114ca7264f4dc809a3ea1424993334e687712c4113674365c39af8cf90436a079ee6b14656479a3cf62e11bd2a9fb67cd9792ac3ed0bbb743650380d39b752f1139cbb60a233fd9bedab4aec5244425e183a46867bc22ac7df9a855b6b33;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h387af982cfa9a76481b69e7482596ab92b879ce2a0814be2c386e7b8d856affd7298f1fc66179e38ec3c10b7133fb9231c94562d9f15d546c9a04fd6d38d3f5d6d0cee3431b6457feee83cf76b59dc4ce5f8c3358b386697511b05b7b0179ebb787d9f6f64684a26560a8b3aa298e436430ddfbce3cdafb347bc5419de936c99;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4303578b60b222ec4ce95e7c7b96d0ffc75d9c8ebeddbd73df1e7cd74c44ddf72abb60624b1fa483a148762b55878f12e77ead8688afd8bfb0af60e07ece7074bae0929debf1bbf931f16449489f51ba61db5875aa693dbd4b61a0f18a20666f6565ac4a01ee01e2475c2bedf351445aad08f56007155ebd9532bbae6db4069;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1534d5d66cabe5e95daf4e5307b6c1808def70ce335869d3923c57191305531a2e4a27b8748182010081f5e4966aa59563d8569827f61012225bf077ea57ef84c556c085484fc4a7577aca5525056ae3285f04ce4f385180317de418a9352c5b5f18ba8321bea74072ecba4aac37365d389ef96e80c21a8bebb2e28fde803b89;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf62d7d53e6ee95d16308b8906243d3e88a3047f23c9ab5a1ecce3c77c553d57a19d64d83b539c6f5a95585a43089871012a9fb03e2a3e3c0bb1eabd55fd8da108bd96cf7fdf2d7399815e53cea0a615d7fb8eb4c61094091d34440fbc552a78b089b6ef28d326c4d5a0d461c65f6ef46089a7d9e4757d7f00d576059e25ca6a7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d9b3c59922c6f3d0367bdeec515158e7bdecb1780c89242c3d5bae54975c6c453807553b187e0798a94d0cc3bb527ed687d9cacecce478321109d37780ffed9723ad9f7049c0780f707f410920619a5c46f8045dcef7d0d63d7e7ade395db09d7af9fcbeebe6b4f9b7d38c7ba166d07ed050dd6acedb59c2a3b3271811d7515;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcea2b4fc8bdaf6a8475b04c54438e82a9b4a09f6def680990d4b0195eb788b8e25a933ac4335fbfc4a650379e4eb7932d5e11ef791606d5b799afc2e8ac437f85b56ee02ea9c9912ee425010dc90512d616633cc3f72901ffa70c50681f67853479156e6e92cafc2823ea415dd3362f46b902dccde03c3940d22b4c4f86135da;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd803a9b31d0f0ece0486582c995bea96eba6b377e51be6df7ed52c2926a6389acb1d414fda2870da4a3547765095a2a8a4f36715fdd84a711796769a0f5f710b9e25058dc660c3593588510ea70643dc34697e947a794abb5390a9dd290aad7fcd11e5dd24c2dcb0eae2535a14c5d180fb0dd7c32209c1b537fb46327df0ab0a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9572c6df99d9ef3d2bf05996f2e327f91ddb830c974d4c50d421d920dde2ed5aaf481967967f1a9bd409af02bcd1c4fa58b68aa35b2194dea915e7f87f36e7ce90bd2d4b1d5b59781e00660d223eaa290112e7a45fd3798659c12839929661b0044a4460d9f4065508d63e1f5fff170cdfa37b76ffcd32fb92f84d64c7a5650c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6adabc2374e1c67a15e360243079092e90e9b520fcbd4d55425563f69c69cfdc09aa4b84552a12b7ddbebb608104f5858237dd481c03539300a64e4fc710072e2add22d81cd52d58a88399f2900056f3582f0ffabc1df768f37ea9dc25ed60ea538f2fd524863f72587060fff63cc6ce6765fcea06f71b9cc81d9bc7468377d7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24fe11f1c3c7a8292fc4724da8ca7b4607417d848a59272b7259ed73b49a912b537295fef45ee69cc9655e9e9416d95ee9271bf1c137b29c0221ae6f690e67f1a23ec3334b60283a5c8dcac7f4e966b546d82895bf7de5363268ebd62a52afcf99bd61cbfaf199082a5ce18d686a4f5b71e44ae284c86ac89ec844b094d9916;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had1d275426116f70c83f7c8a73ba4bb0bcdcf6985aaeccf6e63ec1b910e4903d819d4c2452c73a699e317737a0dd08dfcac968b6edbf180b55386fb2a06083af4098390c5ebca3d7107bf9a5d7c08e998bac4b0ee81c971820acfff23214b935f67692e0f86f742e46b33fcb835c5a3db55f03e1ea127766f4c49c516729ce52;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa3f3d9e20e128d22d0d2ccd776526e41f89604616a339a8fd47501f3dc8f5a544fc1ddf8cc4e95ee94a3e3b42ec70d5de274a47bf095e6aec78392bae49e97de5171191e533aea4e0a100dd53cc3b0f076e93a358798d89cd0af761b5963817dae3808618df2a64d073886d6e3146ac948314233fb24b1b516834181dcd29b8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e1de5d1bfc803f0d48b6eb92822870647c9b11c8e3be3a92c4c5fa17ba87b0042c13c5d559ca00d2ae14e7f8adff818433a6b570b52ec6adf0b51e2d44b0f52245a0005c5dcd626e3fbfebb652806f987314cb354965c83df33732657f58633c473dccb74ab21d095e472c67f59961d5791998236d753284e8bedba085786cf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a7553d5c744e5cc1ced56c449142302a1f7d73f142e46089b993e316174d0d40cd8327bc212a4f7d0d54d8e446757644292e3d2a8cb7114c5b62e7d9745d5e2d2c8162d9cc9a29e8a9d5b16ac29188ee75f015e2424b3e769ad9d535ba6589c9c642827fdf034f7f70f7f0f9ae4357a401eb18cd619b22a793e93a2c2c4e3ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd50b710db2b7c5ee1af098de67a6362cef9ab34cc95f178ff21686dc6b0e39d49ac42acf2e7e60a9771d8bd7f48891775fde3a8117f2ab5bc671a12101830ba81f99e7b179e899f533e4020f8455dcf81657b949036712ab02564aec29335159543c4adf14825af0facf8c3e42a61fdc60c1489da98eb2cc77ee9bd1a436efab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h249d55589cffd2ae0e7bfa5283c4f50b247c84c467a760f2c484b146f63c9b14c40cb7a7fc75e21bdbc8d750d3b0a1cdc6d824783c27ad9336f0d24d29fc3e5578e4e7b292151dee6af7ab7d03e1f20023d35c6e4d5c480e77cce3d25aba98f285548ae80a0fcc177ac8df03d1c1342cab3603c000cee0296bc7e7f6ba0ace40;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22ea90b431eea695b38d56103bd6c094a79a7fd2c2745ec2dce5541e2efa893febc4326aebba8f24ca3eda2a2a07de888a67a34b0691a79f19ee89aac3590ce847fe0eec48750348541b113ac27138495d6e6d8660fe1ffc621078e476a19f32cc6526f9dd1cc130526f3764a06db68f1b0933962fc46062fb082f3c562e1f76;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1a550cf7ea97dc86d19e8723e35fd91539af7a694b14175115839dfdec83819c5a6837764e4496fdf80a25a359953c9c3756029e07eba304514c1bf8198fb004ed772fc9b040f6e9b68a3ca921f0f63587cd4b9d2f3d97e0871a1b8ba3fb3e76d742e44383eef324b6efd9dbea1e1d95991f3eab2c3d5738f54ff66fd25228a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8be5330d6c2f9c8e723448d904c78c0a3781460273c3620b8d949cd36aa4cb3595d184a4bc63abc02d42566d187317748b7fbf715fa61a4258d79f7e0b1531f5840106713ba6c4c72ac37484e837b0da2fbc40dbd68aac947e89e69ae5feccf6b94b4651945780da124c4faf1a866d43cbf4dec279661f569853d75c2d4e0b05;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac352f76904a34e48e450d286db33f172c63b32f00eeb48648444fa17bb8e3bdcbe2b4d79273a986ce3998b45d3fd445651a5eb1cfc130744a71eb77c304f4ce7950645d53d272e5b9fa8f5848857aca222ef9fb1a6b99660ccec37531b0530eff4db5f0e363c83837a189e4dee32b67533a140380622bd12369dffe0f4d4a7f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ba1a57cad2fc708b204e668841f3d5ea43b251ccd0fe11073a30fb5a2d187a7265c304d8103d9e12d83b14177b7d6261d37b2463833d92d93fe320ce00e9d81936d2ce68748065366f0fc56b4769a8ecddc2f7a7441127c4d8df58f3a930e62bd990f556a7bbd4b4753e92b3a7d4966a9b2d5f73dd1686c06311007eaf70466;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ca53f259a4dbd3c1024675f6fb8009a1223c2340c4cfd3c772bfd2ccf35914fd21558f9c622c981bcbe85d86a7d1812f8bd6f96a1187b654ecc1ba2cc899e394f3c86d756e477fc604bcd32ce41278ba7fd3d901aa3dc0adc70382e03a0ab6abd4c848452d4d07ce7c42fcbbff0c37daa4a30f7c6de0172f1ffaf3e6a4bb514;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd17d988d5d1d975905cf82dff0c3f56e191c48cd6ba6dc8c7f1e3be3f2cca25194a069efea8a054f65b393e14c5baaec489280aabfbaddf2803bdd5ee9b40bc2d9499b3c591a6ea46850566f5283d2cf606c81853acf340ca3e7ed5c966f2b7f060f652996d930c08f360943255eafd6ead2754f5a60d65d2f739dc7bd53edb9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hafa4eb0c3a7ce78420280a728b6a1ec29af2a2eb41f8236e0cd2238f86d52d999d6e1053c7f4901f3a4779e76bdaa851bf1200c0379120dc2d2de941f9481421cd829f91482886a692c044e33bb460a5432beefd2e2db853f1038fd6f1c44b6a82f0e8126f2e13623beecdde94d82b0445198a6a3c7dc32c2122de1e00c7600f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc02cc5c9e3fe0dedd4b4dabd09124c62adede109ee3aa962600569261d5d14f7096336e2127eafcb061ca272d1636fb7156ff1f4e8ce99fcb20fed5f8c1d82a0901ff3c02e1dc0db9d99d77732e3cf05250348cd12e51e61b170187b724af82502acb1a160b9273c29e7029420b03676caa13d63c7f692b25d4ac192e167321;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6938a6fe37f644befa801916e8fcd69e589a1fc3a62931586611f9609e8866aeabc4837e940450ac27d697234343e41f0c7e7a23830e398724c33ebc35d3bb70b6215d600a3184717d1ab7bd5277c71ffbdf53e2328d641a7315087f05a1db631397a90db44602821b80445d9f698fffa822d96301ff825fc35cc0d8a60adcb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5db5548571f2600a93f8a2e9551a8a11eaf21ef38bbd9451d7c797a5781431976fe0c275afc5be83d30c65fdccf7ba6ed42302f592de3ef1128d3ef8dd9cc056ac2395feefe474ad8d05736ce9205c9b5526a750aaccca7a290b691d316b5f2679fd0f8067e83d62c5b2916a4392ca4b067dcda7dc7604d3e75c3c15be5ed96;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7500681f0a85fdfaa4b2624511f3ab23893c87aefb65b49c72197edb4c11a0e64a5beed4dbfb0026fb960c2a6adf4296c7b933efbeb14de95a951667e1fc6fe5d0052f6f25097e55d7085bdb55767fda3da49ff1ad1d459c70770f4c8e840978ee28c7808f536d3d450ef2610a9a10baeb5bd49d72e951218971ce0d3e2aadc1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c8486a7b12fa890027a97522c8fe7990fc87def8b29a48eca3697f433c17744f5567be6832d39729ed326323b907b27a0dcd2932644349f9de119f23be88490a78437697d0673386ca9c7f9f28569d884386e870aa62dd4e39a40adb3459780feac5a44f97fa0c974111d80fec4e079e732a8f8ce319c1a64adf0e026f86218;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36a45050ca0536d8af705b1e6b5b2fdfa642f9efa7af4084e5a4980ea31d85b956d8a9ba480f0dd9aefa8221475a9faf98bc3e60529fe9f0f19029dde85ba85f28b7af853fe102aee32eb3868821bfe6875ffed4a7ce26d48d5a4183088832e6df1ed9aebc1d963b5430c8adab47a909247a4758fa75a814ff41f0fdfa680bb7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa4e78e7d3933bb1358ae881cebf8b30939a149c5240ff7f3380d19c0426a78fbebef7408ddc7245e8a87dc7aa59d0a77d6126542671ee8bc9dcfe6a137ddfcf03a74b34ac61f3c3664d3c931e54bc553d20cafae784adfaad05f47bb72f11bc10cadf6ecbd1405bacdde11baef9e5373e1cbf50bec68f7eae536f781675add8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h590fa6947979885bbdacb146127b6bf63ff78e1c5e8e613fad130c0567eaa70d6934345741a31ec465f89de6a6049ea2742ce5dd2d15c9996f7f2d44a70d7eb09fd17bbf39e06dac08c470ede146a417ae91dffb73543f91c248ce7556b181451cb983d5193c4330f54c70bf1b75ad21dcd5c89237ee02cd2dba2b2928dad9f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc6fd16f46678aa357017816d43e9f1664d6158ae872f10b33771338721ac9778f574a9fe5ded8ac65fccc0e1e1549d1c81725e844595ce21a4b164b56b7e6b693a7eaa3a4ff5f669b564c1f03851f965706ecc6852db7515b8894ff75d615ab6314d95b5e17d3f1e62327933789aa10da5711c2feb40b5a6f5690825cbe50d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb0cd3e78569c86417d9d9d1da053bd78804ff8a7bfe06e275d6a9daaf3b4ca5b1c4c0ee52b460454ff245364e3a0cc4a3dfec701078f302b1aba345a3a2bfe936c41627feb1d081c910feb4cae855d7b2a5c8b6ef094e643e38de0d944dab622fc4aa240113b53961959171f27e3ede41700f8b125dd4ebccc473b4763eeccaa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91f3efe074078712c9dd8f6011c986b311a26fc5bbb912c924e21107d260fe913364acaed10f9bf7a5d50e5af0a1e6d670f4797476004a469ead035d273d36ea2eae56a6f0e85832753a812e7150133e7cc6df740b9d30cd7be99ebbe9cc6b3618b82df4188c44c8386079e33a7a2ae8d23adb9ce57cc6df7ee07f08078ad2c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h148954fdd606b236ab5019093da4c8a31a67bd0a9fb76a19cb9976394410cc236fb39d4c6fda7f0eeb4959ee51ba1af5e3278743d4da981ef9fda74d432d99a51fadca8ba6976be53e6b80c95af6ef698b871fcb7a06254002999c66d78867b67193189363aaf7670d460f4ade52af4fb1f609e07c50fa03f5ec23d9715d026c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0a9897f184afd6ad5e0b0175c7c272c07eae990754ed43063533a59923513634bcdf393df05ad3a9eca1c05fe2273e0a395ad52c34467f2429d0827f4923109e2edffb4f03668ddbd5e25f05363263cd0f0f24e8dac706c8016551b4a7206a15a8a328e170c3dae65704e7c0eaa83dafc3aacf97e966b25646aef075a4f8639;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc20a70e3566c6d763515525d1bb58a7184ff8aeb88f279f9522dabc8c7fc3f29889978b062ca1f51e3487139d740745a4587745b10e88c9dd6d25950597841f6891f470ffa8749f230371c6b6136b664405ef40688dd33d66fa071af72c29d551675cfb4dc6e5e3271faa61e3633528a3e6213854cbc35932f635ed87a10c584;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd0b712f9227d574c47cce2a174e978346254f16240aadab14c470c0057c116e4d5d425c9acae1016156072e559c67ef136b1eea8dded4023ac3de4534c540cc9c8c57a1e42a051e5adca1d8dc8d691c9ffe69372e9297609147f9c6f1f649c27258f2aca2520ddca390eaf72b7a82b0a6acbe8d86418098bcf1891a689d8a01;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed678cf052234199ff69839d01133975618eb1f3e1741ca6d13f6582d71020a82e56d3c8a68ceb27971deba0684088413514c5ef812c0b76a164fb671326e08530cd2e12e84a27d16314e3a262bf7bb8aeca848340e5d685c6e1507f009df70a9adbb419d3bdbd9b08529eb4a4c4d8089d655242648eecac2d433c83ba876e68;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e8cfd7b9ff37d0a875730e3d110b389b49a8138a4623fcbbcc267c69733fcd9c63f4cff2a1f376f7e8cf81d06a2009d660c6b650cea48cd3c5c79c754c5c75d44f10da96ef9d562f1466a9333560019dc719957f6b298661be5a80645280fb866854834bc12bc566d84e488dac1910597882c8e365b9d0bed7882531f0c2c2b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf3b45034776bc5fd862d5642d565b98b967f51fcb38afe92a4e3b9a5028beb6f7194bf13f46416e722b67a035bc6e9fd3617fc06cc92f46922c156355905fe79feabe0de24116483835921d22b9fcbf10bdcb3a58040ff27567c1e231fcb59938cb86669927b8200e76f2f13489bc118f1acb59c5d5a63bb5900f9f1e44a14e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce5e5be2661b0241f2296cca20e8d0b88b5f6356cea94931ef3052715c0ff991c372ca72132db954286d611fd82bb2194fc990a6a6bf9169c5e8669961e85dcc07849f8586b44b848aba35e28172fdc8f99f809fce282d4e166fbf5e1520139c849143801f1ce6387a0ce9f6e1073bbbdc9d3f50514e0cee47657ef50b32ea44;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc528f8fb7baaa787fc63f3e956f8a7e0c34cee439c7f85c48ea99347d81d151b110d5cd9fa1f59dd1d38559ded84831f6b760bfe9df05d9b92a6a2c0f9cc2cee81a57b68d05564c1d507b5260f13e5c9d56fd959d67f662fbf6c5e27f2af7aa675e41bb6df4a22717d298994403a296953daf0d8ff353798dcf482ea715cf9ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a5170eed9bba3afe455609398824400ba7aa24446f6c5b1778662cda6ba61d3d602978f4c35e2f4e427be76468132740c2f3f739a28156a48c7caae03caf5c0e9b6207122b02d225d7a8d05fe0693c91a730651b8b9bc8181c20bbbc922a3243baabc98c41f38365487c5e1cb1e214c338b4e4ba50b5f0cbf9d188a77cb96fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a6dbf36d3b7884c8e44ecb5aa382fe7fb05ede9e9f672c5acc015f13e4919a05758da83512a290b71f281445c203e26add7f1706e4e532e381d9f72b2bbc8c68269123da1212191f153fc8fedbe78e9b316a50c05a3a21d87593b818f088d77110802a242aaa8a32f40e2bf51a36e4d3d089d3f048995ee7bca177ad65aa6e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab7035c2dee770f622339ba00a9400f30ebf3e5d98e6d43716273bcb9893facf53a2fcb61c2eca431501986b0b8a7c7dcfbda4ba813d270a40d681662e3c5f63d7bbf45e8d4114bce75c14869c6d947f6558c8f4cf47beb541128471079883478a55cd0f01a68f38b5a367cdc8c77d07f8b33de55f2acf802bdf4ff65068cd12;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb59cfba0754c8e3aa987647eaa4a4abdc9ca021309e3269ff261c86f6c9d95bde0877c233ea8fc4642dcbaff0c39a063c79d2514355f4c87474829abf47542a847d6f280f9f6924975fe3f55e52a5f7b90a0730d79d51332e1ede963cba99c5ddabc38ce478982f3d01270fd7d86861d11b343166a02b683ffa81b046e13d36f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4feca2e727c31c1669a8601abf6e3c7ed7753c9afbab279db4fc73234f5eb1a637abe55d63c0195e5aca8cb6b57eb45907363823238bfb7fc24de0482e849d1b3c808eaa3792df0fe4074de2927adf5f47eed1cd7312635e489684a929f18759e9df826d4729390a5ca37c6e67f5bd12387161c7b882f76841f8d58c7fe7090;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bb58b6a95596f8da347304a48e38f40be2eeac7e3ba1a8bbf4a9e25da5a947668068d537231fd6df0d5e68279d05a93070fba79f4a7df72328a4f3d4d2ae29e681d356c52bdb3e215ed5473e96efcd9f802e43b13466cb3b5a0fc5d969051f3c160f66a7eeff0842f37f0648439a6a07450ee8ca388ce6bde79b156b71e580b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha00de5685a196dbc7226cd6743f05008a6e379997561ffa992b57012a400a337524d56a793638cc211e689ca8b31da7f5144344a1908315ae0e30327d7fb876cd78623ac627f192079bdaf4f0d61ac0a6e0217b8ce44ca3e7c4b1034e76c08600f92106b8795d3e3bd6e10653b012e37b90fba441b981e5a8898f803019912e7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h44e5700f14b9d5139e9d1461a34b0e083e10e9e51786c24ce3b1e3a36ef4dd6ba54c09713c04f61d035ed6f05a61a203a5835a0a3d3d427a5f145d3745e933eedfc7f87ba82b0d012cef179327acfa84ecdb610d051052523174a7422ec90dd2c6b85d70f408f06e1e8c0e4f1a83f10f442b12552511be6f2f77297dd75f6548;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70593e49651916819c9941d88b128a507b901f3daeb39ddf2ce76bd73572d7a4883edee01b0c5d2b8857aee000b01c298c16987345624ffafcb256fa6a69e9d5b391e33d68b50d380f60ca337587eed2fbbc5805d47b00daf4478d06ccc4b7e8475020e49dfe863e07b302f837891ef4008cc96de03426007eebe44d0b0ed39a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32744501ca44d15232e3602742b84780ae455175bc82c3ccff4af44e0b3f37aa8113305e1ca688aaab16b4b39c0726183f6f7c85e64fdd5a8f3454c36521bc0a83dd5ee923676919ed72d5fcfbd3345c0a39c5defaa278207332dedc5ca9c8de1f592940e35f26453ff489309577f5fac4585e9a7d4be7e6d5bdb7dba648e7b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28c83f626bcfce78b6a112fabcf7ea0b2beb564f47514c3e3e81ed6c9405aa9c261e2659d7cc25dd91af82af3da1257649d3039466f29edec79a820fa7883166a494dae5d60d4badf6a9a410419e702603b00c69013de67b8d4ddea112b077e22f205baaba5b2fe436117820e120196095982a9f4c598ca5379f71a6d6a70a65;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3623b1b6222a46f00238783063d90ede76a197b3dd9fcc3a305dc74f5c8e01a19a8430094dec24a0c8652dff117c2e97ca7bc366ef16c582626f40f8feebce65cee567a2e23569f0f76edc1ac80e3dadbe2cff3554e855caa7d40e8bfacc67661388e001fa670aa2a70a1c5a9c5d31645a529793b06b5c455b86a424f2befe9e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbae843b31ecf0f20cebf7c59df12acd556fff110317078267de46a4a0ff1935b290e8ea71d96e7cfd299d3d0d69652a73ec9d3e4469919bc8c9d23d17dc4e7ee632f1dd8b52001a3108fbf45c1af6e4eaf98ae780ea20175c541bf3b6e1941183d663c6c701ae20cefaeb8ec924325f7a8f7892c6a9739ba914bf23a5248adce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e80388d5fafb7a8eafd8e55cf3fd1d5555f6d4237c3b39accdcdd4495cd1f5b1e3635f2e16873122d10bbd818cfb5bbd1d1d7b2c004c359666a75f4dcbec5d0f24f36b817424bd604020cd994ee0ed726cd291f594d76e99b11d2e216f8b5cc555332639f0a3eb7a22d480fed5e652c190b8da233f1e2ab83254300fa5b529e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf9648aa468015c23d4edafb6c3ffcfc7a8c4f118cc1546e15169fae5d45340f08c59179c8351f5726ab405e14b17370b6de0f7e83208dff0c4b3a3e4f9b25ad65ce1bb93ca6fa9dabeb5c193dcaf86b10d4176b70e95e23453588f5cbe8b13d5f16bbf6079210fd4ecc0ed55a5c5627cf4401ceeda94aa2270ef788593b336a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5ad0f93ea6b3e56dbae0673cfdd2ce82729bc468d6f160888702c91be0b9938ab129b51d56677e7dc140d4922d70c1aae1861e01a7226505f600ea20d5896b75a86974c545b6752c1cb6d2b43e2337ec31ce97f820dc3c1c8ec09605b777b4ba1ee9c92f4fac1be33959faaba5a24fc22f4f5890664eaeedaf987fba9619ac4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73ce9bbabe3f8ea08854b8fea49d6a16a592e1188be36a2bfc53a60d9d5ada8e502328be56ef399b27abac6127c17d7b54e57777a8cbcc7c646cd64b5000a7b3f7a4847e95723314187d26e59952d4623ee030caca8c02eeff41fc7e15487573d479066319a82f325b5cf2199925083a96deab18053b799d977ec9def4b64554;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc51c2eb9c581af43a9737af638022cc332efd71bf1f83b768af8aca0b621bb31f8683b04e7fb7c10158c167f67edbe90719e3dd16a91620aaa0fb84d13f25de22ca5fc920ae47d1651fd6c381fceb9dfac8f4f0cd77efbe816014f56acdd6937d3fdf91dba6d876062e37ccbd91936e47c2532ebfad50f4cab98f30a67d5954e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6fb9a9892bce9fd91263deaee41a56bb016f47deaab708d6bbacced8e508a013354731d65f649af09a21d9fc0ef51a39009cfcbd1e21d495e7768cd3b85d0707c31c82999b9aeefab355adc9ec0fda62fb8d9fa4d5756652a3c08e7267e67af06c727687783a2b5713942c13cb131adc94fa94c8f17c1ddbd97390b7a1e5126f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8959176d69b463fd730bc4af15d7789eeac03b928b9181df06ad0088e2d390cf9fb6e04ec111b19381efdf3b543b75fb48d4abaa9882783a3fefec29232622500c0d23bad578753716b2f4e03e0e21713b613b33e32944925178295c2feca1aa365d23887c9dc5b07b5605d9e0268ad068b460f6323b8cad8dfc7ba1aad38f89;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd50d7f728fab2373928964d4d1f83b746f390766e59fa78408d586bea1841102e5d052126eb6504258859a175ec0bdaf32d3526d91d7dc8b0272923c49c1233d98b4b493dbc51ec73421c3ec56ff8b4e38716b229fb85278d77fb578d482123f508cf91ad127fa1ef736a9536b4102d61fb9042280de001f52eaf6efc2b5464a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5b70a46e50069d712c34d391b00de4f855a89d00598fba91685beb6ac169ab387d2b4144f812b8078ec2c620b65238f4af8169620a8f90b3723b6d214f2de5752800d3fcc278107aa7f7e6294a5f1906b9f6bc43760408e31d959aac720406c003cf0992764176d51f3230152fe0b49a70b78e2c2007c7f2e9a3007d50a518d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5efb795f9a59018f672d981728aa62a5224f61bb5331bf479e5d95c84369c794ac58bcb53ef3cf01d46f25b5a7c52a5ccf39c766f9550e1f2086b33ac3122e6bad378a987aaf4ba99de19a01397033fdbec7a096449e480b93c5db53ce953436f3d0e18da5b47b87c7f088b98952f1a4018133d95c77cf1cc24310e81ce7c12f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha41a25914bb4076b1551fc24fa6735da382450b92e27cda99bceb900efc10e24b0496d4775d77a63101175ea90b694ee39fcaa8bae269457fdd79c4a4ae3107fd4e731766330f619d36e05b84a7cd3c076a5c2dfbabf86ede649556240a2cd9ac6c94a0a3dec093b5a82f91cdfcc1c6a928f93dd14695cfcfb3d78ae62f4faad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3a2cf031791a829356c978a41766245922719f55938a023c9bfee5f533ea883ffd7594e152dddb0dffeeee95be13b0180712613aec6b2902ec4896b8e7647080b2d917a7e67a686606c7682f63dbaf44cfb92cdfafc583552ab992ab6c0f2033ecf2a65bf6bc78d9e3db5323dedee06504f81dd1a660d3f7da324cc4c71dc8d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3f16709845a9a66dbdb2b657046deefcb3ac0b929a2028272b91e0b3a092f3e923b7b26fc35228477b3ce5a3a924905e83161590ff79dcde375bff9bdae7215366c6342b2ccc087ba604ac4f7df2cbd8d313458b6b8f8ee1c15079d60edab9c9c0b211bd53baa5ab07a6436159fb375e6ad0dbf993fefa7cb84894b604916f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ad54039838070ad93324de603feb556ed8ed2e9ddafbc7be392121815830904255c277d5f19586c9adf337435c4fe1b8ae3451008741e04cb262fcffa5ed74d8c1b93780ffa7de96cccb7423363feab0b36170b6429dea55bed8538f739e98cce80571a11c887d7b4af8327688663bc8dbd0a78056e1c9d030ed36ce63329a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde7f815bf319497eda50efa7b62b151de65c2682beacbd9ecd50af40515d70cb56afa1e35bdf963669d972baf6e55030763d64773aa95e739aa047a06d93d5b746a2ef680691972ad60290843b92bfcec41053a7297f585a70438a8eaa4e73dce24a7717e579c321a3c043638c992a51568cac607fac6290ac5eef98a1adbe73;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe6e82871fb8dcb516e8f58976f007fcc20c208ba2fdc39033cc51be366c9eaf3cdd26e2fd6be3b1abf7232f06d7b11f5401bed0d6262f579390538189e029ddfaaa4fb50f61b90bb75febdabd06c93615a662313046b07c59af204d5834e5dc9e8e414754a9fa25d782870e4e0dacbf8a0491fcb4686d3dd5e04e81f069f54c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h322a92adb1ea90660392be1cb7a58b59d370ee8cfe0f129ea27731fb6a303e140a35799221c12156b1217cef7a669e573cf2e04a77047d59b9fed0bd6762e5ae24c0af4d21bf13082561c184076d1709a569039e8a9ba383838dd7d17395b143d338f65640085b7b7ec00e2d55cc93c9baa468986bba82aa6b4f1fe66d7d62e4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ee968c74fa23e63e2158aaa4a12c150f382bbfd771053dd15d1d0861548e87ce0964f138fa3f9f14c14924d836fa198f6f66b5c7a60b05e0d6b9dece13b8be0adca1965fb952c688263f76d862c6c9cc9b73bdf5c9d23b49d6d5511f209843a83413a9db3f4ff85377bfd6b22f2560fbc794b2c55b75a2e17c1970f589eab0f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6aca8e786aaa01d8e83168aba89c3a020e92382e85cd15fab5becb551673b50bb14f954665998249ce92f01ffff4f3c2e5a76125968a68a2331c2a0675a3bd29ed031847e5bb3eba9879d731cc0c5424f1c034915c8ae27bc37bb99bcaffd7ce092e16641a3418e60282f7879d0c59b64defe3d648745a7d6c3cd045792a1c0c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5539e3d38237523f619edbe651e62421f31c9c0ecd4a7345d1b2c5c6955f4e0f243cdeecf49d5a0352580d2a2126618205bd586973e22a4613bce2a37c3603162a4ceb2896d85c9301e943e34004849f3880c37c8e5d9f409992460d233fb000842b942788fe372b1a28e4dd7c5940a1744d3b575844148e2d62ff4cfd2e531;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h455a19c50767438165134618e2c54ab81c8c73665bdda97e73437738cdc0d902ecde5ee45afb8ab0d5f867121ebbb478a5c2984bf9391201ad792bd67c266943a2c2073ae164e4ed09be8c29e4eae3acc013d9194f31372522c1d3ee374c0b14cd112011dbad3f8c3e71166135ee28f395a68173084c5cdc945e4583b8df51f6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2dd78f17452164f87b2d839c87bc613c8469e43cbba1dac8ec13363798c758df23396a0d4e85175022bf2aa742a0421b5d3a4a11cd6759c839d0dcea289034b26eecd51dac61434dabaf69763b2dc60020a1998a714a83dd9f124cd96fc93f02c25587b044d93114d3146db57b6c7c911c4aa8676a6c539adbde0958fd1bdff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ebc797c32eb7f47775113d3138962c1d114b0730c9606b35b8a43004f03b6abe49cc31d48270e2b00505b44f49a42f356edcfb756b6a822b68644c5f98cd83cfb6f35471a3cdf08cb80bb79cf06b9dd4b6d0cc666c9ca2447ceb98d7a6044a991364d2433c7683f36d26c4f4b3aef3896c80f69c58345523ab50c372225897c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e1d7747034e0a0244deeb5e3269dee8d7b65869a3375ad3c53be3113a006512de30a31d3545a4bb6c8f7d1d39d72dd235f9efa3a54e7f7d082a0f36aaba56741703c68b4e75aa75e86c81bf38ff03a2df0693fde66c1eb003a2e3cb94a9726dec0b1af18447cefdd5b7172e5f9798e9ab728ccb2e010169339cb7cd65415ee7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a293207fcf4402b77f33e475e04f2981dcef16080071c9268935373853ee0370b1b2682fd8ed6e398265b90903c466f476068baf34275eef023ab30d95c909839c86c68cfc8cb4c8d32fb2721f7886e89f374f9e7a0213d0025ba6dffda2b87c0cd5e33ff07a2d0e179cb7a21f7ff81dcac2fb17bb526369f2845c2fc941624;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he5683156e2fc25ac30b71b58b7c2f2547b8488762ec712126aca47fa195425c0ce5f8de9f82c44dd2ded28f8aeee60ec9588b0225bf397f184fbe02994b77c875c7ad0d2dd1cc30ee6af238086e0346404cede5e412f69608c0d9bb44b5e45a405be7354f040e7ab3be35a2efa9eb17012e7111e441a5dc3f3ef53cca4ada2c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc92e8ef15efe07179121348bc3f0316bbf39ffa3df41b27373befa2416ab3957c9139ad80849a555f2dd278d93ba3a67749ccf96526c3e439cc2c257957f924daf591bdc383f1537a9b579f33783f5fa1fd9ba2a82ca77ca6997ef3cfcc783a3445e2333a37acc6bead8613b1b58b8b600b266a74f2f82e5c029819821c9d0ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8fe02f1f94c82c26f88f4ec02852ba589c868405b429d9d70dc40eaa4fc8d71f233df83b0eeafd364ee0f0c2d2eb61fdba7683acbe3af8116159918491d160147ca4a656988752f4e24c8f6d320b5daab5c560d7da2e924efd367a3a4e5ca77e7c41cf921645b5c641fcb9d6d7e9eac72edeaea7f4a090d32f8061c5a8eb6fce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0efbf410ad2c8c6a2265f7f159e55f45dd5659c04f8985dc0de87d1da0a1d3d023feb5d1e96514b2ae1286d6437325a56d8c74b689bc4a76f701542aae4ff780657fcba1db335a8ca55f0a294414993fcb5ddebadebfc9045fa9a026730830a7704de9ce2519a1ae894e239c98debe8396f8afeb008c04cfcd4acf90eb07b08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4596dde67d988adf7432090ec7dafbfd49d75fce2e9b078ffe8d99dbca6f0ea13601b2800fa0dc2ec06d7f00607c433ef59381b08b820ea3a030f6bdf576d327142f429e686a51d8c974df86405ba7c03b9253c6a7d158cfa26db996475fb7dc48966799d083c7e8f9ed47979839214d845bd076a4138796f27b7075760ebf7e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a53ebb71d92e1c72ca8b579206e74e3da8ae1c2f6eae7b6264c3e6ae42cf34868de3beef7d620ed7d65c04ee9f849579e2a7333ead8dca64b8c0b53c189b71e7b2e6794c801b22f68ab3daf45a41c5f02d409e6f0ef68ef2b5ca3ca4f14d0714513945724c5176ff22ad4fd9854c9ec117313d789419ef2772d2ec880c57e92;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1d847cb800a8aed414668afc748c5d89b86ecf2734d4eda11829d361fbec33991eacffb93ea9108fda51d2883a93b817f4bd31bbafed0aa1db0b38eae5f6b8ad0dba6bec1668ac4134057553453ca252c09112749fbe5e76d5ca304902d9a0b0abba56710795db8d1cba39b1032b72fcac69c0229be262129ae5681877f385f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h29e40e7eb7979efbd3cbbddeb256b11f2e21308c18c275f22aca3f5057d4df061c6da6f530a62560998ac4a64cfa10cb37870c9776054d091efb1f4f33efa6a8cb9c961c5214a52350a8c2ffc3e1f3538fb53215d7b7532bccaa92dd200d13d564f3fe084c73834b3595ec68b91dad3091a8f63a54aff7debffc16eeddd5df32;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbef4db623f1efc9838876bd03b39755268ffdda193848ecbb763d8b08972604ac3e7ba27a9fdf3b254d816c864c83f0bafb903a74acae3fa58def62a71459bc5f67aca63b442d38e57fd900881c9d961104ded14faf4acb6bdf06608cf150e670f81192fee6c6c67e0e1543b38458fa431b7c668e18ab8aec5af879d0599ab50;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e97d180800173f82c32ae7a53977cd68c62e847e42d8d3b4a31917d71b2e4318ae9dedb81678c12891f93d1b98b5845c2ec812c49d51fe4d7bc6fc187dba4fefc6b87b94afe842ea6354899d2e228792609e5923fb37f354dc0220a9703c7db6abec4182bcb5c8f70214839afaceed22dec6314ba7552537f7c0bea1729f0df;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4dac1b4cec2c0fa5a2300d0022847e250ad62f1de58a4dcc13b21c34b541f1dd4030a3befb51777d1cd6234b6b9b12a227b583e06fb8a9451aa37b36f1ac27e48dd7659609abc8bf6732e1efc2bdf19bbefc7cc151aa0351a80c9733e49e1fddcd1586bc5d1f547365af7c4e8270e5fa3ca0a9df9cc047734c280bba39beca1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h920d86a35cbc2d56bf2ca2789544025dae066c60c1f0c58746acabf1d2d12279a2d05a4dd3af32527cd4c5bd12ae97a4ee49adf75699fb969207945df04d2c28df9a85a313be827ef43655a25f44438b55793b95afb724b3d700c63c0e702aa1da45eed10c5cc8f57756a72eed13db613ed1af89633aa3475208f5214d8f39cd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he92a57ba514de8cab8025399a108ad4d6905a1ca2d2c15bd2b2f5e26df7a37ca6f4dea7cc573a0a60fbb7469a1ba76d9fae45b634ebf0b7ca989d8e4439f0839f1d3d7f845b1a58ff3c1973f8e85513c9d4dc6647c28d636ec51123eda5c82040d5524daff4928867530f4835bc740f762a7373b409e06dbfb76e79a08a2d6f6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d6af52f3af60ef38ebc85c85a263ea57fde7656a9b05c5959907caa1f7bd50baa887a2514460d628dde76acd2dbef557d1c5be2816894367a8dc390b61cb4f2476a60cc6de606bd789c02d9fe303b3d30ed16b408dc15995de44355d1aadd98dbd1d66039941908d70709748ae113191afc9011aa4acfce20feaf3ce3f5b097;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haeefe1ee40a420cda15e49441cef0e67ab3fc1d02f716b49c7a6fdb1453a2b4b8c22a4ae2cf7d5a02938f6a41ccb45b27dd1d196595ba57bce64f151968f403a8074d82c1b9caa1063b5191dd24278d8948fb6cd38aac0f14e020a412b3da3a6c1cfe74b3a913f6877d29542a0ecff8c5f5576452d230b1bbe0738f409e99c15;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d8eb709e683bfa9c2019704d3491cb607dd206157b43c45d347a6aabc28df43d1222e8eba24da5e8ba15bd67ec8b57512d80147f9f96fd861b7aefc566ab0e42fcc83baa6dbaee671fccdf0527b653e0df89709c04912ea5b6feba9d2bc066604e394fcec6a8ddf3f97e10bb2d5e889c4622925aed7f8be1660055ee74da9e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ee553f9f7c762e7e40d5f93796d6e224b230e2d760e983e1529fd63c2dec704ed06db116d5b37a27deae158f93ebd2400758637f28c27ecabab082a806fc62cf602ec9cc5286c320225cda68be431ab27bcb25060ca12a49491484cbe425e93b353646d755d8715cb6541223fa746d4ee07e46cb15ab14318ac6e5d6082a45c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he82d06da566e3b94f13f5c3aae009d51357639b5115c835f6d280d3a1a0654bbfef8b785d2e24648e6baffb6b30679344519710c4b16c9b3ebf11279be4620f270455fd7c97088ce78798c404c7e957f3f8bad015c5f9f6a3d3d76027687f16ed8e6722e9ffa71a87a5fd33a66447491f3bf6860f46cb0e0dfc297c4e2f34506;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40e9fc53e57083a819ff88ba4347456ecbb9a40594a7bc99436f620a8e6da47b24f321541016fb74c6219724e3fe68885def727cbd6701530c8322d2795530c39c2395892c2730661a926c2f61b60456ea9fa2f504da44fcfd9a9e53c0bdbb46e5f287a1ed224623c7a3d864af01c87b290c69737c5418626afd60f7949ff09e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a0315f0f3c95af1b661e4b51a4fa1ccab4cc345f78a91097810f2811c89f5722dbbe9bad5f01c887033b225f2867f1d22452640d53e8f3699e34fb9ee8cf0d0cfdf202e5ae6f8998cbf71df2111597df7fe8b73f55075b941f46fa7be7d1f8b97fe97a4e807a3701e9a135cc5446053a594958e045dcd302ba6c6d0ed8085e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81b6026f6d453583e1d6431dcde6e20746439e12c4da1d5fa145b5a603f2c3828a39b529eb438ee9c76bc115f2277acbefa0b3b2bbcac8fbbed726acc3588bdafda3a33cc17ed56827f1903ee1b29d30b528a3b2eefb7ce981b26c935e1d210128e21efd89fc4d03903d1737c24c3cf3a0c1fc4d9c08aaffb5a234dab49faf0c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb73689bbb7fedfb9b5d023af0e3bc0f498ab1e85643a75098d98e4a7430a234e2178aa7a74c1213d421e0840f557142252ddf45dc64c70e216b0695bcccd6bc3d94a35b02d536b303ba2f6a9f2a5657ab58229c9ca86a41d2553f4302c7a5abfefaa2e39555754284c488cd0032c7211419a4e17438b447d63a38687204426de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4b8e90b5105de7d183bbe21a1ac91797a653b8162fefb4a84670a713640864ff8f81348d2107e037aefb08cd897664dd6fc2ed21cc76205115f2d822fbbc91a582aff5ba310bc02875ee62891a0759a16cbb10e0d15964abe2215978772ba8a685e8ebb2dc5b06331d3972084e236b7360e6e5a885fead362777a58dc13090a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h149b1dd6a3c5381c05957e1b4bcfee27313bb8b649c7881e12f452bc2243d47bbfe19ccadb595651692c3f48ea8e6b5e2d6c1ad2f954a56c519420af3cc1a3ce21d0a6f5e2a10fc404922d49fd87f4ce517f7978f72288fe917e9fee797f4ee6fe79c50063beab32d975afe79fad0c416146bd2c0a83550806497cc17492c38d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he73d9d088f5b86569507367983295acceff3972cbcf9d5d804203c7733757475b79edb64444584e0024282c500673ea21ed6d0af90d43a815c2b459884769cdc41a91f3fa941cd0ea86e6af8b31b5ee3af6ca8d482b4b034b6eb8e80ffa67c26c179982f3c2f4fbf93bba4a24c961bddf76e6f59057a6f22f42c94c531f1ee08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haeebc5ef72bb7bca5d5bbc2ca86a81462cc5da710a0ec1900b1448a6ddbe673fbbc5703436edc0e3ea02f8a066697a4efdac3aafdea940b804fbccd87f05967a60715412593c6c54aa05aaa304957fd806a735b87e383f3631ae43206c9ff8d27b35c65a4a1d7afa1f164e05e3b0d27f7a2c24fde7a12cec5ad61d11a0b688f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28983619cbc32a74f68c53942ffc5837d77fb5c74854aef02f5e360ae8b03e34c62fd97b70168a7505fcc87f3c1abfd35f0ddfc8ead5965963a5f4d0d0873b35f17364b81fd241cc88b0a8bf2baaf12ef9f32c841c8e345aa0bc264dccf978e92f8bada23201942af0741f3094f5cf029ae9e4baaac2982e7a7d80625db5f3a8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f553bbb4ca4eff45966921552beeed45a5190ad529ad44179049d8a0b587c64760bbe00e834ab031c757b8f70362988aa9e522b6c3276bffccad9db4ca42e9900ea23c35e2b9a349bff0779244a5535e00e4ea93d978e0b8c26d91e0b6430ac6e77974be1ada239bf6c4008ae2edbcc0edba44548cb9f91422730282434a7c2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h546cc8218bee1137ab966bed87f97fa7a7e649e6e9295ea91cccf13471fbd45bdad128619c2e98eff9629b090aedc3e5e967c4fb2c830a749df53b55dbdeb074e16a6c5d000d90ebfad883abcf6b52642534121c616b8ead061b2a10163c4993e2301f9d720bb8bd1577ad06a390df156bd5873b81118d9fc272c79101aa90a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d3dc0bcf3f95703c496ad66cb79dd851bc2b6ceb5c839898b2201df1521aa75fc2c52a664452cc3ee46bc1a26d1f01c3d514ab43f19111bca3a4cf24457fdb710527f5f3c06f15d1b3491ef9955c82fa0390fb67d7464ccf555090935e2fbf8f2310060489ddc7ea43cf5c23938fabc1e6f5e502bb420159737de6d656c1171;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c9aad0facec22a107192dda003caeed63f0e7287cf80efac82afcc41af34d9614a9a662c26e08b575f1c4248f259aef4898cef098f81d3ae2f1c67286aaf1dfbe8daf830cec276d9299dcc5228a9d9f6d98590bd66e50dbac38c204d3e94da9c2257fe42588ffb1071fa07a607794621b7210202df409be3b04929d9e94d306;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1c5e0bdbb7b1a6c83a6e774b80f202c0b25f0ee453954159fa3294f7b5ee2ae553041a6fce9266cfbf6cd8b19f6b21b34f99d3f7f43475b0e752b4b84309e120e3616a49f083a6dd5ebd3e0ac935798e86cce37a7a47ae4a720167acb97b44981b7d3ed23789a7410ebe64188d8630f071096639bca2ae60cba1d84053906ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd23d00539b30ffd3b67cebc3c2a971c5ec70d2097d0edc875a988a4e1501b5c3197dc9b1a36c7d143c3778360c64f2621f3a420863ef276529331df9f13eb7932a60921d30fa797fb1d6377ad3c700b05699ea7585a71d18e8def50298b5037acfb5a6773531c691b01e5942b651e0c6e0910e4444a9e15096dcd0ec344f45c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf0167b7ad1f854605ec505e0f33a9664e93f340262f9d763c5b793fefa5f5f4c5280743a81b4afbc7bcdca5f83320d47c910057e51cc8f9c86b88688c608f010d9a59c22f00716609b2a8b51df5c51a436b9a39ab11730ba01dd9f04a44e5cea8dcaf2ac065e1499ca0bed6849ef4a975b2100ab593b4f776430fe1d6e726a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35804e48b839c088e21f027cc6a4a9280d80dc8ff6bfe3af5be55859d89d38a68ce8bcf48f4db6884063034e8e15e3d4d2e1de70cea998509847bc771aef76378f8915486a4bbd100b546039b063ce527e5dad39a8d82e5443813eeb13790f15dc34a820bd1b955e803d48d8de4d1d8506e5cefb51790f8a73caaa69c8c1d7c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d27fe15c67af1d1f924ce76c091e7b7fd014b80a94e4456ac39c05d4dfece4a46ef6d378d93d1caf2a0b341aedac67bec4bb614f8d5d9c4695488c58d1fdc785e6fe38d6d4b66d99212dd0c83bd65904041b8f25da191abb8d50cd45dc8f05c4c1ed50f28b3f7e1c6ceaba0fad14e50d1f1e25f77c0da941bab3c827761ef8c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hebf5533de7f9834c64d9794525c582009712426cf5daeb7ca4ed62c5a0eddb758f17d264460ec24c485b2f9118f9ce2fa4b9d75fdbbc012ae378f114f4b36edec47deaa9edf2f0fde09f5809f83385d6d6172f1a5fe2970be03b0617eda3f5edb42e1294ff5dd6adc2960baa954f222739b948534d3726c81e8be68af914e65d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb22e5d2c9729d2585f956b786b60ea3699d84b8621c4fc11b8b52078f4c263ae9f288d8c046f8f83b760c2ab9e58131fc0879a0ebed3ecb41be2bb57e42736e19a7dbc5b1589b3a2707c0ff4266259fae0cce01e34a748a3ef92f92ffa5f8f2e7e811a1ce87dd9fce4e80652dc50299d674762efe35bf5abe9a2a7f4027c554;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb074f3215df02f80cedba4de7c5cebc6ea4c9975723e53002b1e36692f3c1b1d628a8bb887d9f0334f5947f7e4106e714bec0b130f0644b0db5730dcb0b3c8f49f5033a9dd90daab63f7136b0f0813c06c7c9aa5e097859503b880e504a9a40c3aeb338452ff87771b8fa83991e6392411ecf7b3e24ce8fb60b9f4e536a0cb46;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5cc58e088817a168ff6182616256f44b94eac80f31ae57e9970b597e12e0f3c833e00cb464fabedcb13b3409b73ece5ba19c360d35b98da212adaf515f7397d7bdea9e597fd6e88dc1ebb1b27f80ef5f11e7fac387ef549bd57293413e0c1f5e2f0f74529ae89531d170fb1b235c1e3c022541522d83ded13937fb04c91e36e7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7611e010914e0c313a619078bf592c2fdec9d3bd939221a978310c3fd4251716bd67c30d4fa5612da91ed9f678b0086a047a433a86271b74624628cf3bfb02a08bf7b46cb5d9ad43ef2de189f4a2fe54f34929a4f08e4bf3178e68869cb858a980e3b1345e1a7bebf12a1ef99d4daa7e017f010d9b0d3f7d8abee96c99a6b426;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he257bb48ea3d18834414eae11e92f889a465c2042856fa9c1cb3ccd2240a324a982418a39653b6b46b954b4351b9ae74f3719a334487b2b2c7b726a5da18b938c806f4c10b40225d181a0b30754429edc9c15059f2da1e4116611ebecfae49d63e0b679651adf24bbb6d0cd696e400bec8c4a9c18d26e10d41a75eb6cbdaad46;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6a094e7c3a35b5752d99b6b44acf7e91971e542f5e8b758d2fd2a61c4dcd1d7f76a146cda3fa8a6a45523dd42283f7bf882755273aa15662b73108fd368d3333a7796ddd1269b83b09141441e7bb77bebd9c6d70723bc50104c3cd585fb7ba1a762a902c3a2e7f0fd2546c7ef9c1918821e2412d0f8e25282697176170aa100;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e6e7b9418f8ce710051b4b57fd3c9fefc83809b97488b56a7b7acca7118db7e5e14ad34291ddec1b208f28c5ad7fb9c2cdbb35ff0a3c7d83b77d118677bb3e03a343c03cdd93a357e79c071d1d6a5d8dc038af6e655b01dc693527d5598f7a394fc557eabcdbeaefed23dfc247ec49899d62bd78fc48cebc3a263f9e29ffe25;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbfb6167a37a10c799210b925041f063076dca40b91018cddef251ecf87f5873ca86d073a43a5294176aa6a2e5adfdc26d8e003c2d841892f8f0698923c2ad426625a13da17cd74f635904a20af549970da7cd9b677143dee3b82047952ab0f65a860784355e5eeeec7b06d2aaca2efb1ea0a727ea5556b64926670b5189f531d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26b7dbb02fce7094f9bc80deeae9df99f968c4ac4cdac5b4cb9490dd1a1fbf3e089bd8b24c650fa617999a3f5641e91c71f22b656c45510e0c2fb5b9f9fb99d0d4225c102b4d7c240e8fc7efcc8bddd7b4ebf34dcc8a9194525f141af51a499b36e45bfb29c05a126a2cfccd1b0faa2a0344e7a3f5750560468fa242b9cc9037;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38ae13dd1121fb8e5b5f43ed9a1a18664ba685fb0bd97eb8889e4ae185347d52379251760e29d356e684259f62b63cfe123ec4ab5fe41f6132b6ba10171417d67e5aad0105dbcf56a14d8773d52a4672577d40bbb7b767a7c442a6c27f2bcaa1bdcde19943bb3ce358eb277a88dfa84d3662b9bfda38100886e04ba49c0f9282;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b4a9002ad2ca7cb3831a3e95a0593de2ef3d2675b82f21ec7250fd92b92305ab683f886f5b0a19bca6a4d419e600fd5834a7fcf4f3f07cd4c9cb9088a020e50cf12ad26418bdea246e1096b62e4834147acc7db8c9abd010fbe5c1c6be453f19f5497253e0dc4edec5e054186c73028bf73b68a8a3543c253e06ddebdf3e062;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb24e0a3ab03d1a2949c715da77f0f20a9f513b38b16e76768035fd2f289e446f51ad801f623bf0151ec363f8f16610eb4a2df9c20a2c7148cd99dd954aa17a45f89fd5d4dbdfd78a2526488ba7659c5b1ba8c558d8f3d0876da2a5ac8edfc2c78386290d1122bb3541d67acf98457a084563cddf95dec4c1ca5cb86978d68863;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2ba3af58e9b46a1feb8de972148f3527584e93e6a70fbaa609b2df7fd44b1dcf8503b20600275fe50052fafbf8a18d083a6fc5771d9d377c5f594399011d6876d091754ca3a079a839288a10f54ccdd04dd8c07dfceb172631b67ac4e107fdd3fab8bb962aef80c18a445539bb13780f7d69e1dc0bebe2c16fab292c2714d6e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81519ff66cd471571b9c5e5142195f83ea305490d1258a9c562748d5092631de2b589ff60d03c2ee6e0a8b127ac55e578fec927d97bcf12a0c5f4fbee05fa2356d7382619b8462aa941bbfd6ff62254953a2517f9bbf95663050a2d201c808177a7e92cdf3355445aea883eae678bf559b50f80fa539566ad9615f6baebf8600;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43e29101fcfd84d5bfcd2ddaf12e8191863b830296f33c5d89255ad3d70e9567c7d3c084459bbe276703c60a7820dee97af1cce05d1d6325a2cb0c6022f8f13fe8453f40a6fe64997f99e114564124bf363f99e785949f043c0c18d76e7e45c35333151ce598b18ff71aac12a6ec1ae39ff0c1f3340533d208898aa11f23871b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5388d68c23f5640d4c4aec45ae396f86cc10dadc6690cb34da34f119c19b982e16fcf3eb204739ced0083362b65a39f95d4fe7d3a08c1fab030b7cd1ca1b88242d3e671bd08a597cc446eb0cf127d0a739c360c71c92ee61f480a9f9a2094fc1932c72b60cb8f3a8b68042d86329750ea1a0926fd3de37768d12cf43ed74bd98;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2b15eeebc22ceafb1ebf5ec11d29ccd27f2c53b902129aeab07f68bfe7ae4938cf71773ea8790907b0f570bbd2d83d6743ed327a13da6cd0ed2ba18e761baf75c47ec767c8de8ddb002fb32f1b4a703de58d2d991852b9cdae4f43f1dc4bbd6a5bae1c24ac3285519cd3245bcd8b863ded97a07c6e51c257cd3abf073486ca3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4563e42775b5341415284fde7ac25e77a0bcbf3895a429470e8ea91f588badb190ebbbb561a25f9d4990526ee0222d2ab9107f331ee885c7b982ea75a2364b5dbd0a4162d4e8a0c06bb40e606358ec9972ee6fd7a2a2c74083868e0590196b219e7252d7a035c7a70b43b88f833109e6902a9c9ab5d619753028f63162232e12;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27a3ba63ffb4413123b06e229da6d7b9b0adb6435695fe36dde9d328df2091d129e78d25a7bb49fcb4c5ba9403dcf0b1c624964cd018e95507b1c1536d960302210c3930d69b35a4d9ecccbc80f4fbe8decef154b87cbbcbbe456b5af3b39e4e5466a931023296b638e197b08688e224145428fd33b6a180c28654b3de5af5a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h99df6ffc2c143e713b8d30b0c28902110afac5987d7a6300bc90f627263c312b78f3ecd420a15394d13604bc7526146ddd3b678812fb2cfce09f681576107b5bc9e73f655880f4fa237decdfdfb069ec6521fa2d97268c69e5643c0957dd7b0b6b91d8db94cce018af373b8fcd789db4ec2a4bfb4ce778e38739f1290bca20ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he6c464a7937f609836498815022d14242fb29d066a051229d62eda07106b3c3017366b0a586776ae274f26c7a91246b142f1570f2acc21e3d5862d0dd4536ed5051fa1c48790839eb449ddfe874b1020dc636dbd1b6183c5a6b4d4f5ead402b9158b4c04b0652a1b6a550f856c364d7ad2d83fa172d1ad572732bdefbcba0d1c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a4444768be976e6addd73c2824aad1f330784a96a97c049b7499bb1dcc3ca0e5fda642b6bde282b4cb71963c8ac6cdb31fa8591f33b80965e53b927c2ebf7ae551bf7b472455fda0dfb6df8d0030e2b4a9586cc9c087452fdc91a949229b6db6512d36d06415433d99f44238c90e82c42e46bae5cb07cc15e040664bb7cebcf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b86e6f063715ecceece4dd761fe56f68703e130d067c4a6545c408d4711c664749a8847d32270fc9b4dc762c8f59febb3c8a167153d6d7aba5f6fe44bc411171e82c977c24b18c4046f97ba5dd7f7926e73a32d91c4cb633560680f53f5bab4a4f6c92144e2e400f4b0468ec959d7c86955acc169743b211a8b82c35d010d7b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc32b4f3e83928510f7c4bdf3e5cd0e8d68c79cdf5027903a8a7d1b0d7f753c32e5afa4f85d7cee90ce548653574df52423f09bd5f8b78e8dbd6fe958c92dd413647d2d1dc704745733e1601c1ac987509ef67202ce6b83798fbf03d1a5764c5156094bc2f9510002a9e17d15c108c7d0d228020e72460debd68bbbf10c43b0ba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3d24fe80ba549dd025add3db75c91e3482bc45ff35aa0316669c59a2faa7c0822edf9f62b4c61b3ba9b3cd81e7cfdffcf8af09f608918b59c79463cee43dd20f2ca15c63a7b59ffac020d9c89e46c76942a403223981e46191c4dba71e75ce556bb43760519be52b7844d1ca7df1b68405703035d93ad0046dd0408e159f12e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e989ddcc01947fc9b316cbc6f86b0c02d3e1ca9f76ad4bccd6a88740d1083afbff112c9f002a6a43443f06b2dca7de82c0c9494daa4b8de02207a3ef24be99b9f2434c998261cc49d6a673bf123e314d12282013d477efd841ec4a20c9f3f6d91197215c57e49e4b999eb071283ef13fda5a3503bbc96cbb8064002b72fa85c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h965b49667cf652b4055ea9c6cc6644e0763ade470c062a42380b469736f134177a04a5a8daa48150b4dcb2691d7e12cb1d2a66b7ce0584b8288d51d9c05bc70091662c7b2548cbf8a5cd5017b84541a8a59bae490505cbfa837ff41480ae9e949f653640cb0fddf77b1a6b902d5820038e2553ee0d8cc4da9438384308281247;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc66998fc4cb3631010f8a8790f61fcb9445abd1e4d681919c407f7166df2fde520d7fa4cd80a943fea35c74955b57af91e8d57b7d6131cfdcf061d50bc6002501a650f8dbe48f8901246d1922901d991cac7d85d6e5efa810f44dc14fe22c30cc1ea8683c45d47990028b7f6041a22f6def4f3ee052da030d11fdd6533274e87;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1f6a6a4c2cbc3fcb8192325e55e08d525c981f07c28e84813411b151091b6daca5e860754b1f049f2683ecb915a651ed223a22248c551f53bccc10115ee159f2d6b642b533ab715c3cc8827943ff2bc218ea54e2379d12fd226c9f95aca6411289ba1606e567333a86f3deebf6fae4b129d0ab5adc3222db8f145d4111659e76;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd45550f67db524d83ed688d97a32c930bf89fc1a1b7c2454aa7b36a55d29d06884204af460582a98fcb19a2b2cdfd2e86af41bd56bcbb292dfebb5dbf966604fdaa5540147ccc900bad2302c7074a493d79ba3bdd24f628f8405ddf2b34e20ad58337303914f86b3ea55b2d2e0d94811715707e94020f0adce779047925f264a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca7f37c1beed16a502e91e0728f86153ec928c5eee2f2ff6bc2d676ad1614ef1925b6368a1af0982075f76bd877d6f49622db83c7fd0bb2e7b154cd957c341b5ccb8da181508adcb55cd1e8777ccd9c3caf6ba3bafafd008a2f1dbf725c887c1a1781ffe494212bfaa7ca321ffa6883bc1935fcbf5b63dc726e9672a0d3eed1d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f70719a82136c7bca35d101aa0e5dd65c02b53dadc6d86d74bc38292e1851cebfd96f4a4aa2be47f7b8b11f2d92705246b32e2792410bcec93b9ff2cc62fb6371e33760f6926680ec581399d3e3acee07bd946c621200647cdb17eb6c6a5f76dba4fe4f2c4948c6ae1f6ba936a526d58835abdbb5c7eeebfdffb76ae4479f38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h214a9cf129af8706ba9c05dd8bc820b60d0cf86dc580331d9a997d9a2824d26cf5c8984bc5111bd118458e4b94ed953bceb5266da106a566a618bd93ad0732f7e66e6a054282a083fdedcd93f6f36887e46c97ed0aaa5403ad6ee801aea4c482f678076ac8cae02d73b184423875c0b467bb0f50330f9998171ae76b59fba2c1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e684138d5ce16c4c98dce3e413c34580bd8c2ff5ce2ec9551876068b534cf32d46dacffbd29695b0ec0509688379d6c875b402622a4f153c4940f03f48cdc01c43a111234f3cf327d2990cc6bc558a2c040455828da93647033d8efc3de27e257e972de015ca016de0a7d656364c4bd686f806ac56188c1940f619df0d20066;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea3ead813db34e69022df1360eaff100fba68d6f7b74e33dea872b54a9418dd41a7537efdb5565218b84302d86a96bce56730a5f0cfdc7debf1dcb2236aa323ecd7bb047c9df3af564214980780422e087160c0364af902585c5e32bdb6504df2cccd53689969b32e24bc1d39eb0d18ad0886c5bb3b61a276a6f7ed7ccf71319;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h930f075a33d97963586b07dface9c395e158e55f96b08927596ef62a8f09d25a13d0c12eef7f348b1a0b6b0f635b16c0c1d1119e40936352830d3d5e9f9b2a9b80cbb87ae0b53cf11e04d49c066207c88090a5078a8ac6bd4842432b03e97610b0dbe61e8e46cde4ae785d396f5cd5f679a78f7401ccefa99d23d1dc646c0e7d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha383ab63b690712a48a5ec4e8314e801d6c0b030215f38b708012510a8bd0ea687adfbd49bbcdec4c685affc17dea87eab08ea0e3bbd90f8f613dd5088f6795abaecac22de3a06a53776cc66bd9e1c8d7b816d16b51d56211d567aa00aa6a4610a15ae0eb132491ebd8a1efe5139dadf326f3cdedfe43ede5bb4c21d6bdaab28;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hacca3b7949cf67b53e16624da84495aa4cde3d21dec170fa455ebd25d167ad3e72b949e4b4bed5b8b20e85b807460f17d675d05acbefdde0d3fa214d9acbedd4abc620299d873b689b59da3301fbf0bb5707cc06a1f11714d54da59d2045140eece6a52626d09857b51c699ff114de97faf55d8898fa5674ca7c2e0c8a2e5dea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d4f6e108e5d89ca1770a455b2934e758c6701116d601065bc5aecc09631a4a15b77b2929519bca2a38941104cd1fb59d7754eeda44acb10b54e28b9675b0e727991c19c34dbb3c27a0bfda03c67bc370c1041c024b4c38296b83a4a15657fb1b6de6bfbb0b8358315a27fefcc95352785958bce3bcb4bd3f4811a8fcf86b6d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12d4a2242ea67824e6a59e86fe00a683d04dcbbcd34e90051f08e9157fd5e340c88e69bf99cb81f036c31a790feacbfa3fba345e8f3059a840402584092a2601308c011c2f97ffff7c50ab1100bf5cb828a6929161bc13b055667eb98b723cdad04317d43dd224b05aeccc20f269782758f5d2107882678f88f3f5763b980438;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45996175355eb0ffea983bdf84e2ed39f11b40ee38181d179642645d46f94be4b5ddc1da7069d4f0ba4bbaa0381b2b8b87e0d1f6b02924e27b0269628e514248a8f9666af3322d2fbe25e369ebdc5cc81ab29275e75174ddaef11d13e376c511cd33c97137c1d53b6fba653924eef807a5d2fa996fe19a5ee12821c67678661c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h555af723fe12633a22c9e30c55ef9dd924079f48b237af70fd13571192dedf9967801ba6706e09c01e694082f5086b503891cb605bb57156e07cd2a174abcde79f9afff49b86465973d65e57b9e152bb3c097a56e9bdf53d85d03ebd2704dc9384dee59c23e629d5ce857c21ebd83f34afb3b7c77426e452691d01bd90151ed9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc299a417f000863d04b875d8e5d133dd41249d9c220072e583af41d2ac315dac99c19770d7b699d25ef8473f16545a30dc9893d158361874b60b35023f241757c2707075a615296684f2408f96f4ab5e3b154c744a5e1713a7e09de94d5b22437589703b80a93504143fc21e4c194fb5717767a03ca8bde1f76ee599f7a0f752;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50db3fc9546de5e53b68bea368cd4333362bbee6fbd1d6085491ed989080d132bc74c192ea163437cbb619acd3835bea25c4fb62bb58ebae226b4e4702f1ab847fe1564a274e57c43708a344a8c4046cdc0aefc6a1f0e2c8ae9d8ba2dc591f1b5116e5f4d05a6b08ff9c874f37b5354fe4ef453995d3c12ccc0f1ebc51ed2e5f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb924dc39036f6c6043d8c458a4e8a9c65bb6cff97120035159d31da168e12947285d0849b5261204e7e7ad184af05d114116f361031ea2fd35e00768232111e008c1deeb3968c036f878151f127e71044cc9cdbb7f27d69422617fb8d484f73ebe03ac78bdf1c4cb139ae4d7d65d5afb1a06f3c2e0e88370f39729f10938f1c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h273cfb5ff92b4357024ac6824c0e97f8ec2a92b4ed8fb31b5cdcc850f0b7496c61561d2e97a3aaff64dd5669757d1b57ff9c99a6cc2b8ef9c1e815d693cc2ff903af8320134430d22e7e3288bf23735c00f022d1a8798a845319c102d4fb65a11fcfbf6b96de6a658c131bb88a2304061d8616325597fbd001bcd14a232b4a3f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec87bfaa93567098fc19413134e7464c0522319cb0261a14f386a6bdcbf99d065fc63e46fef4ba96d5af563dd622a1ea1f09ce072139eadcf3f0f212c52d37f1f21c23ceadd7b33930f9dd2c093ced03a9381ba7d8b7f7d0768c659f7458c27f92c06cf3592ea0690cbfc835371e8a10ebf0975dec0886e9ec6d77b30fdf46c2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6dad9dc3da871266ba9873abd997457e52f1d504c173c52f0e30f515dffa53c137f6aa34e71a0f262dfe3714a2c5b33c121a84efc31bc3609653dd3ff33d805c4abc23afe29a68b2b542b5ccad6ae4df3d21fa6267a06ccfc6f8ab58b7c38e213cda23e1f0621b5541afba9d66372de435de6b50b2a55ff6656139ef82feb5ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2705d3ad3d9982148d1f88a0642e893dfe4c541314c1c5e126524fc92572273612777456304429e856469ea8f5138f3e596093af2ccbe2d16f8db53cecc6da3fe8cd09317a15de59cb56efc4d6ce32e46c4daeb582c878b1c87f7b7f906011e7123ddbecd8067562aade58f41dc3df0e37f6660577124c921feabcf3d64f2358;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha48b655e659caf123dc0133497d50a98a9756c150a559490023e54176314f44f1911d4a8d58ae49dc3fe5c69b7a73c22966cccd6bd1a17dc9839fe033c92f513147b983d771398709f6bc8fc8bf68dc41e436c91cf24614fc6a50df5b66120e779ec35ff88e7c039094062cceb7ec4d0e5e66b0ccafd12c3b8f67ade01488a15;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3439ee1a1a837d6538b6c8644a794f7f8686e5dca78e445806ceafb6ef164a15a5b7567a0da39818b8acb989d258c7b5156ea9caf9a44dddd8c7a888e18e7fe5140d5a6750567bffd5f496a6823e9fbd2b6406df61e1a70d88146121d1c810016785af9fd64c93d8fdb74d9a757668e483022641c1f1545c15fed4bd4d098ac3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h755b0e80a1dc5f6e4318b7c2c72a88cee1d1a8aaacf615b5f325e4dd7a2eb09c6c5f3ac42955e4a083ed3bda06c8cd1d4563eddf5704a079e77345f38b9a324d776232402dec3844db0b14ec4e05ba0fd88f2f77c60f4bb11da30eb14e72016c1694bfa532bc2d2c71c7298847f311e42b6ddffd2e087089bb089289a7b72245;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf057e1370c4f46cd5532a113cd6cb8b6d02368bdd76c3e7aa5fc255adba9a6e39a5126baeab935bf92999521e16b64d2db3fc5272f704717c5ff78a30a14c01bb417f6a22dff815f080b49a12d51bdebf3c58d78a3c3cba7ba280c1ef2bb4c63b67a598f309c0ea8f1b8ba5cd80717189169beeff1c7ca203c7ddf34ee7649c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1777718443d95363bb77ba94cb2f9890f38f660d1795f23b23b1f83d49e012af8dab1be387a4b550918a7d672ea994a407a200061bad8252c7864395bc8b44171f265d729f90e23ea1eefe3a102aac332347e6f4f29dc487163ea6f4c381b04ddb6e5f614a5f4904e610239c61263c5c321d24799fa285a78377e1bfc56be103;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e96cc3c2f97b6db2457933ed147f9c9d3452422b1f94ca2eebcf19de6d1baba6db2d113146a13d7cd5da2a4a2bafced6afa78fa95e7f0cce94b4179f123d991c688f2555d9a05ed291972413e19a6677ded42023caf1b7576f70d93098873cda46a589670c45fea6a7bdeb65672d8cc81e67974a67e050802e2223b8b837fb5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c0d8ff5ebd6a4f638337656b16ff4f7369c55aad152663c8396bc231b9e3999a36586c92ea664695a054a660fd6c3e15a593eb406609536fbfb38b25c78ed3893ea630b466d0c4960d8126fe4caca29d4425624ebc2c54f8fbb4f6f9270f418a9dae5b28ae861d65e14cb266b1ed7cc36438de8740a8dc84cf925100351b04e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b50c48f85d36a3fa8ce9ff7d81f000b3656b05bf9f8df7cfe7e83caeb025da03b5cabf20b91134282e53f59cbb77852a599443dea6982bf7ba9211cb7a5e2750a8bdfa42aba26c8207e8615f7cf8dc67c26d6f6a80843e15b525a5186fb09852046bf1db73c0355af1d005229f3e3ca2a7af427881ce9c0837065183979d420;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf36529ecc4eee01fa736638109f29dd20de166964cec8142b406d08338249d249ab1b997121c46056c6332f08f8c3d86d967e5ecc78c4224353859498d25957836cbade6dc9002d8a4081cc611f049c8cd0a8ea9bf0d16238f616f191568165dc0d4d1cf2f1050aa93c6ca25a809158b6b01e3b7cef467e23f584c2f51af33b8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbcd341de976c7e5249d3b01398904f0d727b5ffc361491545d878281ae5f33be1503f0c6398500ab9d3e76e0d5eb5c99b697943e7b6653db0b55dde7756cf5c01812836a7f2717c87a72a7745bbf6b8c09e9019925102a94f558e5c0268696c2d91c458ee2442490e60931acceb2739e512ce75c65a3d7142762a3d8ebbb6cf8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21a1b4a35bb23a9de6af7eb6a203651f70806cf499c9879dc331ade91545a0b55b2dd19a4cca9254603a483d29d2faac8522d3df9700a1994da99bd80dd74979341f3c48341c1aa3009eaa6f553b06904d03f56721bb87b29b0fdb9f84cad811a36b45cb85a0c54cd2bdf633fe68c824b7684c5217ebb93b255a58fc1c636a4a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc927bdf9032b40762ce6ff8f1bb341826b6503327809f2726d7ce71f455077388d4210cb7f562391e6adab64d09433a47af6da9f9d9ad3f908a5a22182581182ff72bdee117432fa83a73e86fded9b6980826ad187705429328a5fd656a9bd70c8a9b72f38453b89455b50b83b5587039785a08b2b8cf8abbb7d791a1bd19b45;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11147f97b7beea9702aa8ad05d0b293d8080e7de4aa35856f1d1ea9c8b6d57305f12c986177cc2910ddd48c5453f6efc4e13b29d463d85e51df8a8590afeaff0a9ed1a74e3caa2cb03eff483c811074fd70097447d6197b228e1160c9f38b4f14e3f3492090047a3308264996192384f0dd7d46e5b3670a5c871cb92a0ffef15;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1bce83af5a700b6b867db6f63ae53eeba4382402a3466188763dd2cc9978e0c0653e7870885f1b57af17e52ab8e7527619fadc3b18ba4dfeb9f5600c8cb98a3a4c8a81a2d9d6f10d58ee328368e2282cffb3dc866d2b54c61e4323f83d33dff5fdd0eee3a2bf293dac1e91bc1dfb4db7c37d3610587514c962d874643f128a1d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6094871cba6ca3b792e60ec451fa6da1691a85a7ea6764da6d4581c3af1afb441ac2d51f9732ccea7ba60d60b7440b2d4127e7a8da49acd00c7cdd6abd0c7d5e03a03386c6f7d659c609284155a0a5830a7e26df4f6e142814b3643a17c0b72ea9eda48178f161e058a04c5869657e906a2b7a48f84c4484be2021eff4db6940;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20e5d74c02e78e17947419a36d02964ebde49ecbf2768d357c9e108464f2848c7f4e609f4daf404897de46b6a5290e534a8a909b65ac18da25ef96f555f143f69d8133060b58dac1262572285cbf8641bc8ab8322479b0c1b118f9619971cafd73f5ed61a6e6f95d6054a380bf6da876fcc17e12d0e38829bbb02f89e925a15;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he88e5c4f111a236ef82f28f653cb46330b89bdadc530d6448ce6823f82985a535f0c740ce9cb725a515861f224722b7712eb734ebea52e198041926dedd164156032af102d225b48c01c7b942cf4f99f70afe346de75a8465213212a76162132ee787612935356eaf10e36f4082ab1eb157a9abfc2154b71d1da4c8b0fbcabca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h577370a4e02f9e99e9e8a925fa41e880d4d9e8eb141f8ebc3d0a4c7a5ec49df1765767ea6b45e5dfa7b6d44fd0846ba60f2a7c9ae0921f236551173a2bcbe80ef86bfb1d6527a513560337c4ba318149578a6543a0e3ac76d4ed4b77374ca3fc33451d4fa6e2e3cd88c8bb617af664723d7169ba8cee7f1bab78c06b93ee2be6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha045c0806785d9fcf4a1ed1cca6e4d15ea3b426d013d79b8e271f38e4b4f9812588342b6d42d1e345d8c93b0ada60e7431ec7c89e7c3045e55ba3f5a3e911f2ae496bf17d8f6c45cf8363ef2ce3d438332f72fb021155d161aa3a1c0d2e01ac0a4a6de15e6d2dab70a31d5baed25e1d4fdcbbdf5edbde5cdfd5bf2053bdc60f3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h92e4703adfc91a0f68b41c8371fd8b67f1db228add8084a6c884b6c26db6afa7b9f63271fa6ef58840df9809912a42c8aa7b410b7e9a72d9c133e2edf447a7915e77a1ffb8ed3eabf123e7c24f63331b1b95fdc6a0036815fe3a1b49be639b8676bfcd9fa97f465e31c65b9566b016dd924bf0d2f67f4e026340c55fc26f5efd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71cfedae5a2051e49656066d0f6faadd90da677e807d99d2ba9263dfeddb94b7fd60c5245f971e32f6af3beafe77f81c6ee62386c62afbd7031acd1408eb3eb3435a4a89e3121d2a6b64600f90d2cb20a0a2ecb6de293b9154f13f5f3a7503b2459f0e4651755747166e66f4c657e3f5d666accfcd2ad6f3813152ba5b48ec2e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h981b834bbec1de76230c1bca331d37dda6fe9274e550d67e3a784a2ae39a22aa0500f0356ea80ce9a57441548ae4ac44d1793314b387c2c1dc53a19343d2839ea236e69911a72b8dad6679c1f998290b83d6b486ce8305e581fa5b7c96dc391107684cc02f5dcf48ee5a44265dc9f23bcafa607806c182b696c063ca2d8f9abe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d182642b568e804f900b3c56383be2c026897f2c4f85e73a1f5b172f7253a00d3b87905458dce44f170d4811d9601ede41eedcf0347a99c7bacc343c88248f7c17ef9d1c7bb65572ab604f969833f4d3b5e8bb06a1b35b23982dbe45ad6106f6d8a39d398642f16de691f17b77eb55b47e1e82b3a1bb986ee8bf1a3ece1430d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he80e09b0eee5ee6c8a1595ec32011a5eba00336a7aa20ce9dd98bd3cdba7030e2641dc5a3436263469644dcea0efab8db31a9a22e5361530cac8a69c21dc48a55c511d0453e4ab33082b3bb13c5467bb92d82b132721ad4dcef7db4276a40246d69b6b8e2e766234bd4d888e6a1d5f8f83a2d35f438f06d35fa6ad582736eb20;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h126734911443ee3fa64101f0f4bb3bfafa1a0dbc987f3248ab58bada39cefe951a5ad71140c72c59fbeee4e1b42ac4044fa56183af3aeeb9506039a7df58aaf9952f945f63d18341697999bd1d077f0b0b18e49059d2d96f09af46e102b926f9a883478b0e17c95836c778afa378c1ed75b5fa0e8f4951c86730fe77561072c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbec26becd1437851180bdc4f3546107105967beae79fad12cc2fb6ea904e4d59883ca6cbcccdfe65fd289a74e90f9f3e25ca0db7fe84b59db807fd6819582e1beb76a6a72eee3637146e0b8e548cdc02b3505cc6e3e1985c8920251a39ea744aa9bf4d784acd51d1d3ed43d7a18019c113500ce4659bfaadb94a9c973447201;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4062b2f4ce07dd141bc9f767d9eca842f1641d1b2ac98d743174a844201d0368a0f8ee67ed3576a1b4bfa130c235c8a1fbc38d2a7bda055a565ae3612f80653105b6f25f77a4441a39cdccf1aedf621d6e6096e3a5f6469c8ae9e64cb5b6b74a90612ce2ad808a61cad244eaeaeab09092dd6f27fa1438db50cd1edbb42356;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h720876ff4865113da3a7b82525156384bfefa2ea0de4c4d141994c4024f003ed121c63a7470bef780935d3f612ac1e68e5c3366300d7dd8fda1cc5a1582e2ecddc0d8b4feef52ede21ce647974af495392b21c4d1ada332aefdc7cd385913bb24405687ec410e46fa4bea5a72b65647dfb985a76075eb5d2ba6ba80e5979412c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d998c9bced1ca1e92a85d3d8f45c7a679632dc8b74a6b1ea9029dd5f06a4abade3a493916903d31505bbfe5f0a6c58a9325b8229281e9282976c1bb746a3f983c74e085d5abe2c6929bd3fd15cce4740b7249873473d6fc3f51b368f8987a3471311cb61ec385bb7e0287147724d43bc70777bf35f86c30a738aaef2e436188;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae64631523f319c2b7f6a5e807dbdd04bf0173621b1d78b13a1fdadf4a00da510d33c4094b444e38c9459872f86b772e200c84719777d16a5182ec1a7eac8335b46751c3c45a35db73cb47adcd4a0fd2eb4ab2b3ce017266ae040aca0296c6bd423e8d08017ca0984b275a04b7609865aace131270d5d847b6c8b6b7ae1c10e4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h76e7b42d766bd80a6283164e958110ae5f6b01579def94f61f1277b82b8ef3f930447595c7f8c1acbf28493407f1c49866922bd18276a238009b56e7bcbf4ce9c898dfb95395ee27082951b687b97dbc88362ffda517742e9c2ee10558ec528dc37121e87ce2aebc35adbeae7b3749cd29721bd99bc1ac1711d648d227265b27;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95b3c33a6cfa1c4eff493dfc4a43e96a238446885ebb1e0a8fcbe2eab29d78159c97593e431f6b44c58ae9686828807933ea77cca09ef3faed86ecd8939d15e1a8f154e7a311d3364da7e6b3df592c7a9facd8991429cb660138a067a479108fddbe0749eeac1a8da390169229ab37a2fdedc88a877cc1e874429f57b6693d9e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69f80941b568ece42e48ce40fde7067d4472ebf8be21bcc14d0d1c69f1a7b3b85c1952e33a14a460313f3f3ee8508f87b252c846e51d780eeb0b2a73c704643966ae327b2585ef9721ec554379e82811415a7ec6219425e5d0ffc6302a1a231fe73d3c06fbe2361acdf5667e803ee76336717f3b7642e30fbe3ee4fc703a3778;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72ecf1ec1de921d8f37cbd3622c63e5503480513b9ae764b37d409d05ba4a938abc8234d88ffe3a2800568164526986b4e5828993eadd576b34cef7d6612b0fed78e182404903fa115dda61259e478f9d155d505d6bdb1f895a0324fae846ecd3ebbe1647e99884456a4636e7d00aafac21a865d777f987fc206520ab32d5466;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heff1d06be018e6dd39caa600b528a9d57c0cb1925d4794385807044ca684dc3744985aa5781adec94acc88d99b35d82f428b099a00fac9e8840758655cd9dbbd9301d88b0a08330cbf70bea842304fbe00b2a4a8917d13f4a8d00f89c8dd3a9fda70955158372add9f31ac71895d00ea4f821f1e061cdd66d18b58bf472872a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32daa9ecc8ded14ebaed77acb27452516e6461b004f3223a9acebb3e1b855713bc1c1299bd50e08e7999cafd0478f201241f0a41137d9e8033b4d6ef6aa41c97c3a08e3d2aaa16f910380ef6b18b870a084800fc9c7293ebee0035cb817f3ac91a6bc52ae2e8810cf56b3014b5595983392939793751eb6db41f36e2cc294e25;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca8822a20e98c00e1b8c51d662204e89161fb8366718170478dda36c3eddc4e59cf8ecb7a2b930480e8a99d27c5384c7bdee44e3339248509f067f573a44f47ff95c8218b6c9652e3f4acd8add1cefcf04f5fdadd3565b998afef3edddd87a15af3d24cb5f5fae108bcbd5403e217e5b7b3a2723987001d2ebca9b38d1e5050f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h14c849d1c8efb191fb27fe5a307e076637554cbb6b074f67ca0944326cfe3fad70e517e95d37c89b78dbda2bdad34112963dd7479e7b662207ffaf46dcf41fea36262e0ed5f483dae4650862e38e90745f4869985a27d80ac06d24beab8eefca8c3886a2d02d80de158b8740dcc60afef3c64d16723ea350261980f4575b26f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b4ab572e2f165ef8852a26e9580534d59d9bb52a57ad7fccf3846f61a5b08337fb21244f00914d053c6fba642db506c8c02650e521b08815f5f67512bdb31019fb712abde4ffad825cbe36312402f4d5612b13e6080f6020b053ebcd7482886ea2ce91cbaa2e591c66080085ec8b5cf8b2e2004871f5f4df4a6562380571fdb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfecc03022f4b1eef384ea463f2e50cef40d45fc22b2d887fc730cabba0efb1c1861a61ff271c156394d186e51c48df1004852d7a0e49d737c561221152456e1a13a16c8c5ad0d4c44be98356ce81f88fa6f75377850a3e413b7c96a3389bc7ed951d5df38a7a0d6be5dece3275c87698704e7aa305c65973615586adadfd42d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb486e5bee56a224d4bf0976545ed6ac4cf157ed74eb92100c4ada76641636caf3f77c47f87af9750f0b58757cb7ed6cda75f5c03ac214bf9492d512950f651d503cd9b0a8d58a8cc457db907267905934897d458c14860bc60ab47e9d79f3873891e6b75e312d5607047042d70be495917debe37e5cf9a269d98f30395ee236;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h709d7f4bbc0989e336befb3ee35d917b73faa2be29ef581b554c5c4440cb6fc4a1fd9ef3d30365a55c281926163516c835d169eff8ec022120499746bc800b215a8beed8a3091896791f3662307692aa2b1dec97651569bb20bea9ea75c0868a8684506ba61d1dee41109e6406f70e13df9164fe2d23b3a75e0b75d13fa23efe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h64df718c1c074c016ff27015811538f365d5517e6122a49c50f86b2d39c53163f3c01ce6a22cb3d320a6f0653378c86d8e9cd8581d0c8a3dda1fda6c646373520ae456f1b74aceef0f87b2e13d7ddc3b086717c0d31f5f8d711fe9836ccc34385a15078c741220c6099c3a73a6e0d5b7cf3f66afa042aa27e215c027ebe6bd23;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb30c3efc73f84f28d39065addfc1971491c20b227674d220589c0397729a182e4341b74c745c3ba7f2ddb8f4de811d578b728957f7766822b40b93be421c21be67a4326b25fd2c01a9646f0fef9042972f575fa7d0f74627e224f92aba6dcb8903121c0bc2ff32f4d98f9cf61da86c16f3e0a717286b54c7ee11e2b350e51adf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h734632bfa8b956c94440afe9310fce415713a08a7a8d0393199f3d0bb787a63fe6e900135935b574d9b75428e78898f59676da0e1d7626ff8a65ad7e6cd3d1299039e99b563204f149a6856a51f8ed0bbd30455c44fdea2086c8a1653e315332de1ca0367da14d34f0a82af5989bc66a5f1ba1e919965434ad338fcf39bce2d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9185a0e00a82353de377cb26982d72fd72c9a76ddec4714dae545c7eb593eefd2572814aa10d91dd78146e9025f4375f92b97ff7fc5d626bdf3e210e9a29fe76f7521608b1528c8caf207febd574518800a4cb0269c9c3a659ad9e173b8d857ac53a1c60a174d1e54e4dd1b2941b778f25ac95bad2a6ed79cde2dc4b54ee9357;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h788c75de96d3874faf46c1e5171a3b026252f4b0f2eb295379511ac0921e8f9b4d44ebcc233c7d8ef0a1e0965094cdffde6415472e4c86cec6351a555def55c1c41c00f564bd34750d2b09dab35f8e18cb02d500217350ff19f5e8b22c3628d95a281d718de099c026b7195bb1d22a3dc771e542597506ce0cd4c3a313331ce2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e1a3cb05aeb0abf0263383db66d09c394140ab0305a0d1774c0029426c4031c93f0225914b7fda646d15bb565ac88482a615b3ff370ac05cc72363fb8e352af03a6f3edc70d1203883a59c8e2d975d258e6b77b2e991fb886a354b044d1f823d864e246d5462d6e780c5eeaf1766030abe80026c6671a5f85ec6243a854ccfc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5da16b20f1942822c81c1d44bcbe7f0836b88cd4f4352223c50fc94153fd093484d254c3f1a749924919d4fd4d0e70792344f9e4247f31853cd7459a76e5ebda405f26476f4d9993ebbe6bbe20d0097e803b1fdc041aee948a5709b966c8ea9eeb9373c5a5b0e7eb775215899cb891ad762fc8852b76aebd2b3d2ea6e799da90;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ab5175c0e9a03b7c83c7bbdb0b5c08d8c3900f3d26d2e5050f18cb5366d1d81d59d788b59aef2f36144ea167d226a9a185251b3d4cc3d8477a869479b6b7bed8683cb95819b1a7a76b3569da3e8bb3802321c99d69dceb6c1f9659cf5ad9a46b221fdbd09d02d7d3446d373b7a690db6d8c6250ef07d1ae1214440ea0cb3b7b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h362d16f5500c736d6f448e190ffb410b3956e4f55d7a57306e3cae87df94facfaf3b4752be7704025725b9fc76a6e0091d45b73aa5adeeb824cfb1d3e114f494071245664ca121870ee0f4c5cb66efdbcc06b5441d293efc4d42caf4265704887a06dc3374a161f214e958338a04a8d6399110d5aee98260b6db681cb322cd52;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h604240bf8cc01aaa65d07290926743bf7d06aa95bb95cf12950d98c39f8d56611c13e52e853f69e9c589a124a18d805dbbe45ba407957d596928e405410851a795e6c4ff87b606a77fae1e9e68279d631aca45a809c05ac476d967906c7e00fabd481e69760470b1e829db3bcf289239e2f3c60df76e5f436d7788f9c8663fc5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81ceec42e7612b7dde1f343f0745950e66fba9475a250a22b0f1aa7943f4430cb19c114e4020eeb6e6ff65978e51ed96b97e24f8a8c171499e9e4d306d5aa7cfe456f21d668d645e35103d7f6b72c26ca18221bec4e66773bbf2e94c5a879c07ee95f2315470daba392b1753f2d216476a8592e5156be4990524f0c9c3f6c1cb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he82bdc8bacd4fd1707af99b37e0e87200617044135c3601f212792493b2e8b1ca3e69c0619a942a33c03d0c78ba24bdae33d7afbc34e8c1f5cb8aecfc0a5886272ce87830aa4630bbe15109e0f88b4a216b6a552a0f2dc42938cdf22c1c1e7b06d1d27ee1c14557382e906caa18b9776dcb7d09509ab97c986a5f2e90280cd6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h202f3353fc50e97bbfa372eaed99702352da0eda34639cbda476512b5c6bf849f5a8e00d1807bbee5f4708399aee8cb046e935b0e9f761b8f40472a4aea1aa2111aa4d96767c45a88dd38e1bcf972a6670beeadee77bba680a7daf32f88d8aa15617ee40ab54eb3168a82e92e85950da07befe3f458a2c188db09cd09b3ae557;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5de35665a8f7e58bb11b91bc9902f50b05ace43378fa3f50fac42d4f88516b50079ccb21d3d7d2ffef98212cc1ba842be7a6a2cd1b3ed1c0bf967c7ce4898971d6ab641817139fdfbd0430e2fd13f37c3c035fb6ae391ba0a88d8a1e4dd681f1255c9ce4c883ce056f70875df74f979590ad9964c07df93ade18b605ce51a103;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h206244706ec485b165ea331d7f68fd762b2240b30ac79f22e532619cac4e28d5c32ea8dde08488c9dac297e0f6c4cef8a4a062dafcc9626e2b82f4e89d8387f429333082ca2e3844656523cdcc1a78ba2263f3203064c3c368d635db3e01a5deba842e828c5e9b0c3f61c47af0ba2e6fbd73f620261bedd1cb357ff7b85742e3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c7b29ca898c14b9b11285216a586d40acae820d428b3b3a565a12187353a2a6c59ab29ba7715f5d294fd334dc10bfa423bba58e6839ed70d0f778ba1bd10f2b80e8cab1184fe5ed0cc12ab555f7b65e4964efcc713aa2cb783366fc9299df38e309e23bb119d2b215813704e0f183bde0c8032ecd75e3b5026b1eb570f41e5c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6ab58b3f9d880b93a4b4bc664f7c808e6382c7af35cbdc3cd079d21f9d04cce2ee86d2156258cba1a1f55c1a308ff4729b7194fce0315a8ee2521ce04a6f7d1b563d51b9de30143dcc16a43bc237735fe8d925a7b85edc04fe734ec36f4059650d743cdc235f0ffa3498e37c048661089c9a3e65d92bdff270e8acc740b8deb5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h390eac4066a9d92b9e8b48004c0a2c6163748a86942f6dac10e7c4594c4b97b2e89ea75de82004ba5631675bf3959b7985614d7074867c2e3ca55ab7268c8d92ed7755b316d0a4d5a2a6913de6eea864d74a7a3c83f2549814dc88da4138e39dff09e48cde668fe654ee123e548c39ba6f67389666469eefa65e2870e2a00ea7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8fec14f266777b04ebb5ffd9fdefc1db667a59ab355435907dff251c1e989879e6e23fe995ada790a09c79d958ff2749bba341fd02205b5afc9fcf5206bdd6b978662fc9cea105e9bd9ccc5594b36754dc9e24ba246d554579173a8b18289ae5035d1d4f88b0b2d3f4d54c0e1a4757cc145c3202024072be3309dc5d3a453fdc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1cd25c73bd6e183dcaa03e5cd0565bb9e1caf57d78a5ae3639a7ad8a93816b29e1ba143aa932a92cf48a7069fa37dea84c366d07e402c7d6d01f2f352267ce0e6e7c51150c840f5db67fbc74b66a45ff3d5de613af349346bbae9a271b66eb066e5c94ba1047e53f64ac00dd679f05f2f2e5b7bce3b29186db8a77dfb10ebd5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha188b89163b9322d829d7e19ee69c775e7f1ff70e96b262322917e05b5a220674395663a6f84de732391c700a3a02e4f05a303e727bbb2e9b7231e5442296b3362ba713ce2d4256ed528eb88bd92503ba7613f8333fe14863b9a97ad6ff16b2be112115ccb660aa7232ca8d675632a86d17361518a45c6ccefd5fe2bcc45cdcb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a248a09c75d3f76c08a460fae671444797aadce2a23df9488e60aa4b0b3e50a1a986133646a05939f4815f139c41af78083c5f5193353f2213b3b729a6377e7d1474e1351908b5f2f0fad8214f09d31b2969d6b94b23e0d4fb7aadca70480db9a0e0edf7bdd8fe511752bce77b2917ade4f3546fe16bb5f51f308842e944a23;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2236dcfe0859e82149b037082ad99934dc6d1f9fa2f7c8f628f6bc1a7932d6fef369af5450be0b9f6c8bfd4394cebc85f782bc5f734fe9d09cd41360e8934211480b01469bd760083ebe6025c0485ebcdb001baf71426594c2d9a2a7a99dc70383e2130e99e49b4ac971215d96754f148193efc174872f710597368f0e85ff8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e43c15b49072f5082bde530ece271b0582c7390bb1a18a6bf903cd3cd1abce63a65bf7c4ad4af7eb7a6c820f141b875b3fbe17c697ec47bdcec2edbe78b0f282a08237eeb891168259d54c0b46edbefa195e704c2baae2781a258dc3a34cb493edf5f76bfa4e97b7fd0a66cabe3e877d22dabe1d11f2b71860f528da9eab66f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc567f94ec3b6ea7d2d87ca8abaa882f8a2fa6224c562c457ca3114f62f4df803f247d4e5d1db64c214519cfcd3363223665e4738a6a58eb75b210df4e86a163862a72fc3ffb1a10e4109e0e9d610cf5517e1e5032391ed58f11e7c003c1426ca2b248bdfefd22ede72ffaf3bcfeb21c7a27f85dd117c71219e616248b1ee7c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb0ec50dbeb1a02ebe347fdc71d8e1f089f19ce3540cce581c028819872e3ddbfecd3e3df20e0782f808585c02bedefacdc5158117acddf7a7622519f6949d49d6eac1d7de15cc7d82c10e2eb672b60fa9ef1e1b571e05c3b55c6cdac4df26c03302bd1d9a0356dbda1667c7db6fba43a098a74faee58e93e1789131b1337fe0e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f475c7d51aa84e82a0aa48a5f63df9218bee67b01d17fa5fe87070279bc84918c7088fba144bb27e6e7e4ba7da71353556597e8f2e9369dc5cc8c44d4436735540beccd28ea6f7e7ccd0369e7b9d752f776df4ef2609cb064152aa418049cff091d4b5d7463459c0c7cf4e96cb27d6f02d0e437afe37c5ca64d0c29cf9da06e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2599088a09ac6967ce81a0a890f3f6f413cc24fb3211e2252225a1f5afb87342d0b4fa509a508b52b1b22988d20617f7fda69f888b0c0d93b42db38344846620482149c9e52ee8fba19b015c7086f64fce80125ca8c89df9c6c3ae3b33d55c9e5f4f2d232b4de7896cd2bdb3e1ccbc40636e59e97d863ac58c9b6e777e455442;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf485f1b394894985eac9c11037e605122893c53ea1d1457d849a0ea73a08b99f9e3bdf51ab4f84dd795eebd68db622658d0fb8462fb7c6a193f6c56b4e63180398a5f432bedb84c0b614eb500083cb4af30584a824a00bbffa724ea552f006bdc771c60489e671f1b3d2f5622b88c90d866484f80150260b2d9073eef4ab20d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h65f5ae803fa5062e1ed9402232cb59c500373053ba55732978a216778717bcb4037b680f0d859c85778756c2a3eac2c6550e7346b3cf285722a345b566f622ced95faa2102e52fec75fe599e75a285486c867d54e9aba762dc589d92ed4c4636cdd9e45a822399d7e9176a985a691e53395e50343e5ffb5689cecf34017436d7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40bc81963a1b2ae54fb4129b5c4e1d4023d385f6d829f2de1896b277c979541be3b6df250a9886b84e19db981abc158c1b3562363e88867808fbdc2f6cabef5c154e588b016cd50e266657ea4b3a709c1cd0a08b4fc1121f90b08c819a5b29d29526699dc6c54c56967caec80fe7d9e1cca9408ba5690d5de847cfdfc69a378c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8801e5f3110b1e1017df76747f1775d5a61e76fbf22591d1ccd8a823ba91676db983c58a3ea7bf68d128597af99ac46424d94c9d31ab7e8588cb0dc987384de52b098ca21053f7e21a88f07c1ca06541e478abdee3f1f1fa6173f6c2487b462fda43dfb6224a853a01bc332f2f8c60816a0d8ea824108a295a4363647912e8ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had8475b67d7d25ec5f9a5e0214622cf6a90d798ca172dd12ab8ab4a591961b3e183b00cc1aa54ac33a6678a93317f035f47fae575b9279a5c5ba76938432fbe7eb7fe4c06f161565f4d77e4e95a00205bd08c1a919b31ab4efb3b663f257bdb31e9dd0cd2c0389a0f02342d074a5f0b7582ceee7067254740c6064a0d0bd4ea5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd750128f385291909abb9a851bdd094fc4e094fd711a3f9453c825134e51c2c30a821133948bf044f56f626217b5c4de1dcff0c7da0d3d99b098b65fe6a9e6f75807ee2be0a268e5bc35be9b9d09d8f380a1878f32fd58c652234eaec588f90aae070892b21f88cec0ce027842c529153d4aac992eb397a92e250dbfceaeefa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf35a47eb119add353a01bcb46238fc83b5e8d63967fc4bd9d12f80b42857c9a5f6e05500ff456b1e91d453117b7b833430c0a9d9dfccf28a3f4d337297a15ea7f0a630edf346d242a5d9d88bf162e2f8f12ea414e8392f76aa686ae5d6d948af53a2a07570661d7ed971a3a39c98ef6a9558760ff38d047b6715695c6be4565;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c3302aaf41a5a2f2cc8345f57ac17a3e1e4280ca620dee46498836b96e1a16129d1f63cc1b4edf8b4be00c2e5b226a7204b1da8c721e592ff81375c1a33e328b333b28b878439616aa1285f34661044ca402529ce06c9fa84ab7f365d43783dfdf1d888dff0b61fb29be206be9d1f6f5fa28cd82a1122e9ad275df15236940f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf18e326eeea929908744d12bc7af0231bd4fea235e7f11b46a9031c8cddddb1bdc27128f011f27dc4ed24bc65fa5622ea13e29ca3b89eee76ba47aef9b79cdea7ead4ed08e6442f9717056e214066eb2f3217823289fff0f129b768d5d7ae9b046c090f08a9b3c122cb84a0ca69c36d867961d0670244d1d46c4952b34a041c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5fddcd81d7882f3c4678a9b7263923c2215dcc13683f9bf0ece9f2d3738355db3b8800f986edd60eab94c445ebb0e42f0b65b07a7525fef7e0148a228cf5e6fd489dcf7281aa636fc42a090e96408e14cf429ca7d6c658fbf3854487bafabe0dd6432726a06bf2807106214df3572dbf4e787308f2e0e1c1d1a9a81b9edf3317;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62fc83112fc5f62ef0b3b73bd3838b12f4fc4fbd21597fbec4f8e04c2433b3940d6df2687ddaed6b17664dbeef00d49729fb6fdd24742c87accc4f00c063df9bf29fec82bcc23dc5b399ebbb547665abec00849cb36514caca524f24a124c83d2758b9aaa0a3b752bd18f66d7622da2bd6889b2cb3340da20f06e02d81ced416;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5c4c16045949892660dd104c06af3de68690320d3582c4726576bc35bc2f01841ef860f7ca6ea66293fdeabf45c3bac021d2a6241958a7f795a077db523869b69ada16c243bed3906cd170efc933d3b7ca50ecbac172c6f4dcbe735052f39bf53fac8117c18e903a867fc5a2fe5b23639cdfaed48e974ea7b4d3551bcd0f6f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1411cecd8b9cef160a2e554f311ad4416ef02324c70c1439947b8595c2271492eac288c5e4d22fae221423f369814aaf4839ea6d8d8dfba8816cbb05d405d87cd0d8c1681d5aa02b60d524879e862c4a0d670c5a0149ddbc4d0c4f34e7d0ad31e1ae114ec78aad94603d06941b4cceae325c9f8d1957f85857ac58b70fe05558;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfecd393337a7d97e5cf5464626bba656f9b9eb35f493f2c36fe2c58e2239b78f159403386ab1d37d77630e73c3d71383b8bec19fac9f642dea93c0aa66769507492350b5f96564877f480cc3b960edc22cbdc07cbed85d18a7e445941853f49d10271d4d731134605050cf12d25a8fa7dfb7b785306c2605d99819c196ebdc9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1d99fe0d4d28b921aecb05ce94e7abcabef8fbe6ae123d3b3773995c0b3e4dd376812f93a15bc6d681adfe098e482c88dc257b7d6b31a7b837c350ff9c96e78d5ef98a5347c51f0aa44d2ecefd226c7e0aa617782bbf364b5da02f7577b6e2e9a8b9e6819b2ee45feee398c848fca53baa2e80fa3ca1a4a0bacce3c61b28102;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1fdb2f085a4d4d289f4aa110700feb57f5e53e6f37326780c559ff8d5534558af613f4e9dc7a22eedf3d9af22890a6e97f4813b72b2e659114d88651d24cfa942b165e9163d1e66064f84034a3b24feabc01fd9b95c636400d2b382f8fe78252a6146f43a7607b94c4c9238ac3076ee68d7712ad7d687c15f5624997054fbbb9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h752e90a92f6430493b58c10f690e337a5f3240bddbf3c23faf4529977047b48791a98de587196460c2940f25de2f0ea62491a98d91dfb6056d3829060231d5d4afdd04eacacf6ee18686f22dadf2dc260bbc25a643a9b13ad0af0755e07295193e4e2bedfcc6e839f9d63770fca850e37890f51da56f305aef840677f7d87f07;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4d1b2faed04b583a3e6041f96bb7120204631794e51c8d244e76190933d981b4eefa480a9ee4e3c49973a64167593e69068c60b996917a04bc81c4d31e41117b6e8455f5416f52e15f5a8a81b533de8d55f84cbc7eeb072bac83d675d41a3b5509c204f840bb9bf95c20876b9497f54afcbd10df785679c56c917f4b4c5dd4a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcaedd9f4a66dd777f07ff609c060e5baf0c9a96a22c5fe4dba8c1da613694689ebf6a902a2cef658431172649c7461c05f7a3b0f2bc10e1d7d2b3c19495296f5b5b8acdf6f581d6e592bd2048da9efd28db51ddfc96299240c512c9b27590a765a237f329ab0c37cb0806afc94c21dc993e2f49138b856fb2a6f63e9840a2d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32d9eaf50954ddac7783aee98ec0c3b516b778f41ed704ca3cc161f4868e59f5ba3a5f9495214cb4a12b96b839486e998c3ba94cc3ed168e995446855e32844916f4a1ccfd9fe4032ad49d67fd4b78eab5bc9998460cd85a138f1f24315e1a86e37de0a4c910f5b143a1536c43542c00d792b54184aaeaa69041a7da035c6a62;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7769417ca821377b8a19b7cc4fd8cef126343c42fe63c24097ed741282a5670d2e54c5fe64128986a7977c4a53d134896a2f97a6abd2b20a88e1d2e2ee7067a4a4a55bbe7bade70ba52ad296f55ef5fe4b9d01651bf1343dd33a3f77f504e96ccf61935d04df815e0a607fc12f697acbe99a59044de067416326c1ef769f6b20;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he01234493045d86d560162909586ef8251bae0344be94f22e03f2b965278e303f38c13df1ba49cbf58196edd3d1602d6a9df59167168f75d0b3cb9e807352a917eb7debebf6f12080f5bf7dfe6daca367fcfee0b5e50557afd14c7cf0ecf82e30a689ef17ec79b8f9d84a40202586f242400110a5a5d94992f6f1049c6162da;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha17f115753bbc3c2830294cdb45fe129e1cb07b8909d6136847df1530c19df1bd333a713da2444f88e1f290624daee43b6d91881231fd3ba79a0cf2f3e250bcc8415e93cf440a839ff89d9509c3de7f8f65d0d4db64d30d8a55f951789a536f3830d49ce2ddcecd621b33354e5843ee6cac698bf3dca548fa0563b87761d6f9d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd1ff6ee5d4bb9a0872e8c78146342c68febfc6a0d4c6cdbf8704180fcab237492f3bcfdf4bbe1d04f1158b88a6c930c400d1f91f1a79bf2f2dacdafdc964463e76ce49051a1d2aa861c1b526b596f8ea5959c0f7648bec1a24aa738bece6d094b0bce3a25886650129e410dc9528628d7f2c5363eb3b650e8ae1bb4e3e4cb7a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3ae94eb4178e072a93c14050e6d285f5257816b0d8751a8486e426a491bde37e5c83953ff2f2346a2576e0044a1ada04237428600e6ba143af7fce5a65bc6de4e8dcb9e037b5b62aff854a0d0b5a25b66b999f474e98e3cff1a56d6e20a0bcc640fb5d51983ab4478525a75563eb6aa58b036ddd8213229229ffe92e0deb95a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha31fd4289cbdafd77cb0811351d8919d1a43d13aa335aa2278d6e7586ad8a97eaad156a7427d99d6a909d7ef25c7779ee5ada1f846615853e8fa8de2423a6c0c5e7c094b74293ac7cdf68469f3d5604ee563cdddbd8f2a628f4aeae0ad44aff3d7586a86a8257447e88127f1ade655f3bd281a0f8122a294a76d9981d827c51a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc4f709478fbdbfb2a3dda816e3025055614df90e7f544225fb36999dc0b8ba975c0aeae06babeafba8d0bc436cf649140fde2feec3c2b33a225b89e4d236ba4f31b91a8fcd84e723c6daa8f09db8ed416ebb5bba9634a931eceb648d233643f3e12b43534cff63f2f161ae32ab6aa09aec8cf36fbca4aadef89bb7a72f1621a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h957ea3172a477f495945125dac1735e93fcf8400f92c5b87f33d696c0331d27605c726421484fd97a99862624e8b60aeae637886fb733c1c8449f9fb26062b60f8e024c5f12d493ec98ead20a50119eae2a8da65c136c533787c77e805f622804b02529fdfe69231ce1c0151bc92bf03dda32d54465f1d824a9ca132b30205f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h683934421c57914949d18bd2d5d45bfb7b2604cc8c78b9a0ff65c8ad0618824cf291e8fd65a930d3010643b7bd4ec7c3685843efabb75926db3c69e51807401644509f411a23c34db57ffd7ac6c5881c799b473cb261db23df11fe3bb15e2f924c160b2830c098a190136fa19a6385a5b8ea7a3cd62f52be1c2db13722742529;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h68de8eb7d8927624aa916334dc117b89066da32903588d55b8fe3ae3b5a2bfb29316d23ad89cd90c3f912342e5a3bf5f15ec5fd3fe886947edbbdc48821b9733bb81669cf57db87a59ac39e8564e9a42289ff5fb70b56f0899a7ca819fb0c9a3fed6c5e4813620edcf84be835604cac0c9bc9b4cdd0ee3ae933af60fcce14ff9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7464836b9e3542cd946ce53d4ecc999b557832067fb637f10dc002d6dc84493fb30a241d21de9cd778fc1733634a1de0c0ef5ac5c3323cd9e3339361932d5ddb1011b0523c8e58ff9ce4542771c43598553830bebfd99c2bdec90811ce837958f4aeb5f88c07b582aee5f5c79780ce346764a8676fabb8433288ebe505eb655;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7c1dbc70f414d31bbbc67391ebb9fe8a5a4b485d178883388bac7ec56233ffb1f0c30c2df9dfee1681c63ca2ce5c7077ab32968e1c8382a19b49d4f178833c5001a2db76a48c2b04ba845a49515f20fa1b96126939c9c691912d57d546f7bf286d3a4059dd2b2668f0467c5892ff1da449cce8fe546b27af0abb52594954a61;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6495cb167714966dfcfdf1bd5de06490bd635785baca3de131bc3ab6f8bce31bd9e976c9ac911f1061b04d0bc24e9aa501cb942082158f8d59d0a08f5986c04e814f3bcd4066577cdac0f8fe0de1e7bf6eee6d391ab2c44ee2a57224a0504f56d4dcecb62e4f11548fc3c492e791a25d60727075d87201cadf2025a60e15e0a8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb548a8626edb63369bbdb22d6cc97b345b7d5c63c59d4d291b99213eae2b3449b019b77e7d0752518ca12cd6eeb2aa299ef61cfd7784796d5e812410edf4b844ccac163a33632463b26d4f9142601207b6529296d70e6ca98714f92ce579a7469ba973a9b23929db4c1543f25fd2c43434f6b792f939d6bb69c57e8c58e7285;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf3c300b7f92c89f6463571254eb7e14c5e3797c82f6c22b5e3ef01045c1b662acedb3a5408d8e21886e1aa8e18961f6434a7a029c15181fd0a348c711638c95b2dd814416a8c3b1959d0e6baa8ffb3da8a5aa097e65b86892bb01bd930d56a9d1cd6742ec56631c9faa0522b189b9a9845b0e81d457db6ccf44ba6655a7882b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haec2355b3e49903407849ede7f937b0fd2cc38896a075e659e8010f261303281bbbbde1a60e8e036ee54b00823c519f65364a17d24870794d287c5c6e6d85da7987633fb1a24a5458cf2214a04a0ba9a114af83b7dcff4a61270a2ce9b3343b733f12c9620a58e7db68c6845556b2828624102619fc5d0c97dded58c70e39cf2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7826d163ddd69bab2b61945a53e7735a30c700d2183e3aa6579843eaa26c227c2b54449e0e259c9d702e3975c8add3d00008ac472a3130883d6cf27ecc710b64815fec1271d8e7ea68d516ebb16ea450cc417603b3a34613c10129e99533ddd84afc83149ccdf32c5a2320c9125d7fc3b18d6b2824b8a04bc7dcf4d690e09e83;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2dc86c07ff21fab8ca9fc8a999c9f25557fe76130a71d3903d33d1062060824375e8326cb38cefc2e044edc052ed8490b5a9fc8a3a6048ccd71627880618ab40b52c71df02ffa138b30b7baf2e268b72377b2464e8ba7790b9fca350bc0c1ef06505d9a5ad9fa895bba418ffc2c0989c1462c8b0db402d4192555153f9a6ff20;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d83cb1e8902bc10a90ac8c060b486aa1acbf476aa33c26ce5c8e5af1de9581fdc9dcfcdefbe2c8f5f4aeaf3cfcc5357071354fad9eb05f23f67dbf2aa7cefdf5c31163f156f619bf0fbcf302f20d78d523e8efd02a6ffe019ab9a74a0aa36abf769c51a07629ddd5b0f16337c609d343a71e475426f560a56a56118975356be;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6206ccc0991411645ad5132e54690a2b8bc2e8984306d1b3fbf5e65a9ccca6713da542cc274737becda3b0737a37ce1e40dba99be5adbe99270c791a4692e22b2cf9e55da51a1e0aa99ad2d65c92c39d54ace6f8786e4ce8e50e254c3cf88440737eea3d4f16ebb5cd3d2ceb18034109322f88eafeb78d7413606d251a4ba6c1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc254a4ed2f4bfa52b279101fe16d555dc0b487ef20a658f2d47368b8b0c29ece84c18188cda0a4eecf7dcd4a3189edaa9cf2887cc09b08296cd6e7aed1569d06879c66d0ce6cab344e91c192c9a101253d9b072eea335647724e7b2ec6acab975bc0796224ee37ceb723f4b2a2f4a2c6c97f00333e434fa4422b6b43249888c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6cccd32187720c297606c363bcdad252306f8e27b7b82bf04e501f6a1e8550fda20aef9308a82c1429a444b35e8b9a0f4fc0ee9fc05f3325bbce35c0d1d0f8017d6d335a7a2b121f6c85ebd66f015d54f7fd40f522a4ab560f3e1745f59284c01dfc0edebf1b768a960d1d832842cc45204e31d4709e250c0a7935dd9309efe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15bd1ca123680ecb521055475e02045369e72c6c851c9252c9c0b5463563904d4c809a7ad8b94c8f4a890689f41ded46aaadd6e3ebbb67cd559f0ceb074c742d0be3d71207c48b7e40f99e41be3fa8a6845328ed798fd7b923deb98ea4830ba0539ee6d23dac9f88dd459bc360cc350dea14ce5254aa8f5b3a8f81975a67941f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89348f6f2d03c2a4a21ba6bb8c151acd19c595393a6a4219fb31200b74c704d5eba5ed5e1c331276ddb4dddcb7898c0040c0fc6d07b151ee25f337238de940f4237ed7889c276e5310d4af13d8f2e236f529645482252925488bff4a05f6d18a1c0657c0062d70f9840797a52b5575b0921d32e9828327d2ff7e389cbb8cc095;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he8850c6eee615469283eead067157ed56893da8b801f4f62b9479ea3669c55ef41570f5b0f844e28d424abfd9a7870bb499e8b60e3ecc06010fa1a709fe9a469a0d50873ec933af9b7765aca5b5ac58c9c9ef2c648130876876a963fe7cba963087e188d50e23ef396e4bc49b1c7d6de6643a1eb1e0d332573648ba8a71c97b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbfbcc1159a6dca4f8d5adfe63f01724a46d7dd1735e14a2d789adb1a8226599de8cd318bc5faa6d88ed459ccadc307c84f77f782b067aa6dd61135d668423f26e05b2d1189c685ffeebcc1b4e59557c58be3003c3531cab8cde650857743cf26aca6fc2e9f9a683313ddf5782f9c736cd372dcb6fd78a7c62bd3ccdc1b5ff74a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5718b53c1716e96fa0084c05b04356b0fb7f9fa692fed29b3b9c4205f54fbba3f13aed9fee9f8c0ae787dbdd4deb8638c7451090ba190716baa50550898cf41dda2918e48780a7f258d15b9b5d5e1f313729d1fbb885c0da32d50a98bfcffcbd35ac2f7582dc94cb9741d37dbbc31fa860455b091453bdd415e4732fea8bebde;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54c03474cb7dcc086dbcd1d413f50138f71e4631f079b57506d87571de6dbe8be3935d1f53c79872c38837bf055570a276418abafb9915a145d041716e40fc961a0cf6a6fdb4f914ca84754d71a4c1c87a03a026f5437370a5c20c9398494552babb3c66fc42038380e0f802d06d42d1fd466f2fc3e8a2f38070b73e5598d0be;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h440c085625d9ceef181f4a84e3ca9fa361a6e960a5a544f894a39122bf52ee3893d6f7a825ed02c49afb5bfa7898de105607c8f858283e95a2e10bd45889c8139d252daa23f351d3d16e378f98ca42846acefc99d1b02ff7804cef80990425420c54f1afa05a4e5d7db190203a1e2846350e54e3585f322dcdcd0446cd3426ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e72d783e56f61840e4b00c23b56c299c9773f8578c734aa2fcc6c92947a5acd935017f37af1a7e52837b9b89f3c63927ccf3ab29b4fd86123bc48fd99d18c998b247ee194458420fd5ceb313112bfac38f8f73ac168fdc291d99c48d18173f773670bc973c7a4720ed386a4320505733c1d4afa4dde88a24ad0ba6de9057d82;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57459ef2384723e0bf8053e517ff1c8006b05b19dee552d42efb3b68085df18ec5d0414875390a1b5acb12bc5d20ce5a0b593960109c666974c19aff10bcf15d2a52404c762f569d648738679139d67c44c957909735b8b4a494cd297bb8ecc956a785cc226af3f01212ee136e24cfaabc20b8d11b7a019dc4160a2ba5136f6c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95c079a0923d9e4f06ebafd96884c7445f7c561d67f4960fb3e710397900a3d2a258f6f31532a97432d35f8356b87af4543df58b988ad0335981041fa9278da34998e1cfe198d013b124b3658f725f5bd894240398916d21c8252b2c0f438cbd5c52de483fdbe0b97bfdb5053d3bb900a281b3e4fe8deda426232b2baf9e9436;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5732eeddf5dd9eceea188bdf8320ee9efda18362eff5b2fc791df932a2c9d2220bc09ab10bc4547f342fef1723e5d20a248c80e78827b7efa692cc0ff82a251240d1c91e8885260561506f3facbbcaa14de417819a37c89b8a5b5c3380e09c81ecf7f58b0c0ee985f79e2b193b94e1b9c88cea4774773feeaba4f480c5a19d42;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha641c59a88013ccb21bba2ccd507eb045986c37a6d8851ef477a5e6e069c9ae3f40b7032c059eae8e62178169cef68f20b297a6106bfe1d782782d5440c0cc0e424fac996ace8a6d99be20df77a6d4d315784b095b82e7617f9a11f76221d66f2dabb9cd5a11dfa9832f38ee84d29d400b858806759421c4336a9723961bc3e4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he952f9354e60d5f62d684b2db2ad53d277f94c9910f630a39f2e5e363508d431397a54a8bd97aec21e41af6f806818baf59e3a20da11909e3a768e4d8e2632cdda042c40ee4472ca79dc3ca662f0b16244069064f7a34e0428737b7acb147e77dfe71f547893016d574d6051b0b0d3f5dc28f7d4bb934b7f87e7baf9b34cc7be;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h661c86d88104b593fe5fb763bc7fc66e82bf584e7be8ea9aaaac3cdd8b4bfa7cc2eea5db935907672ef0bae6d98c2daf6436ba002d701723d46fd72293a75b52fff6110a5c20131322910c2c65062235eef703ac76a70742ac4aa21d11f93e9d31aab4ee66b1473df504ac28f682c7ae97d1fb7e29d6d9d1c52949f2788429b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h933a32b8f92b1d80b4e921ebdbed1f3fbc090dae8c083925090f8cfb2eec01f96c787674bc02d2828b491748d6c513727fde638e4126ddb1a44bd77af2305dc586537594d0af5a02ae6baec68b5800bb5116a1069ebc34cde783542a3869e29da9fd9517a86189b10f4b6e3e2d77b4f84ad732aa7caa43b558f5d82a9a1942a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1bd67707228f44c956d18d6a3761dcca13c5ec68cc4213c237d5fe7fabe28cdaebb4b84cb7cf0fcda90f5f6196b201377c8feb260ae664301199e1a92eb8b81eeeacf08420205bac5bbedac551534e095e0050ec202e325deab6123a796f2d232d9a4225a2111b414308b86ad32e7783bd54fc4742b9ce7c0907dea51ed7a662;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88cf1d630b1f87e0638fd1fa8d7ca9b6f5cd8a11f6144ccc750ebc6703c6e2965a9c109f399694f2c973fdfcd78741ceaad34c7ee69171a7968dcb67803c80a18d34b58a976a9b5d641ac7e698c63655c95411e192d67c1b5b2ff6652b1694f7ab77a72436adbde0f11e9b94cbd9c3b48351397a2449dd97ff6b0a8cf7cc3265;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef79f540341be8384e433483ad5d0c26ba853da7d5e11038bd9b36a44695efb8e0b8f22e1ea5d9e3148f1440cecf28e5563457e5d75d274f956fb4e3e07622c4a93a489d451098b3cf559c11e98c7cf00fa084a22800977ba9594406f413619b9ba2bbaa0545de43e9452f90bec3f6f84755016266a4c7328c8c03d95fe39c0b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ab386697076e5fb399592e08f84c3f68f8c29c914edf1352e7a2eb88f05f4dd988b5a405405f51ce4ac98223343d11b9ef0d413d2aa5ce3c9753948ddeca723acad08d82630db6e6d50f2cf892b166d35f5b5068e1bb441c7f0067dac0eee646c6be3032dacaccc1f650ae97e8311689f24e26f8315eaec1947d78ad05f9aea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9730f8f82673fae4859ae82cf1c1c5874153f713bd81700a7e9c8811b4c0e0773c4f82a1f29303327b24a5544fe6a39295845056794f1641eec3dc243cf5e9b1f272ba83f36f00037dd1ba232e8552230eeee9692d7f3a067513d8ef31e6c2945cfba4fe1603ad97e231c2858cdb9c4f2dd797ca15767ef98d4d17f82a67670f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc43742a45b581766f563779a7718468ba63f7cf602fd6a1dcf10155938c1ad52cdf79fa6d33ef5b68d9efa7eb320ac708e8ec6b44a263ff30edfdfa37589d7124567167ad506cadfd41a08e6ae405ccc98f57f773443b826d4d4dd0d312292afc158ad527ffde5f678291f8bbe4a9c1e96bb49c6bf0ea7b6b7c0b07f60b4880;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e5040aa30008dabbddbbc18922f6c00f02b041110e6abeb8344fa135d7dee4c1c3dcf0ddf81e3efd31fb394d767022f57b4e03c5851cde8be652efcbb0ac230634d3b67c6b6cf0900b632b9c26949dc51f7a82bfaa2cab02aa95f7f5d36ac8af6c47d596b51bf2f570258d8b4c75a54d7b6783c1a66545d6e41ab032f0d91b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha74ba47bf814872ee87d8e36b5ae12433ae04e1f6fed4fa5a58e5a74f8fe083e0b2ca7f14b1b44f2fb780ca6b03f7d1a6bcf2016e1c50205f6ad941e3dd142819d4c17e55325819593a26846b973d070cf6144d38e72591ab30cb4104f4e978b4eafecd00b95c6d919cc9e635523838e8dca76b227a7469d1986a6f27d68bd27;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bd8b68fad2280f497bf37e32344c03d0d39c78a70a540af5963c2e9dd990d6d10e6320d3d076fe46e2b38cb972af8f4878a69e29f91916174436f32fe7f6eedba0dfc9e5f2bc855b86cbde7946f9a35ffcd718595949c99fa8c4b95c73d9c6bfdcb391b49983680ff6cce0a5402d134fca311fe44d046c7b0ff0c77ca0a731e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9b4749b016144b123f2ae5b7ff598cf7eb84ea49c49f575f5b9615b1fe3e3920a5dbac2ef9116a606caa08437e5e041546edf94fb9669aa1b56cfd7d0aedfdb22a15b585a8dfe89027c45422f0a13b3038fb7e751764a581311f2503f2118f030a0d5194e999ab265c7a3aeb60fc74bb777c9f91b096eb1310a297a85e52c66;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he88a7d1c495109da35f01b86392d547b94358f0b10dddda215f293f44ab1e2e432d4d1c2f5a48b1ea93c5dc2357fedd924743301a5aa151e74fa5c509606e4a2f73c204e8c951ed6efd7899a78bba7a124275408531d41e3cb086714af15213ebcc560b51fa93488a9aa5145a217a3edb977e2aa91e5dca341de405644d52ee4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdddc35e5a6f62e98c417d1392e7bad435b6896d976611538ab439b1f9c73e80e2ef11edd3d90f9243f7cd4c44074100a26d30a53271a8e797db22a973952de839c8a13d792fd6a4af14332fd62fe96d9afc942ce21ecf3df53476224a9142f6a03b44ef480c610112f5855b76c07034506e133f8425c88bb58e8fe06d16f3d5d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7f044dd740fb30f1ea63ff621064d9559ad19d8dfdcc35ecee46cdb9a97c382fbf982014e4117d77509b4da6028f9b1049e6c760544be62497845171e602c319fbfcda3a39913dc4b8ca37954c7a1b89ccac0c101215daf399ab138ff217b9ca05e815a52fbd8eeba5d6d377c11020cf2b3701762b1883b7ecdfa80681cfb356;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42edb98e60752fd7a59826e101d90847b2fa960f67da39b0fb576ee7e3c430503a3fef49c8f8ddf43d3a4a5bec7f7512848f89ad4158bfeeb6e95f41d1098367ecae3173913610871a01cf91bd2bd0fe08c9d24858a794aa2a0c167c39708589b7d41310bb22969fc87aebc3a85734b1c004ca283810c031a125c870e472c9e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7113afdebd02dd0ad7d46888f11dff941e80b16298d0b9a444ed911f921edcc0749bb4fdf5fa452b4e7a2c7354a53a83828078a14cc46dd540f3cd3007bf8a39c37cafea928488d864d48c23c8f8f6e1812b8d1e2af64a76286bdb0184dab66e0a29b3d4358ae5af29a7b93a80527a335a179758c83f5a3436fde6d1ee32692a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h694fdcc2f63977cd21d380a7c34eab8de3b33e63336323cdbe5aa5977aa6e0dbac448a177c9ce9a91013c1742e65612bac8fda66d42c519f6d954842e358c3e3491fd6c3dcc2863230c36615c5793a3f249c5680102b79bb00cefe32b5bb7838d796f857fd39bca9463a23d8098d05ae9dafaa3b69b05bdadc51f19fe100a32c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9b86a4ba63fd3da2e6f5280238e08d784b034380306b8fb1de2100dcfc97ad76163505856060ac808744fb3621e0ddbf30899ea9727f9656074e63eddd4ef4997d11f27ce801953d799a4c184c7e8ca08eb1366b7adaf6c88655f1fd3449d3e81795a479b9aef3f86f5f460e97541b41b1083b5221293ad4e4d421b59d4b295;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b2740e8c97edd267ea9c703510b3f45a2d4bb81f694cd501a3dd93eb25c7159e2ca5b57415434047f2d67b91ecbbb4c1e987bacaea16fdcf6628195a1fc0de9815810112b9cfdb5bbb66ffe684f69efdac61f4d185eb10ff43c14a57ca971273bb704622dd94f232eecb097a36e63ae43ec0921002a9f1d9a6a160066e3be57;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95d0017cc53ffaf1e83f86dd66aafb74215d18ba206614a62b10af386b457f450261efaa6b44522682706cd319bdd17fcb3704bf950bc7a2a55528eb03878999f765b0306af746ea8670e96144e1886e9d4551c0eebf79c012637fca12980241f17781f2754efc9fe300d74caf92b9670e607b2fa27a6db15fd26f6bdee47f7a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d01d3b1e977addf29e7a2de81ab7289daf60f0bb10984825f7f217339197ab88a205ada114be025e9755e2cfcfb20815bfd8e01a2bcbfedc3b7b1ec5657cff19af0492543434c03bc348bc3d910e769941195e662eecf7eb9dd5f748fb38b971b5bea1aa8f2cf823a7b733ea8122a8c9bdd0fa562350382260531b69ee8bd6a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf480be6b0fb65ba578abbe3ac998785ba0cb25f2cb57ea7e6687a93fc59e59adde2f8c516658b332d3ab42cbcd4942138a107c644a59e6ceb78d0f3b1c4a8453a7539d3ed915c1d8b194206f9cb1f336912afc2710c35290c7a1c8cc669852ee831b9f44ded68b4f4922fcdd3393596142c34f8f0354b6904faf19b4b020dfb4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95f19598496d7648cb62f949c2689f24cf52c4a7897fd01ff5fc211ad7fc44077273b14593346ad77c9d80fa31860844c790482c103805c93290232a6a58e9b1b9cea5f3fb9fa7fc405717c443978220c94af45ba55855f770e8641ec0a014f0f0ffe6c81340f85b77049f6d758b6de720336a6135e99fd7a57d4b47569facbc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8ffbdc9110c62e855d2b9a2bb5b1e516f0053b4eb39c9ae23613c0cd2945e44975f33111e5f94ebabaabc4749dbca276f0037a17e76ee782d6273be9c40065665f7de4600ca38d0ed3b5e28abf382f402d99458992205597653e197f13d330e2cf4c71757627649927828d789159b70960a2359bb6c31ad913d3222552ee8d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd8784eb3080965c493f11477e624f212f8387f9f0f8eb3beb45f431dd251f8cfba69387bd2e2910475f3c2d01ae8a130b3f0699096e7d9d2fe37bd89803a7d0acbc1444617dc65d9dcf9437e4ce1fac921779acb810ccf7824df6353141bab504092953b0bd918272a8ae0bfa97be09fff6f4a27d3fe6d7c1a81453328abf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcebd34e221f4c80c628e25892d4268cad7a6fa6a56e9afc4e78886d6e7ff8d52619864214d9da4a7a4889e66490a767052694b0b9dcd9ca00110b4a3e440803fed7276f60fa2d2297769ce4c28ca51a3b80e4923537d869039becfd7dbfe44a15b1d91e96d4776b4df29f5c270317be377a2de7b49cb9da671f6f6c8dc89e33;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89cb3741d7fa9a27ee5c39e96c9b2f940bac524d49cc759e4d105d2e0ffcabe413efb23220b6d5164ebee4597aa9b55c5e13eeae7720e8e7d5cd3c3c5c4827bf941223387db6486cfc76d03469b605a9c77d417c425a5920d81a010edbe8e3413e5484b1508c3bbcca897e859898ea92ff624918343b2fd9a93035c4be5d9193;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h29305b2f7199cb5b06bae3e6796b906be299935217929955a2abd279cc944b92f3c1a62c862fbae2ed7a47478eaaf5ed097ee4ba8bc4633b9067c93ef84896d351a31090494ff1a723637bd54eac097521dec746e8d5000c10a09a7a02255f22b93ea021e3571d4496543ee023556a8d22dcc8915cd97fd35242b2be1b454feb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1759325e0d057c8cfeec39f21597c47197fc44ce790157befac401629666a5e6ca3e8dea0b0ba6207b88a12ba94a3a553662814d4e2b2eeb3e69e6f73b5229ff2ccf20b1edea990e1953a95a97d854a6a39e727c4d0143ea57ed1922881ca09942a509d9525db73089a03867a212ecc9bc09fbf2e983f01a85c4d16fa467036a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb34b33be71dba69ae758100577e56de1d589014e2d643e513adbbe84b53a5632c86fbde94e346329774886bcfcf720cc3c2291867811f963ef7930b45f295c5cf4e68e45bfb3f19ed7a94b27f48f7a638c1ffe093a3f1dee719f6a178b593ae28a6af3f4d38bb9d26f168b855d655083a2ecac6e370dbb64edd52e22d5edaa0a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11965c2756ebe92fc6033f04f1e5119a0ef881cefb2d91ae807b6890d31a0c89c0d223ac8220c6a5abe7e615e8564467ed30c5c315d7c48592ad00c3324a11418a7446d9cfd7bb1e934d888ee1e5e99a11ea5ba73209a4f3efb3b44e62f23f6eeca7e0b2129ea9c66066540c99aadf35bc89fa831c9548aba3a25f65f0a33756;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10a771dd1cd8472d086449ca0804875564129bd8298fc5a9580edca1ad0f21046383b8f1597c76dd4ac9990c97d7fba8f1b2e0f7ca379bab4eac6bd2ab71c489b1251d914411c49806649cb5a40c361b0c0b2fbfb38678b0c065acfb01f9afba728e48c1e755ba62f1eafd990192784091dd901aaa0a207ca4fed69503cbac44;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6603049ba07fb171a170e38386339849471c2ed8c98ade04909fc5d4ae9376e09c900d74ae8ddbf1f0a19d235e6a188a6070210c2c67c9034cd64ba849cd62630035883fe27d3c2fb9a5246d237f240078e4c0e18edc77025d3b8c16e5c578adfa365f73911d94b4e8bc9e92cf25bf2fe55bcfc8c48ca0fc1a45d8c1fabc3e83;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cb9afe54ba6810683ff5f5723cceb0987dec20b8dedb68e6511efab03f48fa9ee70e2456d9d8938c330e0e24e227590d1dd2442437818a76cad0675c77a88a83b21f2ef679b0a65cdf2faea38087ae6b7a2711aff6479733d5864995a52ce373a04672774178818be8b3c6cceb2a474195f1703e6ce03b23edb6b839c936a5f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfcdadaedbaf79b7968908139b236b2a6163b3f5802837f9852341988927869457b19f42ab38db9469f59b5c72226462bdb6aba6738ae9cd1c616df237f8e909b145bd5db4544bc24eaf236d6d9b6a0bc4c21d7aaca7f0efad4de87dcef34ec0017a9fabf696d8672cb98393b7a43d3ee137d8ac33c866ce6810c816ba5ec0148;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb06e3aee4edbdf45e0e109f3cb7e1b1c10ae6e4dbcb79c2f5754740308ba347ce9591318189629820e4e37441def91cc5c9df81819f4d7653e7840eedffca46537c7afdc05be029be13782c3951f6e52d37e0fa919e091a0c6d82053603df789f41f23c81933c2da73e33a30877f4353f2f408a1cb6321335912ed1e9212cb76;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he37ee25cf1f229c86bfb65964c6d76305a254d86d0889c22a699656a5ab250dc6724a6ed59025aca3c15b2c3903ad6a5a9dcd55c465fbc70306906d94a565d4ec16b734583f7ce74ad2d6eaa250bcb61792bc265f954b4a53db850ff6f6fd6de5b0cb6f562130bb21b80ff03709e75024bc77ea6caefeafc7c0020093c851ed6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4abac4c109f2f64a625124a8d4b94865bbcf9d7fe85e0a9f82d0af28b315381d31df28750040c90e17b55157b9cd81fdf74fff86bd23caf2f399b10b8cd3141006ee5bb948bb89bd2294ef6f1b459a954ea17d056755a06640aa5a66f7172759791a6d28f0637c875bb4c52be830ef30a408a16454315019ce20b57f1204535;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h240bd884de26e6368100a6e7ea71c39f42f2a10d8dc8ebd7f80d34c83ee25f7dcdcf5927633cdca3a148f16c97cc094d94a20ca1f7c0b35a06cb1343d99baa26a2ca1774431b27f23541f23a0f924223a5c7da85c1956881ef947c5b08a6c85f66486c63c3d171c853e7732951f35bc4a1aa0280606f1d7705ba3d69535c5d46;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7ed45327b4f280b35db7c0ca180fe30f470c33ea3d6806926864b4d2c477a178298baab8252a87843cbbc01b2d028a92bd50599cae9a9611af03b70d434de6b77fa529b074bb9bbfe8427e7dd1f914c1cd7860cf7dffbd85aac68ee2ce8537cd8042e62587bb9a76f7fd22ba8318e7e443ae86f7264060dce4703c3737c2ba5c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5810eac67db80f3048d8149ee7d49f2cbf80195c118def85949cf78d2f59fa77deacc040d2d05b90ad01ef6b7ec466ca6f9fb5679acddfec8f285c5a6c7f8a32f805f05b5381c51393f8eb8fc9d2ad5bbdf9b83ebde08cbcf2b400c923683d68f618559676e7b53f9bbceaefcea95563616d1f7cbee0f3d57a33a084ea473e3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffa5f3e28357f3d103fcb53dcbe79ee0da70ef946a4277b69ad56e8834c2f9cc3205ffd773e25373b3e2eb6b640bb53d75987fe4212c8d1515a5e4452d34564579b305e37ae7c09f116f22f3e97d9675438ed64376cfee36da0b803c8b6b363bf82937340151ad51c7af736badbde8037a015a84ab671f1488e3b4deccf19b06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf86c265840aed7046a035a07a89bd9eef8035aa3b289b149f0c0d4d6dd77b41feb676dd982b0be0249ad01e2c2b40f22e38594bf7a16a782ad3372c74c769a00f2db5c17807f4c3ac6ab1f4a9441623a34eb766c374160388546dffe8f35b0297560fb6352db5b35a313b99af5700314fff6c92e116980ba1f28c9997b31bc8d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2101def5cfb55345ea0ca92277ed211e37c881c569e8a7c2597dc365fbadd69af666134ea80c61385bbd5a933faa8d25a2adb0dd630ebfab0c5aadb4918f92bd04a3d2baebaf6a690c85918a9117d31abb56cf5f3796427547e381977543ebd4194f473b142dac244611d1f0b67e4d62f32ba7ace392f9fbafde199ce74a1455;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf4b7a84b080cf81e0c25f8f9e918abae14e0e85c788af04f42fb24f1e16406c8a5cd2da3c8df16124bcbef0bd4569c573169fdb86fd8aacbbdee539a7fbb4f37b625e7f8d9c278f0633089023a1870cc56a54a711ba16436c624676e134f15ef2bdd7f1c5d5a5ba6afb824271fda9e5be17ec5c5dba46bb86235c5aaa6936a88;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd40a15130c7c3d025464bce7bddd41f89843585ba7093f56235c239f3e51505447b791d353769b58428693d82cb6a57abaabb00d70948e510f1476dd740f6e2e397ff9963c70555ceb65599df6ae6784022a9ec345d2d749b3fe7cd0f83157745cdb0a9b0406f903c51324d715940a34ee47f740d97ed207b668ba54e2dfc3e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1eff9181b64bd960641ec304940760430fb2df2a7fade0323f80917bc7030db462fcda1854ca36b788e7fae14653d44e249ee861ff876693295be7007a015f8c426896df16bc7375f5e6eb03dba58f4a700aeb61759e589f1fbcf160ca54ce5b9d6b7f212545904b86db6a153d0b9aeb628ef6dd322ff977d538487e54cb1722;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6cdd9ace5b54d27f44f5aa0f08b4d0c9a88e02dcf807ffae2aa5a3a4d81cac7cc7bbef5d404a8213fbd129ec0b978e7986d4f339b5ddcd9738191c8fbc3fcde2916d48018bd048d6300e678a7ddf76da8ada49eed30dd6a3c6c400e256c220d27287749203c8e7b6e6721e03a1541d6f02136966f609e55344cc52e72c143bcb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb499e4933fcc425c4265e8252ee2a535d82f743d0d2b6382a8c25a8dfdc35b2211cfc6424449cc9b3328ff29a6ed87fa4cc41de8ce56ca90adc35760d90a5fbe2f3f2fa5355fdc577eddd83dc4d5734e18ce8f641a6511445a57d1ad32fe397485514379d4fd93bfa4dd03ed019f544ce35f0ee89d929f512d71a3635d7f9881;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h271224efa3e996cdc32c8234e6c7c234fb1dae12ae0225d142d30afdf06062a43ec67e8512901281ccbd6c043ad9d3c794095bf0d42424920510d9b42b527cfc1fb94900483eac362956f956f22707470435046073526269f4e5e0e2221f6886ba7c52d826f5b5804dd42eee556b3d346975ebf3ce9d5c6fecc841031d61e87;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85329c3bc5ac18ea1a6c04835cb016a009391bed036c6ae1f44c02e84d9bb80551684bc3787638464915afd3d4cf89818168a01006c42f782079e1822bc1793744a4d967114bd85d66d079fc18652ffa860a65a3188de060ea6a0d2507a58c04a2515369ed101f534703a656701621ff67e473feebe3d7616f99e78d26d69959;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72898f157ef4d3d52ae4163f371cded4fb4e68aaa9e6f9d4cfff2adefa025fe2bd8feb8172167c879bd5c85de39e53eef83dd118c80cd6e5122b99481d5d6aeb4b54cb3d21c82ec08f843b07e03fed9950340272a10985688fa6531620d1294f64cdcaaa2b2e0556045356aebb8980b6b20b0aeb3a8b502a9b082af690a03a03;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c72c802c87fece305b01ce6e419d728d0f0f289311ef7a6e5961a9056a493cfc9428abb6ac3124945cad55b702a6c2f619074d65e275a971904207ff25afd539229466dd50ab65df60f9614652ff061ff016fb1023926f86a5bb8fcde5182acd589b5ccd637adf585a8c6888aaea6253e8f8a3618aad3c563c87b014cc04a9b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2303455b8c8de0ee8586756d57fb1b73cbe53c198159f2c42b7e048d90855fb96c0fff17f3a426373bdccef2b8f7d5e80068107d76c639a9a307a7169e9bd381f3c3bb759ac7f1fce86024b70679603784777496bbc9ab21c56e1ad76f7fb7ed70e70ed20336edd8ec85683f89d27c4e00f1817d0a2c6cd065c3210b016c43c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22d44f1f86f6c39a905cc3b0c124a06a85fcc3af1dbbc3cced96b2e3a3aac92142fcd509b4bdc4149f0f8ce790e483cd29078b3f54ae9cfdacafedccd09d9d4e39a87a7a420bf9ced3d5674ea17bba06e33ae7cebab52f3d215cbcc1517cf29e7c81d58a1c67b05330d6aef9d9c34351fdfcf24c3d78b519e3e393c3fa148be5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4236510df43934ee238648f36a4af168abc86edf5756936765ac8519551a1ed5bdbbc669d9f083ebd532bd5eae38b6e016980b25d73d866490b942bbeaeb4ebe0f6cef1810fe7cff5149145cc6334c655115afda16de54a14659562f92e6377fbd75a4c0f61b4a56c030a0d5dde492964888a5f05da3402116c160bf63c099e8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba7dc66fcefe3f55be62cab952090ae05e3ec2571f7618e6d9a2971e94e21757c8ca3470a33beae4e0138d45439579f571fe0ba1760246afc4d50980ff2b2a9c300fbedf240b0b79a1ae0a1ad3f09621c98470f40c86577560b21c2ddcf3b9f1f1e02a44ccf0fd3f8368c7b5846efa2d5fc095484255df8cdca58c111c496d19;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9c842e7d5057d599588d6b2f9c3f2b973f73f47efb388eafa684c8ebbeaf269a29a279a46423e31f57b76ecec09281199d506db33a7e1e6dd05b3e0583f384fca09abb2ae7a7ad8b42747fa3f42417f0eb39ea174f3be4748ce59132ddeb89f8b3aa9d3b93dbfb6425362c69198f174aebf5b07546bc2562954577f12be8b3b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h318d81b57199f60b13746084dfe4dc5472923b4affdaa4af13b4b8b4746ef8bac6d1d247a0486dc2e2eafd65f8212eadce26b2c535da36d9d83676190ba74e679e12631857a73e5aca686abd352d4ee89590a0a88b33dcda63d14a8167495f2c0d2176e09327f97dbbdc281ea8f8112f67f8f5991cb7ca740b49540ee8acf3cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h654f4b2dc3e540e7f0d788d457898471820f3f2da593c59513cde0af6eac6d349805433641be9b6a5ede95eb46134fb4879a7535d8225541e23a66d57be6ac0721c0f9bf521133ed8414b59503de433dad09205b211b12b06097523e7c3aa26442899aadb956672cf8d5778b066f2b08c441c40d09a6551bae12945b72e89444;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he06dffa936378bdf91aa1d7c996a5a0fc57ad53778e61ce8f57c6b1accc5565ebc33eee741059bc1aa1c906e4a795938b7019b8e1f24606f639b048dc93ee943807332a87218ebe11f677702eaf18d89aa482da60ffa03461f1ff05119052376e2e3308c672483eafa4110876253211be62d2cf487d6bb0400f5b001510b0027;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e828e2cca33870f96ce00026edeae41a1425123b9ba558aa925971f72495f2405ca876e7659421884026949db0f82230cbfbc2964fd3194665e7d85c7431877f145f8ef88fd792cb545abb0f68f3b9437f03d286c37563a5106d813e3026e55f0dcfe6a3d726691f696653a10bd176a9ad0944b9eab3b9526c349c84aebf266;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b04430148f289e38d44ddb377d776c54517a0401cff14f1340b8e7e7de9c24a9bfc400c5e0baa1cc425429a236af70c015c00add37f5c5b1a26c111c8d501200013f4222c467cca82e91e41feeea55c257ee0ecd5957605e3e41684093e7bb399c9eb0ac58773cef9c5fff86c121f807840d5e33cba1e78044fdaacdc368a86;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h815062497b55965a64aef7191535b2811cae48c57766d408b62d0e1e9c355f4bfe9e0d45615b92cd6520286178dd6fd538186ab62cad0367e9aeca92702f2888389eab6535e7e752cba1f2ce853932648bb71b3398ab6de2bcc8b0ac511296da67a15bfc554aa081ea89f2d42b90f3f3a82541aa3b7f7da4a79830b6de6d80f4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h651a603280b71389da6ea8c24dd09720266a2ade73705b8c7101714ba379826adae02c369cfe861bdc51fd6deac2d66575af901ffccae7522b35c076f496b05a9409425c51940889d8e8f1f3981850d0be3fb05988dbf5eecc10d8a35559df4c190d31bba4f30457f028d27ec0fcf2fe22925203179423da52130e092202a59d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac79888863a779548719db2ca04bed017613395e7e7f84f9a147aaf77f67bc98f4c5ab3195f5dc908a515d5941c1cc61e8b656454f8fe58e9460fbae9546d0b86617b20f4e31e39a3b253423ccf63008455d1c542907e2f291df4dda5ffab53adfa3285ca5a4991998844ea0bc8c09a5f640bf51eb96a42102f5357c98972bfa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab1f65097e011d14a1f8e37a13be6a917c848ae07c1414276043ea9e411118cf24b7737663b7e407ff50ea0cacf59ac033ca50d58b6ada40b11ca9fdcfa0ae7520c8371d0174c12a98913c491b5637e3989e4cdb0df6d008560ff192879e993abd12929174dd784005f47cd0770aba72fdb003c2eda1149a5a8861ecd4b0db3a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6269ac498c92a7c7449054433c08cbc059eae9dcb002654ac29c0fb21d5c1b1de05f4e7c372b7ee90ae87b51fe4073dc8865271c33da64e01f6bd39b623e4c2f80977b68076e07a782019564f6d8f6c605257946a0db41fd5c04b79046617e304812bd117423090dcb1d0be04dcf7e3edeabadd6b20dcdcda4ff2e4d6db5fdb3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5cde5e0daf74a5b0e6625b08e1c6c8340183ca7f2858f5c4d5d0ad411931be8ed245a8ebccb498d839e5091e1a4143fdb3434e2e74feeaf36a66328642f37d7bfe15a3578cc4af4610b3eb9df4ae3793623aadd7f83e2eb340000753a7feb638777964a72a2af290b3fd5322b9987a83482a226f8be78c481b7926d711096a02;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf068b79c768f6be6fe3e5178920455efd4120289b8a1a232dda0d04dff0ee5e9fc57d7a874ac132f82edcef21c17c1da24d7084022ad3683370c557f597dc02a7ed1095e9466d26ee7d51b45d3a623f7b31deba7161bd641fb47bb8ca82fbd5da90254355a57135c4987f6bc19394af4b33794e85f325966bfda8acd614440fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc17560c1b4c38906d7c44bafbfbd4e34eb80c44c27d16414507921c085f92688ad989ec9809556432da5ed1b4574e9967a81d5a9b015b93fb5eedc96e8e678ac7aab411bbd203d11b459fd6841dd2d65c354ba3f16a5dd73140f96fa83c261841b841f31f06dc073abce952a6bb7255867377428393e1f2a74503b251296d80;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb7e16ece2a2b23bb4fa6997308525bd6fe251cf732a92ba3092b82ec56df13ed4be3e22ae789c2a41c1cdfb69569e55771009a4a59e3e0f958c17dc54ce671438c074dc76fdf957a7e3535aba21f59d1bcd1ee6973f534737b78e22898acf011efc24f0f5bbedc0f8b8e42798d8f8ceca7f3b266df780df06ccbd96d9c183e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd66d82d3c6e34922ae969a150b144a3ca5cc99eef4737c7896aece1cfe1484e8fe569e44b12755abe4afd2b47f8a7b4232778e4e8348927cabf7f68bb14ea06ee4d2f72054103d7dab289ab747c9dfd3bb3877a22ce005d8f1a0601fd70c3fa6f509ac220224bca69aa8793d83aafec429d7016ac6d5fed05bb1033925607d5e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18b31cef7ea0417c09c20b7860f5b9b96f962433004320a0318cc3bff5796a797e7d556ff1803dde256bcac6a2d440e1b572d8a612c43987b7cfc93dd304d3645c126656fca4d3446362a7a614c1320748ef66aa2def658fdd77cfdf7f6d4566458fdba3b265ae90e75038248eecf8ec4c1a908be5fc1e09526ea02336e08cdc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42ef0df617093b81c4be69eafc03f8db14f1f3510dc81da1d10645dad7ebe8bd1e999337fc17587aa1c9f4260a8159ad493fd1b582029181204913ccaeee78fe527c57d9072a318f6199b9be2b85e5d3b7ef199d0c287b69073e1fc7ec3515a45bfd6a6377959e2ba626247aa03e6df641d676963539a7e8bc50e4e2e3277629;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2c190defa94a92aafbfcc19bce94525ca26a74c19656e49f900132cd0be00ddf966d6677972a80f47a759a3ab019005e3bc35db1113a1ed0a9d41a496b4441e76d157998892c0a23327e16c186fb7c0936b0e81f881f371854411c4842b71e88eff5f81b20889c8ec1a4a95713200b2f16d619084dd056b28594aec9f467744;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha98d9b64c37c3ae32c5b7976d238461172fb8c7e21d7a77df8e4d4b5b6d7864a34c1d2ec9e110b15b4504f5b2559e420452ae3c9233973a19d58f6e84ba0f5c25df74dee50417748fbd7309ec77a788643998c254304c35f8a18bec90ad702027a0dbcfdacdec25300736a89a350243a58d107ce2f8fe0712d0c6e3919297cdb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2652c59b8a7bfc01b95008f22bd6c509280c09001b8d83e72f587f937fddd147b3aeefd235afd83cc1dc3313f4172788ed8b84fa4ec6cfe513bc01d660db6397ab2953644cb1b6bd081749e131e277b8aa0b51d36f7dce2d67c80c7a5427b7f2d15b5e324a2a31ba80fc81de7a68749dad6f58e153d2ece32047b6cf7c0a26a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74c6fdb69397634c7d0aab5f864f341e243cd015f16a9d5901ce675ba57a12a360dd483838227f20bfa47176e9157d5b068d0cc2f6dbccd4d7f3adc0c778075ecd6e4d27adc75af8892b17721f2a07c33aabaed0f0cbf1d82087689b2a9b6aa26faf7c8dd53916c7bcdb195935e313ec1f20b0031da243c8aab2aa97b5a512b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ca853f025c5d6439497a3bfb0cf11d9bc680af973b11e674e61e9275bde8fe5151eedf6fc9b21993776f6307919ddea1e7c08b53a3712f1c8b093107a14f4c2e51d70ae6ed8ec8cae661556d1a7a477ec8693287348536f644a284e0560e20aa0e78756ae67d7e2e4253276257bb512478fcc62e89d953df4dfcf50896477f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4e238ec25f8cb6ee3b82302bfc1a921e73d9746537543986eb5bb3351134fcf543f0d49ab1c3edbd8e84ede2a2dfbf1ba0085d1e202019b3c64cd908519f32fa663023effb192eaa7a4f55615fd3d4767282da3c7f2cdabc78baaea7b82b11fabf080027f2fd56ccab06df0e74919aa99da4a1be2d7121cbed09e8c78e110ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha28ef7714f19e5a12e63f8bf7d21562d07736fbb3ea09712aa60c3f1ca0ab793fb6cdd48f54fae735ff6f2c9c0fe163b8f9dab434ca2f7b1b5daf3c5f21e3ed83df49b99c16e0a93a83e5e888ce86d1f71e64f02f3f8ac2cf704d59927e3ec6dd4a1cd057a2a66caed294fee26018de6c564daba43e884bdf4fdcc4b82ee723f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h783bbc4abff72b9ea4b64e334e12dea459e2be1725e054bbc969c2c35f2cb3842308bbb379ff0324700f69c5fd8fc6cd3b5a12e80b00cbfed89cec76be6849ae6bf811e201f6a2049ad57d6e05eb0d6857b307b984be1fd0ca7d05986f1fed95fffff4c4ca0ca05a2a6163aa401ad01cc3e282fe1833c4c1674f5344a665fa2f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he237b46f19011a11860f08e381563f5f48c38314803f322d07a64e4822e4ae6b985feec2d6daa83cd6353afce25a559b0e03588260a49832dbb8eb09f482cd4a74118d9ac08508a39b3cc65176a41d1542bfb19ee51e4e067fb12b4b868f23f43faf1a3449c6bf6700ff636dbc1b4b757a7984218d7c82149f69fb372f7518d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91efc1c75c6411bb1e1be566ae0248cd947c3635aefbe3a96d3d5b91d365f78efda78a4251d1f3398ea119c992278cb2217b6987c7594a231c7e1e17d231dc9d934e1151910b87cd70f5cabc633fb6bf21977adc0da62be52e3bbdea4199713ac4dc71fa449c7f98f2936fef4de8f93da5583037414bd8d0124927c7012713ce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee7ca216bfd7b64f5a74a208c0c678a0be386e55659d2967285f1b0204bdef5ca1a6328f32954d1ba062943dff75530938717ac3a6b47c6da533a4acd49dbb0ba4e7e91ce1ddc0c6689469815c4309b0440127a18d4e652cc237db507130cc02f5f9ddeb343a6cd6681f80a60400a966c3bd0be829862751e70eac98d9267c5a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19711e99db96f83783500782a17ca8e6476dfc19b6c308ba7de6642732b2104babcf859b2f7d3e5f3f451d3c2b1b6227312b641771a9e973827922d3e111b4e5cc54bc9d9f16ce516a665175886758b2576795164c506c8c2d8fe218482a7f724667147b83d909d56d734fba4b4f301ee1055693214d835539a55f58a68d545f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h874e99273f5ae7f2da258c5c7e9866460bdb4faa1cfb1bd63cb2c6d8efd2bd268eb2f9c3d44f2e2b79cdfc78597d8d5f2a8831a4eaeae3b8788676ee17c17abbc7ce029b277e966c24876c0739c1f9bf020341331932aa0c869e89d2dd2ce1c7176d9f48fd0a39e9a5d0abe8dd341f65b9977a7a35bb28b632c0a5edaae16f54;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4c34318d9ad1bd319f20f32ef2c11e8d36e93906c2fd548ae1c5d4c1374fdf6a09d9a535a15dc24eb1d3c1b54c382c639b4276e9daf5e44696100d3fe69dd81e08320d04e3b9c9c47cd791a6e87bc4de9062fa45aad154275ee3dcda88f6200485f7864386958a7e7701e1699ad2782231cb102ac98d031bb1efaf4ff947d5b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcaf3bd071f2f7f512b53b929896443f2e2d6d4677f027328babc7c233654484a1cc62d3a6da31096fa40b7ba576b72f6041782d92bf9f46173658f05a26bb3e2694e131ff119d04abf01bcd9063630daaba306b81c31444bb288e8af44508d6a1af6549a4cad29a3b7d675d0565119a075a703a4aa1db79bc72828415dda39c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h29a1fea1599f82aa826a433fbaac2b83b2f129a81adcff3e2c94525a5f78ed52027b7680a83bd44d5a2ed382615ac93c5e9baf635ca844f27ee12d4bb2c0a77999c10792a0329894e0133ea087bd2ebdbfb818b650f1cb92a8145841050996511cf7d67a0e3f0656d5be7e85908bb06e97be9afe76246899cce8add059971e5b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h90d4243dd9fbee206a8da63807b65de282138032e6b9a3b7b8672a160d6797da98f34183327df6ed31ec484d4168bb8ce9d25a95486ccda89b95f70af4d5ec6a0975fa803c1fc82162aa493f8b1203a282f734f8b607c6fc727b85898b93617287fd73401dd2338d11a8a0e02d4a23fc54a2f78dd062fbb881d8fe2a73b665c2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35f994179bcea350f85eb36ad58aee7eb1aa0572f370f40724bcce2422176b4f74d5f3aabdb99964292c784146b06c3fc08d52c2fe203b78fb8067f1b209ef93ba298cbe762e9b5987d8066745588e136f1b3b909d35890bd11b118915cea43865b0c20184b8fccb0b709e1cb3c96ffab1cec3e2097e010d940ed2c148664758;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec372f340a37266489af2676801ff828ad8cdfed1e58510ee64f4570f9eac3890499e22744343cd56bd1aef2e8aab499b305ba6025f0f7a0815b89bfc509a9595a263a9bff2b42cb7bd16abaef3a21b42f6a5eeb0f50cbe8d92e1eb60ebc43caab52b983a930804996c2db3c197d7c80334da1a2075d1d048648d4b72fb3c3a5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdaec6c017cb85fe75f12c68467a5f9ed23934cc98029e74dc744e96edfd66fa02878648e56e7bc327e8622e6abfdc0d5336e95b82297bbcad94d0fc664cfbf14ca2c8443e3aea502ea4b76b14d4255c6bebf4b6eacdb941964ca8fb51f0ef37ba8491acf4e0fc836920c2307e8fa60aba579906f277d271547d0130a179cdfc3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97e52d78039f567d0ee1da2dc229aad26822557e9ce5d82676b81aef0b3b9bf62c1cf1f1de74e9e555db4022ec7cf87429e6eb0819fb698a2fb56d9867438d1138a6247fa681b66601305f4a67bda3be267945312c24262b60e5a0c420a97ccdc84716f8e9c21eb64ce1c00e9eea451f9dc05c6ea915602faf1c1527fa27b937;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ab63b07f66f01e9ae5bb82184dcdb8e3ba91f54169cfb8d71bd18200efd1f7d34aa45eb17e4fae0aa821aff580c6369ac5097c0744ed72cd88c1d6b6c030d56af9cffe8fb1ee73db07d7f9b9df9771af76426a8db1c5cbeaa028de7859be9e9e0c0fdc1b895b2271507d3be0408c8a56195b0f524689a52097c694d6959c7a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h448e03f9ad3738653f1c9285c3f1ad2a152e88a42a8740143af8eceebf92b9131d19e1f93c402d180dbe139d99fbbe8b46209f3100df5ea9fd37038981f9a1896803cf70b37626678a0a914b8c3ab652e5c5396802319a6e514451c9476f3278f504facd6e1842413b4442e32a1bdb0b47ad46bac73df9573308701218dbde7b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h858fb261e5a42768d5eefcfb8be3b51a83832657728cb2d1494483158d956dd67343a1949f75fb8464d09e9964c8ee93d869bf99b07018f0ab66fda3425d95d99f1b74c2e8b3de6640350598043712541e7edfea0562178d92253d514cfe920bf564a8138655ba95c4a7d6d4c01774e0237837dc571e27f4f366ac35ecc9e990;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5b89ba7969936c9e5fd20a5dc8e1a057e03073dc89563d8d707bb9f76c2e5971fec87582196c6fd85fdb05669d22c7e0cb1d4de8384152f1cc4112cfba8e67a44dffd70e71548b0ec502c0d54f396784bfcf7bf97d3a8ed582de7de7e3677ee954ae373c732e70fe1356557ad551297f32c8fdfac1610a5cad8dc632281ea85;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he44148d38125eb2ff33f5dae26c1f9adaa42962295810ee88d6be7ac5a4fc83b0558bd8e22bd948d45660fe2b606c350b7a683e845dd0e9363559c44b4e863d1eb7e52e40d7c40aaa892bcbff476b3f097569b7e51f888a1e8a29e3df693f89b438cb0559b8898a9e11de9c0b4a1c6c005bfec0fc2a71ffadd1c803f05e5aa81;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28dec7b82015fa5b4c12d5ea741493965d2a0f4fbd6c5fd633b82a67f48f4680f7ffbd24e3983c581f0ca8589dbc47bad1aaf4e1cce850045ee4d08aefa9a549a73dbdb9bc2cc033bea56985a7fc353cbd7dba1779f8f17c9fc33f87bd37354fd2a6b138d392004dfe3138291923bff12ed19391136b64228dd82720ae709327;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e7240c10e916e5216e0d29fe953f75fdf019177f216983aa6e0ebf8408147c5669b9fb8ebbfcab1d255edd5553dabeb198cae2e1dc2001661c0243ae4bf639a2a59d7e5bbed1e4b892bb5ec4598968ca4b0a885673ee27ab05e0716c1a8d82c9ba46af9d7da5aa59af817d6f9d4a5456c72de3ec7f910b874f81bdabe2f6d36;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b2dd6002b92fafe319f6e26bdf1c6752476db711eac15dd2fd50e4f2b5e1db926130ec82f0b24aa049e82940bdd793c734e74f9e8a341a01f8505e410a029f9838b7e64f9fafaeacedacb1b737bd27f18b8717dba97ba55c127d8ad530207562ae8f72e7ce7c38553624b71299ff9294f6291479ee53d7439aaa6e01f39fbf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde5e758bdabbf12e13899d1d519b02dcc557c91d58075458092c0b5bcc39795dfcb9523828150f4ff03a198d8dd9889c48dbf9b9341f62204a37881cbfa9af29b43f03f53695ec2dc9580172e27b007388552d47a082fdf31980cfb30d903daa90f98e694debc935275d5ef3b53da556cf6f694d3b470c2970fdcb725d1b2eb6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf64787f0c30b4eba2e68e676b5250369621b016368fb0265a2b03f8946e076765fccde0da9729c439b4f124d8f21ed0e12e9d8703ab8f033ee41141782a51dd5d3e5ece74594c43f6429a6cc079d7cca0e4075622ba02eaeb4ef75483518f67fc00b06a3c3734b302e3b5a1b0ce64b26270f3b07a50e94ae3f2eb7ccd7af7475;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc4159023e1a0e0a4b5943538e61584838e233b4a061f0a769c8dee09600499553a613e0f480e8bc2bb52ab9a0f6b67b1fce494b43ed8eab1ba307bc5a2c0bd47cd6c0ea9588056077b7768d97da61ca5769060fc57d250df2d4520f704bc54dfa39f06cdd7545229af964f90e08433217fb2ebab6048ffced32a94e3bdea7e5d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97bd1aef2d078d36a299063e05c0b641df00086e326cb4ff458fed10e7e9c0b8ead1b445271c90d4826ce1a19ef052341f68c6de56d4906d30677565cb60a9924ebee636e174c02324e09ff82ed442b6bfdf71c57ac5546cff84894b74f125fe830ce9c68594f8e576a6e75dd06d538c3c0275fca6a4b73621abdd340e92967f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1810d433897badc0d4b7adf6b8d532b04e35185537d512d0b228da0e053cf6ddea981d9fd100b64de2003d44ef462a84e5eceb0ec04936e1bdd1802c98391c271ee6300395af43edc771b876ae94c3ab17a92a2f7f5d6063a695f5b7477b87ff6d6c020e8da80d3b1429f04eeca4ad054f38dc709ec117a8159e8316715bcf68;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79cb9d07acedb8c42e4026927d9b63afd49fb6197a2f0f30d9accf7ce13c34807066432432dc788562617dabf78982bd6e8c170aaaa75e7aaa45d01800cdc1947f7daa15516ae4eea8cf5ab3a60a8ced65256c9223e8527b36edee2aa54f68909369f8ed727f38bc2c41410890fa7b7ec0f1d7cb32a272ccab16adabfda823e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74856c2157c6dcff20d30f98c50e5a4e2a1b2f1b43c7a6196336042c447d6d55d4c9246c31d8d240446782df36d7120bc26606deb6f629cd3060abd8696d11ddc0ffd322b6dc6667b99e1962bc975fa853f6649f8aa61a4946b01d20226c9aa10a689b50d0442745624d84b665cb6508ee3776d0236bc7cb880aff36bc24639e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9cc64a099fe7cccedd935948daee6f05c639780c53bb0db678e7cd0c9425f62dc3e8e2466d746dffbf5a569d6500ceaf3fb8c1e6b5b970e29ae642470e11b6d5316d398357cfaf725218eeadb2eef13e87d9aabcfe5283270ffa7c5e901e3865126edd8fcf90833eb3cb4198b47474b50383f94577bcd279f66273745418b780;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c15f84ad5d88202bb64b619d6fb7e18721782c997b18037e4eb3780f3c52bc8810f9c38dd961b3b4afbe7c5739d52fb9bc78a21a9f3f14b17bfce7cf9169b554cd0e3a4210a00ef9b4b2463c05c679d87e6c806a5d02786bc399406e7101b55046f8441d7326cbfec58d69d4bd5a6672db5c00326506c4badf46de5d2054790;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf64b7d9c56c5e43b9b8fdbe9ff17ff115df4b810f3859fa8458612dd39db331d883149f5fc1b72dcdb7ccd4aebfc4327def024957451c74bb6a24c464b4ea9974deb904e1ff03c0a2e105cb631badf6c54a5f21a5b64fe14a3dcd1fbc6933d4c4386b93a7d0d221b74870621592822798d09a11768d5b81409fdc7cf5e224937;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb527b04461b498bf24d3690ac08d68ac50922b3426ed078fb71e8b388395390d320e8097bb07f074c7d73ba9f5fe8205bcf162c7b178bbdf84285886db7ce31d3ac36557fb31e15a14154f08e5efbe3b8ad0ed01f686ca9b0f8b92716696f294e87e53f1fdf62e1819b2ddb04b41c8f9d10c34c1607d461bc6b9a25e2daac9a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d724c31283415db215a145c36aff6c1830c9edea893d0a19cc0178b27d6a872b0f708934cddf74841dc369ba50e37914e43f388db77513707346763948b2c1cfde5449018ed5153267ce057c2c3cea2fb9b46b856764cdaa94a155f13b2ffb5e3441a9f455b1078729e5d3515741e88176d717e7bc95534b996cd7eaca0f99c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e67677d828ab52c88c2e7859a82d90973173cbd7b1104d378c85f1d3d5c938451d19983fd7555261c217956e5747871d6d17e16dfe3fdfc830678ef93404d929635c9a81488d743e7ea706f76c24851e043327e9639f5d70dd8124e30356ec4ff72c72592819ab2811623a04aacbd8d4b7aa6f602d194bef7c6d686d4b22fd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9bbc496b96d6d8bb01dfab27b6705f24086002b8fb967e51a5448aca66a8f544f7ef56a43fada163c9d1ba238a7f53d4e8adc423d6b36d0959b32fca8b51375f058a333a2d9560c7ebcc0439863e98b1c14b257f877fc7166b65bb2d79806c56da9c7fa2364fd4069ed3887b940bb406cbb4a81ba4bad731caa06e17c539e00f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h645a802f6efa85669d0de5f16aaecbbae40a554814f6d366abcf0ebb43233ad3f58bee566efd55ae2d193878bccfa732cb9a98b043451c41c522691569dfdd31e247c16d13b44d3f4f2276051ae003db332accd0f2eca6a07027d3df567117ea70b400b18a1beb95968a5151762dd85d8be27eb4697f02945792f9e314e13f5d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h250c0eed31cef7d9557f6da393055115e874494963b8714d78fad88b58a8a719b73d9329fca7a808d316b3e5b5cfce931ac9ee2a8199bad6468688822bddc2c6e5ead2ceb2a3e4059d7797f088493ddbd168a63cc25359d125334ee77e063645eedf441087e77b1d85645be43510e7c19de996242ad61a24833e8cd7aa5fe5c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb50bb88c28a810b7f096a9bdabe80e6e8585cc3c22fbc8801b5123e13e5e7e278bd2c81250873d71f627ccc74cfafb59aadf6aaa59cd853dff15f64eec2aededca1436b998fb11dd14b7df02b886d6c71134e5bf85de50cbb2c3eb620f99bf17ebc5b1b2654af6027693a9adf6e6d024696d6f08c6af70b4d4c0873dae7571a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7912f9f0d991f0291d7a04a9d25f83d555a9fd44503778cc387b41ccdb2e2372e5204d3047945ba6d746d87ddb7ad8c521a1659792706d7b97a78e6a779a0bd4eeac2ce35064e0d046c2d12b692732bdcad0724e64ad8d0f0163110591812b57e3442a0bcd1356f6226a38adc2c7c806ca682e5c11e841587e15eaffaea5bd7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8498548714ceadd26f6a9aaae031666c8d8c7bff54a2d3cf444626d21965ff65b5cf26ce902cc248fbcd500d2d68f69c06e1f5ea92bb0fd5b92cf80e5b7825cebbe9f1e7954b5c8ce237d26d7989961cf41d8504461bf8e5c6698bd4afbc2c923442ee9d84e53f297e4d9258b05a03e2bf2c393bcddb7c291ce8828fe83bc56;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h376579b01b1671ecf5f45e6a03951f77ff46c1c7c823b8004cd5b581ec31c6b6d44cc45faef05893cec61f2131ed2a951328c500688b01a5be77016104490db31376aeafc26c22cef17d8655cd5f9388a4056c04563439a5d4b972f876980456c723370eba69cfc0d6ceab878c8db245eca2de8eb58dd79ea0f62c50e678ea8c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h593e551b0fc57ac3e0b7c79c25bf1b3d6a506af2743483c79aa76798662dd377c52df84c4253171736aa38c08a91710961dabbe0d0c8ff900932fd69b3b150bf60633442d16f3626bf1edcf863a41a6197edb232249810ce8ac74060caa77c02f5222866cdd8d1609c391a273a36fe623e86a9e7ddaae2da8207ac91c318b731;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdfdc31c3433f68d4d07b59f27842a19b96f6caef35235ac7ba5bd051c9e782fb01f329609b3feb144087b1cec17de17dbf238170bf5d155677d775975723cf9859a6e439673a4546a68befd67181b126309ee6f7bf9ec504e3d1b70e956af23ee8ba4ef971313f69f00b7949f7c342f94045b2d82d495da6cfa469d5236174d8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd78f5446263c2b0c69f26e5ccc0cb71004f89f22edcff4e4bce8022cb924e8279d6da6b6399fee864993e80d824416166b2bf77057ea87b8ade5dbdecbf9df5863f02d02f4ae70a768ec38c3b456b2fe3486801d8fb7b8feb5f2592426dc1c7d2e891292c7433e2238b74bf5f4b42cd6be7831d7e88e7001ea58b790b09a9964;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85a07597c1295496c5fa66c0eb02939d8a22e11ca46e47d06854d14ee49a04e32b8604d7d227504a58adf0c0f53659e285edf935bbe10af1981de862aa910cdd1e0e4912e5f3ae6d1db5423734b3babf0579fd7cef44257eaf7f02687bbd9b69e6e8982a3cc0c48024b3bb0eb30842c1cfdec0abbf5955d2f1b2d879955a4439;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbdbd57241c384650580716e32cf2ead78e45f83e8e0ff50a14d70ef4183f6153441e61d04d5213460197e86e14c10c7e337b6bd10b7346a036aab1143efc2a6cb52e16bc2aa8cfe41448762810b712edbde469385eb38fb26a7424d13a9fe891547a7a81938b3fd7a5b0e2b33d750f753c6891e2b903bee8b698ab7c9790a49f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd41da3a81130e5423263d40be767bbf17093d408683fb720878177d8ac04b30ad353b147d3b7d99323c14d37ce1d723a2c4b06884a0228438a522e820d86cdc2d3cd72e1f7e7aa0ed80ca105ef11bf542f1c65e91bff0abd8ef74432c2e0d535b0fc7a633f15f344c5589fcbce81fa4f868587ff140f33cf2aa2b05f151a02c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5da16a6588d7b52fa6fa807c3559b02a34723a7b02a41d2d99b3d3e44818834906f8b7f2ef3e2c4b3a91e3f60a338b15fdcaabb9795b09f30c93ddefa7b3d70e7cd8d8c14797f3fcb8cf2bc713a6f603a2b9107ccc0ea3dee2e7e0eda43172b1a3b24606e007957fa55df0f58049014375cc41816ef3bdc4531dd7389e10bffd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h45e0d1ac4bae037f66ccddbe13cc6e1a43a8504189d23f014f2cf1b7497186096fe4acea7248ea856cfed0e1c79e136c1c0b767cb25fb23dd3a0130d8be8f57dd4882fd433ba6714a535161859cbbc638f3c298b39818f9799e0062e0e56624ffd1abcf8641a67c7e909ef8aaa8f7c347dfbc7bbae1e8d06929adc349373f26;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4da40a71c94e7e01ceb7d291fbdf9d9ac1b9bdb05f44f8aaab5a32a4d09e0c4d500d3c408c90aa402d2f57e77370ca4d0a6ed6d6c4bd673cbe5e1383668321e76dc6e99c967016e148b4b7fd1b7d4466c91d5d07c914a7621668150623976454b5850fad0a242613fca8930df37593193d174b94e368a3a62a09e7e411b14666;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha1210cdc44d5ed35cac4ad7e9f4035b526dd26f9caee479d99dfc03cf9e4445b397ba10112e3cd5fa60b50f308f6cd2e3446ce2e9673322ea9439427bb963b11806f498ef9e9ed15709b8e07baf077e272d1d4362c0ee82aaabdec8fe32fb9f8a1784a1d36cc02a1af236754c3f473fd4b63e431ca71e2cbda7b58f1d37458ca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34f4cd315a2aba3589fec91e26dfb6c1acd743a2764b71f9bf38f59870442fc000e18832db3cbb32353ec712ab6a8a7e7950ad272b26e34cd0e22389302fc469162489ffe9c4901275b436f0348900f0586b2a883d6c02828a3b30f3fdd4c8f25e61adf43afd2f130273212edec62f509116b2f68f501cb857bcb2474f1b9314;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfbd90e0d9ffcef6f1cf5c4a5cd96cd909e348f1d70714d6dc37ba2d4ed7a08d79db8d66e62e6d8039f8be7dc410e163fdc25ec965f9a0e86e5b186d4c1addd4b872269c0b463e27a85a2253faed26b2117ac043195f1ea0b8db8e42b3ce44384b6b8b85de324352cbad912f91f201bec40e4e5f4a42fcad0bddae0a5f821450;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha582fb2dfa361dd6d9e1ea4e0ef85878dd758cf590524d675425df93875d98cf184de5587a26076e3643516e95e61d9b2c84ab7a6336b148ef520ceab3ee49c9abd6aac8dee203da23a26026d91cbe1f19a8938312ab2afebca10b864580c8fd79d5e9df64bbf01287f8b884d8757311df3240f193a56cc64cae4ff5f9c2240b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7eb71c6be34141fe4cbd6103b8cfdfcc493345b118137f3d8c4772d80b87b568da0dc7c14ffaf4aaac37be4df78212a165c71dd06090b75ed93ff53bc38e09ad0799b9cb8a6797060a035b337b01c9856bec7045c2fab873a41d29004b86ba7e5e9a57b6df54edc25deef344452d1a88482d87ff5ed8d4d99b970fc30e6c18c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdbf9fd9db450420881d17ac0aa07b080b42b7d34ad6927436a96e3bb02538f58a93bf1fa2ba6002a5f9fe83d81fd8223ad86017d6dbdc4c01e9e3ce3688f35a62c76fc6975c2d2da5479bdbbf708a2dfe290d39ccbc35de12966596ee5859432efb0bd83007097c102f5b6fcff19c4293e282ede66cab7624f25a9811e3e2538;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd55af2e2d1f394d733b6861edabbecbd90577e83d0dba476cfa4fed80be23766a8d77ec6538b1be80ef498d23f965a9cfb1c6e835a9b64b531c13308fddcb642adf477a852c4fd1fff3187feb8e2b092a5513e10a7b2fb7a0a9c34520c4a0dfce9310bb579a1a632e48d8795d87a134b96c8c87d50b6b49a3144b7a5c2d5822a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd55edc50221a319a714545078878e4280610a53402d9aa1862df3ed1cbe768f814e89e3096ca23007dec567f37ae2438d24078520acdf419d1f66fcb7072f7ec724f808d251902947a7ec316e6d18d538d5cdd964d03807e18dcf85f9c70a01cdcbc05a3ef962585018b790dc3d62e34900389974bc3babf551c6712d33c06cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h287f165cc8a6bbf5188c5f9ffd0c406bc1a9be17b544fbda2ea20a8a28f4b06d3462567640d4eab695840d48f8678e8226d469f2527ac8972be5d5ee2665dfac400488e567bc344b6e51621896399580356ec9ce684727d9716f1df3cdc92da9f67fa0b16c9dd9923b22d89fcde92fedadef772dfadb85ec18513804d06e4203;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70598c700599f939b8b0dea7ae47d438ebc4c8cd151b258496b5f5ac2ab85fe156f5ca52419037cd33873ca25a9c2d7db963398afe254cf318ca71e988267179eb5b0966b154f3b84bff98c383842374d21572afed9ce45cf7878e71c90c53e887e846a724d6044830fd00e965d94bd1432f284645d7787aca2608dcfe12935a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66bd7c036ec0c909a5d76e03e5209a7df523421e05c8282f2aea0a8ace7b5e4766d5f54ae7eeec0b94f2ae53008e0e664922a0d915c6ab19f3110f79437ca70775e26f48664b7ba228796233a9830f10e4ca9836a52d70d7108d883e7afde28fdba00e21f0025d3a35123606fb1684ba8709e316e6a0779169dd79022e18cda6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h167f1076cdc0ad585bc62a5148ac20253b65d85be7ba05e4e32383c78a7eb720a1e78c889da3b75bd548c134080964e28b2faa4e3afb502fa59406e516b7b42e55dd252ff1c246b8ff55d972c5096d963bec6b7595b821f5d058c6fcb63c332cf2a6e7cf765566e46a9e35bdfdd765c7e28d66d777a1fc501935c05fa6ac57f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha714aff7d880dff19475f96bf0017b8d482e9ff2dd2643f3fade855810d5b1525c6a4cf7613dcab3d6ce76060cd0e3ec944698e708c273db0caafd17bfa7334ad17b7f4762f86aa8735939134dadbbf41ca5c575655c7c3f5204d810e18b2ea64283534008bab2a5fe3ac0450dd02c44ca23df387532e7aaf5b2856cb6f244b6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94940044277f0d2a701cac27def5a07a913ca5c9e0df8342c36ad4f8345adac899221b5a051709fa22c1192b3dee64d75a36e902172837b244b0be532f5c010d6f4a20f31df781f46e45df8cd2f74f6bd8e11ba35f915ebe43889acfb72ce5905965e025d72bfe18396e22bdae2b5a00c61bd9878d6402684c05ba85aadf458b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11faf2f4b9dd69c7ed2648cd55ed0ab2af17612926688d1f2bbc9ef9b2b0b072d1ddfc35875a6783b070a2b80c15881bc3705a0cddf30bea3277ba27e5b234fc5168cde10a3ff12d60e4a50f565840c5ce67700036f455dd140d411c494448e2a2720aa8818468a5ad3a21260f908d6e505dbf83ddd999b791ad4546b8a7688c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62891e129e613a5cb3ace3c6ed282cd8f474b3638a56c05e9a59a9594b3f315ab2e594d99733a54150de5952926df239139d87e84eb6e85d5c4b9d60cffe165b6e50ce95dcf25e007c22604397cec3572c9dde34c099f780a74041193f20125b6fc0f7fd5f0a05c2007e298b829140c977b929ee636985a82c67a00d1de0ca4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h193e2f0ef856493bf400d18194059975eea9cd9d5e0493cbc0eb2bc856eaede8dd893967e6fd514ffc6e3a7015a236557452190f0bcc53e2ff41d8450ba472715a0886e54fbd952d1f069d5c90b470b92fcab1d86f2a776b489bcf54e004c12eb997efd7c5e407e8832b3c23b7041e4a1807e68da6d454feb86161e855f10be7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb610b9e559ab4b8d2e6032babb1dc9f40bf36e4a7e9ddb4a2611c9efcb3e95507427a455a0c6b2a1c8822d04b251aa48e3e8596009dedd82a83f3ead23cb99da92f9e542b70321c39ef35374689bd7c058306b7813b9d69eb9c6209dc2b8c6a7ae9564eaf04a1efa2cbb25674c2c549789369ab937031b35f12d7d3a526c781;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5bd2d8fcb824ba02c5d51295bf3743aaca92b613e8cfe418c5323220cd0e4855e1860be56507e3dc566f896cb117e9e455c8464b8c8d56e5b729de7e3bd34a391e284ae7991f268179a162315cf97c726b5c7da8e9eef68f225cdc4afc91f8f4ceff336b46f31672c40f5b7b7b7617062b4cad9427946ced97445640c4072f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h95a0af51074292d931005ae178ff408d6bfba44cc9ea0744c076168a025cf21ea4dfc6441a55f515599f6e37259df616e4cf71ab70f49a8038790bd7625182ed24a3a6bf36e14270672c369a91c12a2b5e793dd6fc83169e87d341d0cfeb4c67f98e912f02045e60637318989df0dfa6e44cb499562e96a8bb70cfd4e8d0c5c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7ce6bad38f0556f61960a6875a255540d0f62fba12260dd861aff4c8126296c9fcfea0333b92967eb4f0d7c6139c5f935ef8595b7320cbe4d35c85712f3051928fb6a9c461f3f8c920e398b49f3c9d7c9a07bbe40383c4c829e7721750d45537755eedcfd4221524391b1ff97d181d9388aaeac38e5d7ba8af9a4e26a8d77a5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h717894212c9b26d4abecbe1ffc96d841896f3e415b21a6673f552d6eb14af9002de9aa661c668353eeb626921e5a6e098c39e2018db8135321eabc1d1521207f7119761c758e0302de7406c2183a7ffaccfb66301820dcb2e1cae3a96320cef619ef63994d36dcdf4ae58b75a73765a5ee169d66e5048b8a82deb8b2adbd1228;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6580efb27c7924546181dd1bcab051f7f048b8b45da9343630a971f918c5b1105e229658c18eb1fa7d10e082d1d7245006e20574902ec173d78aa48cef49f2c118d213a42dbdc2e67ad4cfe225fbbceb2e594450b1c70be8418c772da584e982ac2ac5890d32e33c8aaaa1c0baa3a32db8e35819c3d1120864a78105678481c4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd5032be3c4b9bbedb567ea4da1caacca3e84acfbbc52fa15db539bdd1db90d64ea148c665dd524060ebb01294ae6127f1f8a84eb85924734bbe1645f8b7d1a3a573484b1565d05dabb993da67b8dc0bed4d19055e820e65901447f88bcb884ce240f3e1baf59f7a2c965cc1d1031d9f28e671887807fe67ab64fe28fccec5cb5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20f2fbc61d0ad00c571e0678d6aff91d5c280b3d357b7516020dce3dc4e372e3fb30eea03f15565e968196e6088f1633853061d2c291f558be62e80d4e9da963e34758b7f086c2d7bfab73de4c9db9d830e3d333eb00784027b4bf4770ea54e18a3239a9b1d463fe0052149046da1906aa11329696a95c4d5fa10ad2b143ca42;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82248b4785ebb0d57e42e6273b8c4527bab63f96462dbf1beba695dc7dd2db89eaf3e7ce13792008f8d63de5fa8e4fcbe052bbd3229bb1d0fb8db2c83a360715dca8cdfd972e27445d6b8dd0c4c3a6ac3054854cd820280d4841c13596b37135818a637bc2f91fcd18d39633975af82ef3500e5c50f9b19e774f29f68ba457db;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81dbd70e290686ea79b30a37f8fd81ade1ef92a86c752837261e6e0c58d2126f9d17e1b3facb3e8b3320f913195ae68db804ef7ecccf7dd451d323d48baf45c9c85097447bc9500c5831a0bf8f3759471910f2d3c831000e4cfd58dd74ff27385bec69615a2b6835b0e00f4e3a49020c4cd9f56868e955708616a952b2c28709;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb71915a69eb153cdf09cee73e1c7b18844a21ca7ce139d98bb1a62e28e73c77ce447121af09d2afad3726898d1d70fa01b39a53078a259365067f839e2c1c982a40d4557fe71972847709a852b4aa6162ee7103473665184c95a7d797fbd1a26892fe7d094e9b676aff449b551d96b3a434bba2e20fff23431e54d12e3f0dcd1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e9084f069d4e059111865168259649ca1111f1655ea5d17e20dea759d586291a3169357fbfb60e20db3edf033c28a79f5373a5f1a051d93630ade5cf20fa7b6afd21259cdafaf07b2040ca1cd288306ea23fadf2d993f1bc41089bd90d07b8aed3d8400ceb1990bd370f36badaafb99e491e656db3b403526a488a67fd084dc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h87fbe95bf95373d0c3fba7668f6f8b03dea3205726a1e0c5fc1a1c2331abdb2ebbfc7a967db714f6df6c26e016016f86adb24e916ad48f7e4049ea9973d509abc311d52f1ed73f58c85de55517d1cfba6ac2d803a7f6c1e4a8951a3a75580e145e6daa393320241fae0a014123227154bbc38cb77f65808d37702c0e66620e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42a577fbc8a7e16d401b47f07be86add9876daf0cbd65fde75c5efe710f8963f2961cfb5cacf5964b4f3d8cd414da3ecc59b527528f937627a49f6dea80ab74f3eea98af999909697df71a453f559cd1e15d6314b946b6b4756ca09a68512d16423d3d1c66f424482c6527e921a781e62f3ad575a7e6b6900164bdc4cdf74d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d6fc53284a04695ae96afd51a8ed604fb029c00d0c78d75c3afa98b89443b8c78d7786945c27bc2baaf5def3b2159f84f55d97f20de1a668eb1718ba8a5b0ae11f994e646097820904bd9058a9486978cd821aa3122d531577783ef69a5fc6e7c3f07a8bfbe6077dfcd1afb262774f16e7f7ccc42c4efc583495bafc39c1d60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha6ac20cf0ac8951dcec1d1c63ea9d6e46f2a0957e68c1f67c415f036bfbe53837dcc71ecde024c181432e8b728d0107d30cf269144d6ff52f3b6bf0ab96ed0b2ad2b558135dffb6bef8209d9fe8673f766457745299e67fd4b79c933dacf755eaabf827cf418e55e65407c18cbf96277dfb9e80e02e8691d562c384bc875e834;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f0398ffa49f697484e37af18e37212754abd788ad289c6062c75a4de423a37e0a70361623fe2d40461a18a3dd7f998606f32cf7eb2cab2d4ee925de7e7c7612f40c00940dde4e201461cb551d62358b592e23f81aab4d770cb3f3f2c5af5e65f41101504e4b9b9e0c5bfd82e284beda2b9bb8c5304f17dde050000e6cab816f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc2b6d63f35e19f378712188de01241d32bdfe93cb65c5847af56b1160119e166f018907ddf1a97ed22441474ba34868b9bf87a576b189429c1eb4bdfa1b075ff45c426e4d7d81192d4c6b7e85cac6040d91aa8e8d29e38998d63a5406918bcd1d12c55898bc7aba4fbb38a77d60ce0daa9e23d8e52be728c36a3be39ad97486b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8dd42bdc615a0cd6b163622009cdaacf92200fdad082b404278050b61ce6d5bd3dba209588f13e50b25995290c32b930fd1d0ca76412bd0e0c89f8b0e6fd69e3950d5382c4f9024db813844451e5c82bd0aa2d195fe4323b1cd3db969cd14a96f953663fe88a554bddc21b9c2bafb1abd6fb156148344d32adb79ab2afd7d9b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h430c74d5414757ca634e0eee8fd5a1fde6bf50ccdd3d0e35492c32f97e0d2a57fbb05c56cc39631e9d77cfffc5bd8a702a355f7c398929bbc90e83d09f44ea9ac96330824a88fc85e3dec271dd10b1a0c928197dda2d5f6afd8fe6e6e391d533c5aeeffc40c7290d532352b8506a175b6275aaa5e9a35416ff299ade064b3452;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae6fe74b47851c3ea0221bbec469facda853369d0238977dc2d9bccbf600605296884580e1fc434c01b66df0eddf41b67bfa08de2c2a64f74c035d019777e2eaf995d0e56b0a73c5633456e66f5808968a47dfadffad6c3b673688bbf09af39507619e934e7c7ca39bb771649634d9ef4f0116ebd68fc0bc72dc84e37b61172a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd8b4967d8f5d8a0af9973da39a57b9835ccc06df71517e620bb919b7267c0013f625a254f9c42fc604d8000fc39db940babd4fbb64135a74aced3563eb484fb02dd23b867ceb1fbb366b9e1a7b46eddde998c9c22da3fdc1a2cf2a10eb60cdd708b7d106e8673d6a4b0bbbd42952fa8f68e9845dbf7adaeb84f2997a0b1a8f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'habfdf4a933d9a4f57ae1ffcc8b84793aadd3e0ee0b8a73f8c881146ea5fa92e3d500c275ad2ff9cf78261c8b03c150e482340ad96cb27b5e1cbe89b6df5e96b6090ddefb70d82e9676d5592c5137acb2154645682f2bd3c178382aa71c0931c84632582c51456cd43c601e1dd70a4c91bf4353dec3df66f8b0cffd31a004990d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2bb02f7281f99d00818fd81c30118ebac303f6e7b4f58a6dd950b7d1f73724294cfffabcf8a995a53f2ed8744e63065dc8a6260f05fa18d0ecd9c0c60a4591f172eba1c54e99ec85e90b2c49304575d66dbc6397400ed65e000cbf8a11552bca5a41b8d53f067038ccabbdc135580962a2d1469e8515e46ca60bfec9d1a01fb0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb66a579a5fcefe6ec3dc32968bd4094ed78f9729940eeaa47b6edcb1e86ab1f0caced4958bbb415a0db418ce587772813adf15347b83db833cc5741ae6be512b211b98113b4171ff0bad9710633ca29a5760f9defd46d52c7f4498ff5a7918989877aa6cda1a18eea2b12e81d37e0a0d58b68f63dfc586f9dd1be11b9c2ac012;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4395edd563913d98ad81bfd3fc267a9bb6d1963d3d45b98de4800ef1b5f7851494643b0ded67861b4572da78367e85331b1a627d8256a5073f7ad11a50c68d34de3186c246bd5eb437ac8b7e762d12d308a140546d56ff6e508414edefe358399e19220bd73a6a64f95118fcf675cde9415b24f14e04a274227f220f19bbdbb2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb7202946b1e848439d26f5249689d223610cf57882d34147fb77ce449b015ef7f0825ad4b7fc1ea34d4d01291ff269e4eff04031b29a4fe263bdedd2881436debdd2924ec29ca46c885ad851bf1cd470b0c234c9c9c7bcda3928bc550ccceeeb9c3536d65919629da68edba602ef8b46dc55a2c34a8a8dd8b4d4a5c25057da1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbb73671705f985f7222a4f5102291e1f98721777bf254d4f7f79571f2096378ba68d5645586ea1342aec0c309b5d9946f4a4686b722ed78f2a9d6efaba787e68a1e362d39fe75e11bda5a927c91f713538be60443a990d8c1f74c18e51eeacd4d7916ddf63b499026b55aed23af8b372cbf29b0a704c5823886d4ef06961883;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea375e209eeb90b66adab54b0939c1196a3f4c226f6b6487e76be15c123437384debd4ee516a926b6178670017214c2ab299e91cea80b1e8e076d5cbb32c94f2e83e78c376a5e6619eacb101907be24be1f59e295a150f62f4179989ca346c900ed414af120a8ec4679f99f8734807e7bd34730dcfe8e61a114fa2bbd9593248;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf05192081e905045a81a0fc8352f1d9753d6483d633ae5bb436eac8959b514a4ccc3c1a892f6407fcd0bc7860150164c79d30f68e09d00bbad926a4c018494f975f61dc159f6a3a226976c8851306a52fa0290db2548d98b6c0e20e2abf5bf11641d1c4fd4a4c312c80dacd2b1baa34ab6b6151701fc3b96fe41070f941e944a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha97122b40a2f3aa7f13ef300d483e616007d1dc78860889dc15ce6919b1c6314ffecf743ecfee9d99db45dc2af88e23bd008548052ff6a97906fd361ea4b942f2150dfef50545d4890327624ead8752043925af0a9bbb945d9b1162b4143bbf7c67e9a110eef2b2d5f9e500ffda16d1f71a52cc9df60aebdc31bf63389900a11;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7da84db7370c8eb5666d72a473945effdd4c1e6e69ea85b088fcd70e9bd25d4d1cd48a0e92dfe7626a52f70eb249d2fcf0e35a135ed5edc97157070e233c5111a2abe9844758a93787b59b5d2c8e66db39a5f419dc0ff09574692012fcb5659d46042d630dd88952266288507de5c81c5eed085ebbc8e0cece5209c8bcbd5ca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd155f2ad9361ac0197766c44080563e69dbbffc309bcf96a40378bddda04ae52a4cf69bf3a53dc91470490271d3ea63f037c483af89b20177083ec4650997bdd914e94baeb707e21d28be390e5834f3e19ebadcbfe9f9cc2486a1253a990fbfacf87803728a958089bda78eff9f6524fdebbe9c1fbb261bd88ea2405b2c0bc4b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79109f59626545b44d811c2d8c7237c8f94394be3ab4b5bee41637b5e341d270cd823122dfa1cf8cf3623ed5583ca62e2349746bd476a6b5e2fe640f5c8fd011319a6f77c866fc2f2992a9afa8d6c0719645841c4c7acd121ff82b5a4489b39730624670af8e3bef9a22cc02668e600b84f2b9994c4d8d70db9e7bf34b979ac1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3520cc98d232992e132d982eff65aa2c91f309ed3d97989dc60cfc17066db141194b5028b37be355b31457e9d4cee32fbe43b164ac1ce055db3d88fed6c633c29585f96764b03b98c52c7b40525024b7e8c8dc0827098cdff3f905af39aa4c726ef4c5ae7b427db5cb5ccb53a236becbae5f9755d1ec6059881fc4c0d9f74878;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4603abbf33f9cd75f528f4c3455cd4ba25cacfcb3200933afa02414f26b588a6593f2466030a1238449263a81104242ca7203a8c60adc3ce215ac804fd7415513de218816ab0c7587700c28cd6cacda77d70b487d89c857126e23613210b0d6c7953d155b5cd0100ac2f8197518fd82445117e13b4f8777e9b0d8a62e3a9baee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h192573beeeda38d014645ecf773545d0d6586c9b1ba763ef5f3a556f0011ea3ba47e24fadf44fd291e168fc1c97aeba75a486e3e93981f38fa4d3d7b0d064276135b64cb8c6ca7a3d43587fe2515ff9bf1793e84832edf78a8f07ddfa0b6a8dbb8cc80dbc0b152c39411ea1860f1f1f9ff809cec1f684090a1518e2bcc30d276;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa05a5935da9d74096585f9df1d2ccad304977d22be8c3781fcc27bcc41e4b76618020cb882b60dc6770bd1608bed409bfe0a671f56aab602c30d7bc903ea60fa9d83ccedfd8cfd74f518046fcac9b116a9083d05ae2fff2bc6c28c4f515299a2e70acce1efb914f6f5bb06e51e181a9689f73b67f3da75c96f0a879163373be;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe7bbac7e308102897a723cf4472a41eeeff46515b2ad1dc809c63000a6b225faa1d503ce211dc2658de956da83be64732bfcae94452ac4951efffb2f9cc437283e33309df66e90508e8247ec4312eab5167619f3328c5d371127dea651bb97280a398fa5161b7471067225f5d8dccb3463e381d50d0c7fcd27f5a000fdada57;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5ba61e46e22c49785ea9340b891bbe4e3f2aa8338da253be490fffbbc980025ade8ea5831b9d601ba86b221270e367235b93c64d03dfc8ee028596cea6412a2cadbb4b0538e98caa1b146db92347f2e36d155606becd716d0760bdb4ab4533c90e86629670014ad6d6caf2a81d55345564ca657ece10d3ffd486f45c27103bda;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7abda170feaf84008c29ed1ef631dce707d99e6778f3e75968c2f96a4e2474cbe9ceebf73367925f3b490a34c97cbc1829c42ae1036a0f115c760820feff0e4557e6ce35518f277b7c9b1eed2a938e73955ade588b003ebb9b1d4dd379a2d5afd01e923663caa70bdd0fe29391f54924303defc214158354ef897ae4676244c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f63f3313dd99f257d731f94f96036d3065b250ab0de8123b6caf9e836c6da6dc3aefeedea6e19dfe26bc14be93af252f7ecdaaf187e8a01f797cdc3e9672d3c5ab2f38fdee2ca679b735398a870068d4f1b3cfca2e35fe4af226cb9a231197b51eb4b4534b6c4694d51b359bb757aa7c9c9f73e7756cb04dcdbce2c9a322d81;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9739de649dfd9f7034553eaf88f344704eba36463be50c2bf3d198695c47b539b60aa2d31c93876298dd2fd5e4c19682e2a7483f4105a9a100354b3cfaee14c32d18c84ed5104e6d1d3cb0c79e977a634c45edbdf783a49e87520669cc8e89ce1ca232c6041ca1d1329d0b292427d8106bf1e6d5bd9ae49f9d67a758a6d5a8b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he5fa9879ae17e79d3d73d8b13ffc467ce63088957b9926ef1a6cf3c38c1a191d94b45a648fee94ea3963d3fdaf284eea2782373af227ccad022a228cdc4b47f512749fa621cc01f083bb4c28fdc677fdff12fe5ca5d2b55408582f8786888175db46043eca534a413b6f167accd0086a5d44186dd0153d08ad1a744a0585fd18;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec8699eb42df155871de4cbc14fb0c2d7e7400ed13b545aacca06225efc3413ae146dccff8add26eeccbfd50e627a338afccc844cdeaa668124310bf6e33f445c2bbce3cc830783d9ed87eb33456cdbabfd2c4b921b5cd4106342b62405d002a2d030013a51c8af8d3ddd711e69c473778bb02df7f28faa20e77d57500205e1e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h904af9ab382161d14fd1cf18ebed4d69cff20a855df121549ed9bcc74618da97d99eea17bcefbf5a31a672f8b2a70ac7201e308e87b95d05e915b5610cbf870ef1d4f76d10cff970ee3a4a7b45587c2d15d7e8de4717ea5bec4e6e33afe1782cde290ada0494dacec757ba510a52fd9957df3ea7a937964ae7eb3ea736654da2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24cafa531150ad14d57b6c97b9c92f1efe491bfc177f871377a8ebc473e42b18c6be2c8d45fa8523947fda1d26fbd67b6dafc4cc2a1a19b94e43ca07348b6027fe7e6ad792dd897de8d11d03f0d48449006c65b93a2e99cf3a7a7afff8a8769992a74f5c00651943977a88b45a70fb71c74853d9e7f8f9bc088af7eae7983948;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heafccc66727c97c79520644e72ba6f9d7832c2ee63d28afa1d616932d6908fd1c131bedce14d69fe1d5641cb853fdd83cc91a8d5f3f152c7bdfcd26f75684481b147f5874a04362a90617b6e9991f00a9a536612d18c37eb33b96229e4edcb52e3f9429712024b1a6d078e12f5285b112261531694124f46c7c76a70037bb622;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e6ebcfaa8cf9bc056e1c5fc75b4a8c67ac715c489c6ef32d244f6e62cd38387f55ca2ea10bb25a156b40a5e55f2c258ee92d0e8be754f6f4ba2d60594cd76be9f3e0ffb65dfc16c66fbf36f1957382ba2da694b0f4f6b00221854e1c4c2e0f514bbfaaf7ca88a7f38c97e9a39ca7f88fb3659aa7633c2ea791de987d603337a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h646ff1b3e804fb4b95e5ccf606cbcae88a1d64bbdb2c77a935b957a15169d49713882d744b9bd9ec7141c018107de6db6a283a71c7d50ad104545cdb7703485cee12c5418d9cbb2c933cff3d1592ed91965c2be2e1ee5fa4fae597c65196474f8eda57c3f60c47f31acf8d5a71991403bcada7f92d72db3ebdc740170db39d90;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h218141b615b6a2bc137e86ac8f3ba1dc56de53601376d6d6dd5de9f02a936756afb8ff8ef42623750a041a56219a43bb21463055c8309e7c5d6f1aba7d20dbf8ce834f2805e3bd33df8e269d19142144d2fbd8324572b56fe80644359a20540d4b17daa2c438d2582391ad1dc8ddf30928f2ee5a21443ada5a3d728e73be0ff6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3d3ab1b31ec620b0fd05c092d521f6e60c828447866bb6a469921b9f87bee09260c4003678f802372b8cc9d3eeddbeb3f67675f3ae79e84f7f665b17e55f1554271d073390b206333f8768e0116b907d390979d95f4587e513672484acf0bdf5894ce31db781ea72976e414b13ab7e88ecbdfd538fe3fed2ec9721ffea43b05;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h468f2cff24a667458416f50e94e51dd2a9b02d6f66da4b7d6b41898075dbbedb9afa69ccbbfb5c12d0894e135d8ac6e5b38ae247ef670430e836836a1ba860167bdc1e62142e916e140e8e9c1cc07e5185ab6e702700b27966b11aaf8ba583663b220adb91140c4dbd29ccd1709f30c045b0248c8b2fe789f9260eeda1a34514;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h99404728286c470a7d1b0f8c7e829311db11bd9a118f631c1d186839e3da2a93fa9046af39ea8eb92640f2dab9def96b0d445a3433e48a2b7773216f77f1c6334af0d10f41b521caad432127596dc7b56f6439cb1918fb44c227a817b14f83029bc02374a4c2660dfc260bfbf7de18e09edb83fd1a2f3fbe27f77c83ce811558;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47ce173e6922a9c865945ce1b6cb06146367b17f94fc8fd66c0868d8dbd85c14957302e398e425ab63168ab9afe2595115a312e2485a6899866f360fb8df9f79703488cabefdf992dbdad35a21b576397a0605c7ed4eeb49ed7003912b6f2eeb4df9fc11fdf327fb11dde6a41921de0ea44c6e6f15b1cf44899e9129a898deb4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20201a3adff03506bb14b0206cf616f6054d435d78de71d1625a36e9a5809db4af3d3b681bb6880b4a40316f701f8e08f1c9a1057f10fd8221545286c7afd6b57a0dc9b331b4b6ff82fff85f5c5ea503513e7a6ebcf3b67751f7cffd0cd54b92780728b5c2326ede24046565bf477d0ef5b52d6fe46927e2a636e0657abb21b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbdfd7c8557f7489952a43849e7b50f6b8d906bdc1f7d45f402bd955311b7a12735beebe2d4ee17bb0af43923af41cc221a5df77e4e9c41d72db39269e138797d246bcaa761c0556b61a88cde093830dd7272cfabcf91502d71398cc26e029271ccf27ca4a3f581ff058fa1e01ca1f10642b491972616e6ff1c24c53291d6667e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7bc4c641d3a74c168187291dbfda17fd0199a51338276c8d0e9c8524df6f52faf895534ee63183e12ccf3d6a428f009031f5018ad9e2ee034bc61c5ce9a6d4ab2738bd89baecd096f83bfd1f1cfe0b34002e5cc98a713950e35e90f3786f5ba077ca61b3cd871ede6afba09371aa8922d17379972d206f2cfb19f5120cc730db;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdcb12859f1ea62e76156857570339c8b3edabb20805fc81c531dec6bd75918adfa6170ae527b956184b823cb439569263941a50402413140ab305bfca15f009aa4aad0c5d259458d3397a41f78e1f14d570b0f4b8546fdafc783339b19b1c83bd7ef62f507d29e62d86e6770ce22eb55bc4cdc5a4bcba3c88584a2fa08b5aa06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8716b47879107c48f075f3d638333a612de01708899684caed48d957380928d595ae517c953023ba312ae87706ebbc2c4dbfb27b17091acf16ada949de571348234294a121bbaa7b7b755fd62947bb37b82781c6adf22daac7868ef4f79fff9d598fc0f59a90b02d4d325831dc3aa9ddb182c763f793ebb0c5a7c19021b7d22;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h92d0808b83962d7e12e7597999625bae43a25df528a0ac33bcd89c5aeca5891ac387ce518f7f8d1871aec176f844d684931db9735ab2b45a3fbea529e155f6a4b89c6495dc85a2e57d53a322915ebe53e6372a735ef9fc9ea0f769cf98cd8519faeedbc89c88803e5ca6b3ad13991c10ad2097505ce27f77364f181d4e92bf70;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h287c6f894a5ffe9e4f78031ee2cc0991008bfad36f09dcb727abbb58d8c65735ca9b29b67d24ceef65ebf08dcb9e224aed3228949f5513ecdf3abe826e12b45b8293cdb6e58ac3655830dbf570a320dc9e90b59ad981801697a145c9cad9d1d4ea056e25f8a6166ebead0237e58dd5bda3e4e071af238ccf94054e7615dec551;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfca016ceffe4bace2cfdc6dc93ac7c90f7240f7341a9a19e4067b99556f85f82a581a240eac8f2dcf428c2f8c60f9875d1b8631e6cd02ebd09ecb59c189e298f218e8dbd1499fabd1db1e3bb9df6a768c4a089a45d215c4a29802743b9ea28106ba34d4f6aaf2c5eae40a5447b927b714e77ab053b81e20346c6bf305c546be4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8a0a79634a0f48ac02c79d4c92cc0d33b91d71f10b3f7b7cc494739bee3d8a1fa6481b0329acd2e78b90e7fdd1d5b2c39a8dd9b21c2194e280a388fc5326c63d46eeaf39d304e0c8056342f8f20a9f99175f78a705df02dcb7283e05c40f68494b241422ba3c6bfb12f34401b715bee190dc88d7f172f06496b69243e4bdb8b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7860f312d78747d747acd155e76285efb80b71624bd5edeb387a7f954ad5cb78997dd1f0ad790282100ed35fdef2f8391fcb9553248e629c4f6c349a8761b1d7b58cba6844caefb8b181c8c65b658b4f28298f9dc63539c153c0fdee81332e58a14a390672b43e74e1f6c114ba5085d1389214a8f7a2537c016592a5eaeb5dfe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b8a481475f27af62dc12526d8d5081c6f79f5578b724b6285897a0a9fad568ad6db6f160ad5fe75eb980b4e14e197bcbc42af66c5ce9c544b06b90d32d1411f12066dfd10060d0f6d664274ce87406706dddfcacdc60ebc0dd5fc7467ace69dedf70a9b57e5e73fdd131741894e6f6893ab287357b5ae9b4965ac6d12e649c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he425ad536ed9f0cc6714e41c978b9cdf9ef4b79a9224e0d6fb3af46ad2bd901241f9bc4b26a06109552c9ed646a15c92ba9b101c2192b71f8663a8bf5b744738c6a4846a0a3b731320d603119618de869c5c5f67d9bc26e6613c0d4c0435027fe560f5df6e499e84ef9cd2528c596f11cd9334192dfb29c94fa9f19a66b82d7a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b1ca9b987278717813ff713e149e2d2e1625ef8c093f1502715f28cfb5b4668cf4cdc3fe776fc0eddbf289d75d086fdfd9639cb5ecf3764cf59a0797b866ab3111cba57c48662b269efe7c44870c6df08b547908c538ec42cc3e8e935d8a9c519ec2646fe47a9aef5b640da538ac57b50d1e7fdb2e056ac2963b398d940d630;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7fc1115b915a0c9df6c1260fbba8ce3f34d940fc1c00423c2606497504823853d904c7fccf6bb78d291506acd5c450221c12f3b371ebfeb944a494ea334e35559e58066356e003a2ee990cda37a8abc3933f8300daad7311eaba62fb0a4ea963c4a483668af2e9b3068e8ce7f41759c1340102a68b36efc1171086591191dd60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h29b7bdf49c0c75effa18f721d7ed042c914d801295ac957b49cda48271cf9e98ca892066dbbc1e2c8bb38d0aa821ceb1e6919cb1645f5035253488ad1c54594c18a9393ccdce4662c706b193c4f4530852c9ed2e7e2e4a4d2759f55bc676522e755e48bdcf3af18b8846050d81404112b21b56fed8dc6b19b70d0c186e279bbc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c46f6b5efac1acac6f016e999e7f370934d4a31fc7b029c9de4671639fb0067d15d6a2753199c3fee3109740014b188601985ae09aa3de5226a88cc28193e04ab37431d161e82c7e4959447cad0bb0227ff45812058f30298bbb6cf9aeedced1974fdfdf09168483283705bd40869566ea6f39d40e522bd328bd89b7a81360;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c21037d43004ee1b63c2e7280aaeaadbdfdaee36812fc73211c5976053496080c4d85ab1d310d5316971e186bbe25a242f1652697a0398c3d099e0ab6cbef89156bb416a378ccaa319aee66089db5b95880d73a09f6fde02b10840cf38e20d472906233eea82e0324c6c4b3fbff0a0fe5e1e471244cce7aa380de4113c49418;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h672c2b91a9b571342983badcbe5441decc530f3f504d2a1248515d36fcd2507918e4f79fd5afbd1646eef42158811bab496166941ebf28d51aff78fac6caf598dc300ea0aadc48038d940b7496be8abb5e0cf577e546c13920d4ba0c2816ae6afada04e511b05731ebb4ee25406e370396fdc422056b471377b762b9cc3e4ca4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf98d00bc39ff0baea27e38e50deaf1178e7b8e3659e3932fadc883acd6790ed3609a39cc58062dcf0f97571e61dea52fbb45b72fd8cea995ce88b910c86081427e5a2ebe801151e68236b86ea993673108b8d844423e5cb5d3eee2b20690081516a9fe5ad345f0c67bdce570c09014f3869dbb6ee3bad14b5baf652f64be2ffe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb53f3b60b36a415d3979b6b6789397a6a8ec8c5bdbb1aa0c490f3eb1b98a7b17e4ad3aaa431ca8ee7b9d5ad99f8a7d631a14c168118b1dd948dbc255391e00ca12471e316d44583489fcb75b5268135cde5d734fb1f8f8e68b4fd1360703f97f64a827961fec5c89661ae52c7f8d83966faa8616e85e54973b80fcbb77138146;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h96280cbc38a19b9f3047210397d1f573796a0674209f8de4a7f4183f15a015f2832ffb65da9d8e7d8eef73a08f0e9250c3e3b996f1f13cec237dc563e29830168d23d1089fc736410fa13e721025de36fab8a1bebcc988f3bb1f3f3778a293b20428255d12d48ef77b1b72d50a031a5778de424ab78586d791983f7554185462;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde9c800612c292194a05a6c4506ae3311868c1384d04b9cdb4565dca03e534a0a963579198df97b0ed89e706c735bc08599661eb09e7d2a7e31d2a5c7760587d122506afbc82f71a2782d458e18b4d5ebc73ce0c00fda33d6ca97badf507c19b62eb9ac8d0bbed3f5930963a452e8b0c1f0b7492f52e89494f95cffb3c514456;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32bcbf893421d38902ceddabac9d463ca2fa397e226894364d68538e8ba50c439598bd3d9724157ad052588c361e3804536038c1cf4109289d8f6dbaf7a11e9ab35c76e57ab7f17c2c1cac92f9fdc5da00b7b90181ec691a7671874564d80d780b9a4fa728fa9261890eb1b205c2bbf229b583d7d6a259dda25bfcb6162640b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba80480476d5ff358f5efb09806684c86597721df82a92f5aedf4d8edbd3efbb5bb2194b43cfd1c51aaa2b392edfc3f90d64fa46443a06f931a08e3d6f6b70b540a4a9056868b9c0d6d931420e3684778a4b596231069a7a91ecd9d1c1870e7fc032ab7f5f4fb9548b029f5f6024744e0cba8ce696e8c85dfa1b1411135b37ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h393257b5e91525d811743df2083c48bec741f0891cb3590dc3533692e7a2a86386f59c8dc345118be9af9b7da2573976cc9feb1975e446302dbcbc28c36867df0cb93b5d4196593cf2a9b997950105642a789e7feafb14d240d4360e1297ac8bfa3a95c86ad8b98fd025b709693c6920b24b2f707232a1210ca959d275dcad8e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfdb29dbec0c35aed3dd56bc94ea19445a9e9b4b1262524a7f02a3dd60add09ba4d105d95823390f49b02088614658e1098c6f5a00bb0832b0975c41c943021ee8f322664d88440937494f126e9606de99a31249c5e8be57362f9be31812eb20a2c305ebebe5ecd9727a13d133eec154ad8e2b8fd82fda0d97c4c588104e78a7a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5de9260f42f5cc9deccf9a36fe3418019da6afcb2c76be5a643caef4b69b9a24d28e81b1b3bd897c7b64bda6c4b99dc9e7fe9772af8dee723c18801619a0ef098acb41657cd557e989bcf9b193b02cb9a9f3cfff07b34caba4761fc33ea32cad07a3192a342c367a886ee8cf4f5a9a15737b08bd73c822ebeb3831b5046c058b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h691e5d8944d16195e43c935d2bbd7e1c8b425a3e5a372d2cd193695a9af59a80b15f7dc8d6b56a2200c5c105f395f62fee2018c837aff1789589b4660f8921f9bc10c389324b50a1b0304ad94bd741820c0d1a58d5535c98a2d35557dcfca60376d881e5484b2925bf5a128dabb4adcb63385b4a8fbc9acb95de9a74ae08aef8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2c6a05fc6ccb072c22c7e33c87dfd85df6be296e28d257d99e473f8833a03629228243816efdee5865b8ab310028dbe4c669c486c87df0d74919cfde4854a617fd5f6d20d0c97d0e3f82e4ea183ffcd7c346abc01272e09bdd415ad6a253f5bed3baf32d57389c16e50c8e0b2e79a2e025b677a59f68544da6654b78d1dcacc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb764b5e71a0c7b371efc76f570192c7bf05b5db4818996ba8d18abb4f231c36e1a931a4119f8767d1380f04ddf9fb0005e082c6f692affe0720e8a5f8b9f9cd25e1c79f06e3f3fc6cb9ccfb19100eea3a19a067b9388d73ffd0b92c00c00142239c83e47670db3bbf30f8d3d34e90aa778c8078c85212b2a173f46dc9be208;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1628e06fcd4b76faf08352df8c807be4daf318e3083465df463a236bde11ba18b755427d3eff5fa94756a00e7752033b4857697288ce3faec04ba05e1b7d6619f4b0651f3bb2490dff235612ebe5c15c090db600af5ffb578f3c73e1ee8f871a7e9adb882322983585b914b01e6e991d6a5259bebdf894e28939d4b653eec6f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2580d10cfefb81ba43a926651f4a6fb3057cc5bd57e20f9c4991a75eb616d0eac5e5a3cb0adf47e768355eef47273037792a751097e206b9864a30ac4f55851ae8f3681c50070da6905017929557cf3f88affe0afa09c49cc1f3132b9f189fbca86357d0ad3106f8459cbbd0c466ba7f701b21bc57ae80b11ea0145d83850cf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2f3795ad41cc65549606aa63ba6271a37081121e93bdc010b5e2b68a45a0475b95fce0332232a30fe4daaaec33cceb1464824bf49196df6eb9b7be3e8581b96decfc2f8a1224940576838819c318a9d777221b2b84622364b740f3e3bc3bd521d9ff4e4ad475a51590cda74308d8dc8e685795b9d1157c6e3b7125e1947badb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e9a57cb12335e7b2852d42a076bc78a51882979bf646ff46f22a791d9530135f0ed220b628565577a95ea222ef704d40e214615987f8e41c8eb0d36b63001fa432fb6a1651236f084d14391c5006b0a4fc50c6c2dd85b270d6704aa6ae0caefd81ee8397e1ab10fbc361ff20d6cd494688e6c8161da4f360cf457c8cf295091;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0b37ef44d5beda265a7c33172c00fa0d04b4378bcf4c0a62fb71a796cfdfff0f259757b98f98bf6a8b81c6e3c1996b8dd0c93a8b8f13c8a0f4dafac43438bfc9cbe3007143d3f346882b6a627005c6f85910487b23f90b5016f5b6052ab1788047ca1c36611adf8d5b4ae8ffa1c6f4cbef0048afca4e8e3f4b6a5ab187e646;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20b1dc4bf29d92b7dc6bc98e81a7d69010625de3cc869cfd4bfd05bd87fb498bb8924a4fc83c6365f4cedc4b3e94a32c67c7df9569d798cf793a6712b801c38378d1bb6aab2b97a4ff92e72c4fae4962754b6f73a7ed9a4e5345d9c05db969fd61195927c88b252b4858fe597ebd32e4615b6ea580e4c9e40c94a044ec08ef4d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0e2496496098e3cf817598a36789ffa0c913b678844f18e43a124a81f31523402525a01731a5fd35ce7725926d4e166889b7a62da5d962b50d417215c9657e164d53fa72344c3c1470e2707d4cd705b7b00e809688017df9deea07337d3fbe3c3f16d5e8e6acd40d7dad69b8a3bd1ec4f14cd1668052fcd45ef9fb7a2717c13;
        #1
        $finish();
    end
endmodule
