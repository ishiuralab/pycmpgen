module testbench();
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    reg [31:0] src16;
    reg [31:0] src17;
    reg [31:0] src18;
    reg [31:0] src19;
    reg [31:0] src20;
    reg [31:0] src21;
    reg [31:0] src22;
    reg [31:0] src23;
    reg [31:0] src24;
    reg [31:0] src25;
    reg [31:0] src26;
    reg [31:0] src27;
    reg [31:0] src28;
    reg [31:0] src29;
    reg [31:0] src30;
    reg [31:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [36:0] srcsum;
    wire [36:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1eb9ffb2d3f44bcbdaec0730528473efd575bcafb92cf026b35e25f4b5b0a969296d366d2b05956f606c2dff28f336a83afa4bd7e93d61ad51f799df375bbc7a87af89b7e40e4c24223c4041a7768cfdb3a5f3941fb50578a5c035a7ed532419a264ac9b339fd2195999c31df354c13fc4a3d7a0caa3a9c001f6a03c4428360;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18c3a1868a9a4415f19fcc35b1d845a1b29f58e0963fecc5ab9160c3b6d46e5813929c4c3c3df00f02b1ae5a2327df114f9ac74fdea1da25799200aec4e871d89100007a82ead8950efb771647748c25fe484de890483f45d57bfa316595e281bd34b1867ab05c889779a5291776aaf7bcc0f140c59e399c735b753e2723a3b8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfaf1eadb2ac75d0cb7122223b5b3927c144404a14c9e3aec4bd358822d18dede4388caf1ca34989318610257cf9ec696750031fdbe5357b12a72db696a45427b5c1835c1e91ce4c6e3fcb4624aaee63890aaed4a5208d1314d49cef1850d64c407c5a63724c5bd8dc3b9b1dcd08a47cbe6c4945226e4bf6b565eb8adbf8531a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h154f20b89923c3f597a7f68ff36b1c30d5b8319fbb2e7abc9a4d0ce3ea67e095d1f55e78b0ad4fce8dadf77aaa8e1d0ec8ed7b29f73e233478acbdf18382d3dba4a8471526da92074c07d53ac707f76135204fb763bf15d97f1562e18af9b29d2463156775b62f50dd57f1e907b9a7723562836fb61afaceee7e767bb5f1e82f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15c1fa3be08ea1622599384c96b75311ff634e195ca4a5ade7829aae13040be0ee4ef21641d90a710c4ca1f07c15e5221290ff9d3810eb1e4a3c51826264b352578f8d06daa491b74a5ff544ddf72a7451e48837449f8d3e324fddbf33f5452e97c888dc660729466bfcfb92dfa84a3271e8bf791ab967c3517c96999023111;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb92b9d251705aa9ded9c855b1201162e147784cb8007b0208c33cc851ef851515bca722ff702ca4440e01ecf3d18ecd32e8662ae577b192f5da15b2394be5cec36ee0a4db672452589619e39e939dd9521d1b8eb514c67adbe7f2d41333bc070f4af8a57bd4bc750b2a1323ae86cce0259c7e67e10fbf7de27c48a103a65e230;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h466294ea2fe564b077191f05423f80e1c3e9b377656dddf65b43d76ca4854a684cf64558254bad4a1d49d27866a2a504d5572dafd9702fad069fb2adec492bf4ff4bcaa850cc85bd91e9ca68ac3558f6e0ec8e3936320586d2d97cd0a28ef01fda564d4abaae924fd7281a02ee097f001b5d83a9a19c36a2c1d04319dff2858b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h224d5140e7a3482c89627889a52df1a9163b7e39b850552f92af8999508558fd969ed35063106496b09293ae618424d9ed3a53344bbd75882281de241590eb91f8b2af2a3fbfce19533a471db2f0f48041463b20f8e593969c1d8883459b931515f7a7c6a14e0ab072694188f283756620f13d7c1ef649af4e55a5ef571ce0d8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c769511b955ff1bad798f040f0e88884583e815e3dc0424f50cb517b30ea7562b085ec00279b8d584bf7d81aa6521c1f01014768be011b6604f1001701504aad2644300e6798cad898cd17fcd8aee8dcc5c51b119711177a3d952ad81b92e4b61f0b8563d0406f5190675735bae8fdd10a0b290923c5209e993952ea9e77b25;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2dcb78e109fd1a956ad61a08fb976c13db059d97031e87a46532d9335660556470e2b0c79e013d2c8befabc9f338cbda85ee0b71f8db083b8c260884983cdb55a87f2643431b4451497d1bcfba4d952d3d34931fbc52cca835a7fa4251eb607e72b1e5d0cb7fd3ab331550cac91d245e71902f3c5e1808d3e4ead81819d985f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b51886fc7cfd359307f70c758a74fa343499c290af52700de721717d72b784f4065657a8d46bceb3a946bd8b0bbbfdc89013bebdbc4737cd3c3367b5e2f8b392adcd8f5df07db0564272069b71436619a04966f08679f7c8891f4178e1386e4aa9f0e3853b7beeec17f19820f73c45e87c778b738ad4a13722df2fedb7d5495;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1fb3ad5da07a8712b081066167ea0051e2d6039ca05c78c7d822d862efa4caac31f0d15bab178f0459c85b1d7b41d06651ad265a79f0d0adcd460c806122ee41310276aea0ac531560a494c6d6553d823e8fe44425cd18630d347f0b5a0682cfe00b7ef47fdebadfea1039dc3047505fa511d87791e7b08f284e2d295e504c03;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc012296b3d52ba03783ef13161cdab911f319c6a08d6304af09349b759568e9d3f8a9d06c14bab82c72151b41c0caa62fad1a9ca53fa4314d224ab556d4bf8a001f5f851246dcba0154df8a318c1f31991d54f2268364104560c6705c73461d97018598c7eee2046178566b6c58b77c82101a9e976c22d5b25d97541b3d75f41;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h795f7dcd601446eb88893dbabfcb878325b90db091996f1f8f770a386ed14298053eb773db8bb768da748a70260f6b27fadd25d0d9d268688a1faa4d7292e1240b280cf983ada5acd4ab4ca5f9c891ba290c3f66ce18e70a674b4a86607e91c48c40006a870e5dcfc5668c426fe8dcd89eab44380815228449097e1b4ffa83de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6d99e2db67999a5d02986f4952b23a00e2d209498404c003b4f587cf63dfb4fffee4c9ce2c7cbc5768952053531c397aef8fed19b4769da45399e714930abc7eb29a757dbc85df0992119d7a6de201c825eec6cfb4650bb8e6e22c9e0f59e7d429b5fc3a45d165a3ccdd881b89e6746d008a650ba5299b8f281f80328e7b6759;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h947f2e5090d2d2b84743f40db843ab6d510eb7d066155b19ed3408f606f9ae57bb9d3da817431607f6e75177661675ff4362a048ff48147131ef95dbfe74613a8e2800c5fc46999e7010fb1e449d442a7c39be6ff4281c00e36dc4faaf55f56bd6ec1afdb4cf2aabfe61244fb48555b3f67dc786177a65ef76e4a4228ade4b08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd60f989daff4a3c95f2bd4362a45a8410ca0221d8563cdc8e1c7c8a1d801c77abc9af6cb21bdc4b6bbbe645efd64f3b25e4da96782c6d69e84c416e37e2f20fbef158cb4f1c82d924b166d4e9f9199809e6e08a568ed680d93dd12b4255fba50238576685b164376f024b9d5030a4c9466132a4b43ff3e5edab9663e1dd5dda;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a88e67a67b8443879a00fbb406c38c9fd42aa846789f36fdc0229bd942910dbf383271be9adbced80c03100390213136edddad8dbe4c3ebba426c0d7307063f7e3e5b6f037400f49b20bad004197550685229fd9ae536a4b716498f91991b7ca7416fe3c37c05043847b62effcffe879c6a4e28c15216802460b0f6b3107829;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h28849b6da7ceb132e10fb6824d0b0e33581dbeeda87b665d2965846010357dcbd9db67670da1764e135ba0edb20c6102eec49fff6a1d9848cd37f8fc09c51783e11746969e442935a1b839a18ecf6fc06bee67bc0f92afe451299e4c8da6699c3a8db54e6b541f954374fe3af0b6f4a8549c5e72ccc2284ed8c0eccfa013b8ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he715fe2aa0b84ebfd947195f2006fa779def6032dc96adc73e04f9b8903e941704602371119d4c52e1028f98116e7e71fe49065c3c9a255d7753f6cdc8228fde84bb4c4e3766bb14d10e2d6aed8a351b61b191e6b3063c17ceebe82e7614aaf6877e986d09c8c02d8a508211aa9a5a4a03e3a2625a7278de0d3e6d8183228c08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha485c9cfef7c22de5227cb4b0c26fd694464d57c042e566496b02a2b30a3780dde76cf6821698ce6db3437621df0c1f05916a5045aebed1e36e6c4c378c4ac6f31de38198e69093fb973992570cedc327acf5b9e9a976851920c3ca36db6b454e12e900e93db316fa2b1848cd417180bb18f8dfb7957cce32f1c34f878991622;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea1f4754378b1a55bf02786d59e7e3078444bc0c49509c13bc5d04b61c145e61ea7b32e9e37168f7ad191f83ee519ef91ad785bee9a2cdeeed6b155fe0746a0e7191d83bcdf3c29b8f32a3d5d863ade7b97554798dda8884303e973e0d2d3bba6ee51f8490e791f8bb7f5e33ee4c2ac13ef2ffe31684cf3c99709d1763466ff3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha69e5559fd8b46f9ec569e5d5bffc7be6540c39c7204d81d3150a25aeae778b2f80a9bc51ec8bc5d8f2a8b0453c04780c16c81cf3d5106e3df5e7f4baa863b37ccece081642002d59e0b185f38819cb87c9ac13e648b8e757a78a5d6830295dbb8106bfe7199e9b80d800a3d002256ac2eb7efa4fd84c46950e7a6ff804db23d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4a44d90f30759ff76b122f3f4b8b387313d64556801b55a7636e7498a21b050fef7b82c0cd275564c4283777a62819e71fd7e6b7ca3cf209dec6622c79a2b88af29fb1aff4034e71d4aaa3d5324e01a75c9a551b08a5c83c7ae2f1728cda26602e5febc458ba4956793e5289da90b983e9ae7378d3b02b8cd3209cd4c51103d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h207d4aa9db968bb6f35ba18b7ec65876ee72e741a468e72f2d8a04468c8aecf5fe8506ecd9812f748be4a3b151718960f8af0e92b2035b9b0ffd459ce2cfde5082f31e279a8cdc9c954d51824062bb11bd31ebf258e89bcdd99e1f61439ba5b72811bd3130e54cce6d2a0e52e33da2b4a9f947cd61a1ca325bf2537c36465edc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13b5d2284f44b09799d62848de7e34b96ba892b8cc3ceeb9e5ec7aa4d5e5c8684f1eb84ba30fe04c32039268315ea0ac149a5733861f91b32c3f7c0ed37638f2e361c80e6ba4e32b17ae0450627fddf96c9bddee7700a8f099cd1597cf2296cd381b819c4df3a1927705ecb58ba9f50d8d9106a109f2953b8a119a5b43900cf1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf51ddc22d8d64d62a2ff547651f6cd2fbcadf1b40c06c41b0ecf126d823b2cd039f9f37b978df45bc75dd11f41783a1e0cbb01a68254725c8eb2a8be32ca5425d15860bc761f7501b4e8f01186a8120735d918b761cb0ea02c75ff3ca80450ea172a6322c0b37b6327d7180f0a1e0e0428bbc9693692fb5e1d13c63efa33210a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8ce47c388323d9faff6161f6469b68ec3aa38deb70252e32d9f91050384c9533bab5b38c94aea5e7f07177d16befe1b7d1ba544399cd60339a0e35916dacd82fa280602203cb065ea717db49f0a411f1ccd7aa8004d08f351a4b29889ba116e1d0771c718e6d15032f15b0019a39b551a05f7cf04bcd1a0a8e1dcfa0b34557e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdcf7adb4146bc284a02e2697a87c524dcfa260009edda954d815dcc2700c03d32df762433f275f66d96b966f39e05743634e3e93dd6cabe11264ec581e653d61e4ec85365fc8c4064d983bec483a7845f799c894b154862980720896a166b4f6985a8c888ba3f411793d73eb70585f55cd31a6cb9c69fc96a0107a8939f1c325;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc76ad2dde775b5f9bcd86e0e3d899f1ba85f0ce88710dacd546cad0ecc2811551caf78c5498d70a561173b74f5f889a61997308e0ff6ef8be3b5af819898db4c5b6b8d20849545c18d89d741c72a4fe621f930ce5427389f98e77a499b7c61604bba9b54e51eeac04ca1d2e49ab44d7fb71706ccb47197b1e7350358211e671e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13f6baccb24d9df603dbdd5fcd4e7fdc1bef530be3745282c87370e478242b1d2c43745e859aa3986fd7231fbb55874509e7b79d8785ed6a99eba743948280e442a8dbe468e2a8b2f6406273d7051a7290ea1e99421345e9f12db70690a1c9f9baff7636deb7e12c7d2f5a2b3516bb1a7bd034373fc19fdf9b3c2944d6a16317;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1775fdcb822c011c19f0871bffeffc57547f634c06f882dad0770c0b36fd914a9115b5fbf5ab2410619ab4702c8ef1b4a6354736f18aee6b5290883f9489e5e5ed072e90cd7c108918bdd69176769a1e100e2a2d2e83ba27f142efa6d3e7576317679f4d8876a7fc5609f3a1bcc6963d464e954adbe7542bdf68d73287348784;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e8e8d3ca491dbf8342e8b863ffa5c9254c4a75280d94351a8ec96cc6a5f0176064cfb0cc0030f6b68bb92a4220ca3353c3697e647f7278a7988ea04d3a41b42247925418163975777edfb1519d753e88591cdc2e473f4f2fdf3ec480de2b41fc85dee19034aa1f9bd4a9f9f659eb62e90464bae9be545471643932d33a4b409;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h77be10dceeda1d1a0b57845bb8f7a2872ed814982ff9676239b83bdb9e4e137c0c016d3026923d92ca5e8e988fdb304e0be2f347e4156b68c687107581d49b1935c69d527f9589e9dc7ed9a11b76406c855f314c2c882dd19b52fee757ef664830891a8952f8b069402d8c07e5bfd788f7a8ae6e6791ab3b571f63d48ff82f69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1ae9fd993676693c9d07de27c3240055b780b746a36c9ef1a15384611f660e2adad1522d2bc0b3f33a0b50846f46467b87eb86a58048358c95ab79acc6c258ad5faa99f01482279040ac71e177a3aa097c3988756c2ef9e65eb955d3b6c1d51713aa71d9d2345d0178e6363f3cf21f42682f7007938ffb58a4b70fae4ee59e5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd10a51745297f669c0c641b1bedfaed2b98fb0954874d26cce30ce03899ac56e6c105e323ce9c5f258a9b9327dd5bfbfa2ff72318d0cd589153e174df1ff4725ae6c012ed1f99f95b631b771c217f82f2d51a0c567d0ea0dc244b32333e3989bdc90bf6e5974b9026bc2a1db7827b7d83a65aca090a5872352fd10203eec1709;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d78525be347090b0b5050584965b2c01b718089ee62e4447a5300e44235a869e77bc3efbe20150090a95288eda84ed7455d817fa0cb2644d0160bbf57d72045f4ff46e16941776051298f5c9519107834480a245fcc1032a1ea8bcb12031b0202a82f8904b20efcc743eddbda3c0658889aeaa3cba53dbf66d58d7f17af1de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heab21c4fac4967f9c7d19f6b7fe09a0847684e5f43f5806aa20dd15e3635a65f200b70a6fe83fef29cf8f15f57b521f9a6d88896ed03531b5fa8edb30f2d120d1bbc4810d4c3313f8aa4a5c2e4c04e88e4a4d3f03a8a36ba45d4f5e7766dc3a4fbc884d9b070a188b2558e300e34fd24526bb04e3beb2196e173d743b3297faa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h492d92e10056760e78bab7deb2a1891c96c7b90c6aecad7c724f546031a105dbd474240289be2fe5bec44bb55ee3238a6c582e365065dba55f1c3e1ddfda3afe060435dbdafe5c7896afa86d35e28781e14bcc4f563ada0e80bdaa44e273267e160a65cdca58586c8420b6c120fc4911ed2b8e038c5843b0a6319c3f1defb32c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he27dcce5990e19d658c41922c2d756fc895de348d7ee73c13c2b64248e65fc6f3aa5773d7ac3df3e139466b91ba698d7860ec2afbf39f713ef85484ee58ba662491b56b88a22089423b418a5195ac351e3bbadf5eddc93e3eaad69edcb98ab72cec74c11779187a68cc5f0d947202e43417f752aac1617ad69c78bdea8dee2de;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88ee2d18919a29f2f7e2006febb24d1d856ae550e84b8ac0274fac28f752a71ffdb7ff3264bb8015bb6ae614d63a32339f247d45e4ff49c17c60951a87d1e0a0a30d02116dafd66533cb6b4f815bed32ccabe394a1a7daff8a82390baa2c806936a1defdf203f0a4d29a94e7551726c5cff5043a4f0b4400dbfaabfb81a7ce57;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h354f24b61b7fafc3b51e9d7207a049c4eda2297168eb38b244e49b23cd7053b15dcfb3b11ac436d44eb86e56dbf59ea80dd97935caaaf702bb1df8c160b1aebfad3e0be029866915fc233d0b221b5e3cb7d6dfc7281f7fffb7119164c61ebff67dfba49400383c1f99abb467f6042a2a705ab8999320e9add5bf43441a12b9d9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf9fc18f6bccd05c0ad6d17e8a8d753a77f7481fee7d23c375dbefabb61e541a46c7a9c16e2a2389558d22a807d3416451f2c100e234fdec691d7eca739ff759dc6bd32d5afa5b60bc1ec7377504a8fa4c60815ad77c9fde828db95e87bca21a477c824242df4ac501a7dc0496304a10545ebed4f243f01af1367cd7e4fb3179d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74858c0f5448070a4cf806a1c031e374503402e4d1f6581b0d42b46aabae7b39b965a87d3f0e086b6c61ab643eecc53f8561a7442fecab76f4e13c0d7e6fc68c15779d5e896ecccdccf16125c8f18268a9779ddd448b298223c06e5ca8aa63f001c9bed807fd8b75202e284138f4307b6340fbed62aeafb9dd5a0149972786e3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52a412b7912a5caaacd622aa44b671cd94e6129abb7a9760f06262d40a856e2b54d7ad7e59771606f9c61e2bb98b760ca415b08aa986e244bffa11cc268b114245508bf99cd5bda3ceb592e844080b0614c8bc88220e6b6b513cd94e4ab3bb1a0a70dc955ed5abe6ea9185e7dbd0ed2bbfe10d2d7e24d96cc578bb6076ba0b67;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97ae18cebbc2eae01ce3e078a6b9705dfa6a7181120103e60a956ce625c77f5e802e44cdcf824641c326c07ad6f1b6a19d17b609795c1fd0789f963e9b9d038cf8e723d606e18d3320d6318e3b76df6456c46aeb47ccafcb2f51056693cbcc49c600c4411c485e40df3b533d6bf5d6dfafd3c10e0c8839a74228ddde013ada13;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hecb451529500ba52787164ab4fe6027e0e8a1d9528601cef2ef996de6ed68d48e23d87ebcfbab37bc87ba3b1bcf52ba0417f23f21dfc32046bd86b602ff587c69a447780b40931a273390a6708c98286d37a519018cb7f8d4dcba22cf5e76b187b8599cee7d2ad899f3c31b0758144d89f83a428b6298c33ef7aeaaa4a0de10d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd87a52f99b4f7f70a34eb2c7104c936c16e9ec58f58657cdfc0bce129d6008aff0f79f13b398b3d4357f5fd6a305562146a8044388217d7d69b98d76d013a6df6b2f467e39ea8d2d7e6987ccfe21f557a86c40c5f33d86c05aac49b69fdf53bf7ef0f345e969eafe3bcbe1dfdeefc279b80a057bbda22c6384bd7be769b207;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c85fd8f32c83fe589000c89f8c344aad33cae50da169a28e55ffe4793d5c97582b358c70fde775385c4eaac06e2f103a6cb3ac47eb3ac2da835c9019c3b7280d0ba7febcba312880d134b1dbe1fdaba6d416ca572de51e61944ba7445bdf6e722a40b4cedd7ce90da6606fce86c645758c80804c2454c98cc921e358c63bf03;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h76965d97438975189983db393f6866d334041b8bfee860b320714c30446c66dfe669e7caae14dcc88cebfa98b0412eb77247f260bb9e933c566d4de38198b2f6efd38d15ceedc937cb4414ed77b97eab82a40599519b886619a18f7a353b3e40c85435a2230d14415174f3855dea64d30edd89ec9d1bb053d20d55ff86f27404;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34f66ec606126a09a5dd9f82ee9ba4e592bfd961e865958468b5809ad2e1eee456907be689e1dd28a15b87997bf3ba31d42c6eb973819fa487a4cef12537c768d6fa082270721f44ac64ea36fa9394f9ef860e85584540a022d83143b25d74f665137a100815531cb9c88ce45f7ed829a5e2d23e8afe60c2546b975c13928670;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha78dfa3d286665e1d22e79b426dfb52842892fbec6d8936f60a596f313978620dee6552365db049f944ba38f9cc336cfaf8cb16913ad513d86b6a88cc3b8f4761bf24d2244f97d2260c211bf742f970cdacc64e1eafd7665494d2e82906983b387c1f6d5b8e270dc1fd64d80ec0ca7f3041472dc66d5d6186995170fe70e249a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0d34d0397770d0ed20f2973f643c18631a940d2a0efc99624df495fec0a04c26a9bbfb31c9f53b4258f44200440390852003b21e9fa70f96a707077d638c1f1b4813edb203aa14ed7ec2cffa642593dc1596f670c792057ccc423d1cc19e4a78763d40c854199c76fef7b31e7a1f26d9d0924966c80e06a2106c860164a2ccb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8b8e3b8367076ec075b4f394b1e53727ecdd69172f12a8499e930d3f4784930af8779dfa95af738778558b2fa723beb5c6137ea99e0bcb1c061042da7f4c193f7b7b18965f1aa710068e7911ae8176542b6da157cbc8a0770a7a7fee6c9f440c5d3222a251fbe8bb780223060b3c74c4257857dca0d1e21b9de35e04d76b52;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd9f5e791aadaf5ad380104fc8c59b6c5393a714282725afd7a38077a993ce4c9425d2a9026892d4da732d2f2c36836a4b428584eb734dc3f165604f461a8deb7d0bc52519d2337de8ed17020b6f5b17bea042bae3283a4a3a646cce056b929e6f325e94b8ddf0ee4474d9f7068de04361709c7bd4c009b92f6c2021b60b3a4e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc83b65895ddadc9b4b71f50508a50b204271ea7ec7785aeef8a945463c1291eef662a132aa9ad1ac248cff58f2486f19fe76e16228c301838e04171ba4d90f08373fe7feaa6cf4ac7631edf602cd70feaa6173287173ef0e2eac468c19e3ab27d8c60c4cf8d805e06c37741a34df71a349850ef8d8d03c95b760efb2ed43d0a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38b874783a0a0bc8f70f1aaa1ca5b7a9d770db2f1a42e9b27305e63394878caf8b0a1ec4de76474a73a0c9f2c386237b0055dca116f51691d7493832f8d20bd2a8536f1dcddd462c443087e5af8d9748b7b8deda53a7e6579cbf1595ba1bfc170aa6adfccb4c6921ae5f7e1260c2c04e6c39988dcd0ce0bbcc7fd99f9a3831c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcdfba925cae666c26883f29ef4af9c4cee9ebe019616dc7263322cb9ae3477dc2176fe14b7e5f96861c00faafc363738235a2e0e4dcdc7af7e1b3f8dcd6f494b45472a811734421c13874ee9226c4d8997551ddb1f619eb87ab217c0d3df5cb0e4d0f7f12359249b989d19fc9d1710ea297944758e0d8781c624fec21ee5fa93;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11ce0fcf59ff451092ca2e0543c3f5496f142a71c2f0a4a0387cbabf3ba8564fb313692d3dba314b697a72efe4025eecfeb569dc7733294506d489146968e5fdc666522fb44983a39d391ad2417370504c76056e5368b6de15e8dedd2e76af134db0f1c8051806aef6aaae2f2824e3316d5b527e0d798b7e2630140ed4d17c41;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82676793747fdb5b46de40a7e51b61df6fba81baf2f5d1b78356583d2e0bad8a51ccc9fd53a3f6878b399053f617ca1c832f676dda1cf6be1048d754ba15704e156bb2888ee8feb9d2a4524cbd346b102aef07d599200affe7f855495e3f4319d11201d476ffad18cdf8283ec034823b4aec01310fa0afadd99d303d2049595f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8683b5fea8733274f512c532386163332dd9d10b1ecd63fb2a5f9eedc7b0f95dd8a737352c326ddef8b8f78585233e8f1f94f9911c41fe47647be8ceb44d41c3a94623e8aae28b4978d183b6219c22ff044a7df787161f560184a0eb3fbd88918010893f385b998158865c725ff3a1b8b5ca2d5bd7790ccd5cb92dbd3cf8c159;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcfd13127b88a2304f85815b7f53098ef05d6b2bd4cdae1963fb616299d7c7d870780bf33d9c530e320fea94d1ee7a732739eabe6d874a3909b1cc85166e5683af0c52b1962dabc9d80af4e4fed500aa13d3bc27fc9631c0c69622e93ba8daec15e3c424e12e1d4ed25a3937543c5f5464da415678b893c8f6213ffca83c306fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18d7cc9d36b4ece7c59058c2988e920c32095f77799d8f96f16dbe1338a56618c0daee1c9ee3b7129d6e93d97f0fd2aff6f474d07e7b0219e81df8509ce9539149262ed236dbb4d5f10d945aa9c39c984b0aaf5094c110e44e48022e8d69484e76ec0b35cf7b7b2e74d73b4e925804d3d81dba59128b57cbe939611fce30e6f1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2fcb0b9b6844416b1be80f5f9d4e5f5118cead0899a106f08a280efe2eebb2d79a84ccf8539e9dfe0738609ab9b36d9cd002f53c26f37e1b56fd80a936d3883cf2a2b18c3ba9553c5c47e079963305fc209983d4c30497fab0f85b117e1ecb16e105aa1ce19bdcf6ff12626ae0409cbadb5aa338aca1a929269598620a9c2edf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed932564497bc1be4db410f50487faebae560f00fd456f860ef1338ad8f2e738a414ea7ce23a347d69a29ca39205844d1a05fecb3f0784bd6a217ae3060fdcfb900d58e184006ac2e3f97de30f53052195abe6b155abcb85b5506ca5abdb13aca7a243999058fe4b33153ce5d4a10da8963906e3d1911f1da2443b305f14afcb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h29abe47363ea001d1737fbd9af8ba599c06124d0d0505a9d4e2a92258764fe9ff69bd5ddd380bf8850143411e92258294725fc3f7fd5080b508a4c1dd1f75ccbd05b0162795bef59b0e30f4fd8c7f36695d8e88452bbfc84915cf8cb98e8183f2cc8be828197acb2da028ac2432f7536dc6071cc1064fb946a3a8e606d20bea7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a4aeff1c21f36edf3b9c9703eb78a09aaadd77eecf688cad97453b15aae88bab5e6c62cb03d77a4325aff6fd2c4f7af13031084b1431edb3a025fc98a68bb036fee7a258b77125953c604ebf349f86c77582fab2ad407b8bcd51cc77c14981f89240cdeb522d062b18de2b0fe0fabdad5c98e62c5c5c38bff3ccad65964d560;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb127e809044734b67104a6e5bd013d16d57c7e1790b789cac69ba3d5621eab56bbab6b7c3a8d1656116706c7c3a514cc5b3cae08fe29012cbcae3c00f815f92c1da45967cfdbc63ad67ef861edf114d3a0e1f3ec961353f2c3298b4216ef5d31a8ae0a7feeeb2f9fda54489a898a84cba22d3bbfc41eb7febfeee1901bdb1e1e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a5d775a7c921d9a42549103c5eafb427d59bad58106bc71e2bf90a1fe6fa02e0ed6d784101be6a13c1c1709b5a97f5e59ff63ca1ba3fa8a6f56315c2fe0cd2a79ebe4b741effc3ffbcb3d70fcf58bec1d1b704567e253a9399d6506dd5b631b1a6bbe3fddeab85d751bf158ac3274a78f0a77f5b07f0c5fa3eb0e679c27d902;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2bbaefeafb32ef47260166031b5dcb508a668c9a646f6d0faec178ab9196b0cb0a8f09fef63c3b27b0f2d1201a8fe2ebe147250b49555bb10ab0d58df0f4fd2c35ada55d7ae416d6a280fe04658aae6697b6a70151bd57e744066c01362d6e7532a229334eace87a36fd79be758ec6d5360a7943df0dfd5fe59da48f4803a43f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcad3fc9bfd8b2eebe7cac25293189e1671d0ee43138d21fc581df1dd6465a3ab5c5d7b946e0ebc5c7777d0f56e84c444a7ba4a085dfc63d576c24538994ba8141ea84c3d5c6456b2d2824b53b476dd54d0d02f57d1c5f35ef117f0ef34d6204d1677a9f116aac09cf344a270133eead284846795381128a8ec8b153426ff0672;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfca9f696e97e881b0259765317d75fcc006ffce3e4b81f2d5305dca6b8e6d19a2cda42f32abdcd5a776a7430d3122c3fe07b9a496693b9b2f9c3e8576b0c6736d96a73a555a38511bce3fc5d8aa5f95e15cefd950df92cdc744f2ce93e89308db8fab1da3e9bfeaa74c793b581a3b28fe21a36a9b1592f5ceaac002469f5fb3f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66549fb3495e5b9be03a80cfeddc8e1df5890ee6a6afbae5ec250a1a64635e459b4041109846d2c30115e8990a3861f0de6f2b1f047f2c48510d5fe8522572923910421d5710a45177916ad12fc6aad6b78751dd6a8da3866f3adf82096efdf9be1aeda8797b77f1e196faf5ba78b2fe583ca7d2a57e2b5fa1995468dd58d4bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab811880726912fb2bf5857083f2fae3a69f05b842fe8fb78380b0b404834126d37e200b4e5477a59b82ba2cbca821dcf73c2869e6ba9f418db1eaad8c37035388b75503e02177fa6591a3ef54118e09ff0479ec1ebf58f20e39ad48cd282df7e887e2107e0fe99ab1293de842e52e3507471b978cccea9122f4f39ae550440a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3744f72d204dac0cb5dd28401995dcc7f16db9b10448e2d8fc492574545d51a7c0693d5b8a4da444686bd8d8f8cf219da968f85ebfdad7ce159058b9f0c0960a0b2d0e83022346eeed4ee907e799954d9b23894966edd721532a37b1e9f3831be611085cb2b476ac8011bd3acb00159b215472bca5e14fd994b9e131c12c23c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9dfd7a438913d4f664989bf0bc6758e5f503974fc3eff0ee78f9f25abe2931b0293e91ac078368e2e0e2b16dcdcebfb38247ee783f6c0620169f62a95328d40c41ee4a8ebf424c558de2aa3b33bec76ddde4941544590fff73f0bbee8f1303c8ab36724dbbafa1efacb0f5b286ee0f36f5dd19b1799f83df77c2cd673afbaad9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c09cff334ca36b38cde4a760e546335637f6cd91803499604a3cdbb7b193707f02d7a2ba6a8e09e7d0b0ee122e8424f1cef72f963b8a84f4f5b5fc51a640bfc1d2d8325a018b382571dea70269831209a06911641742a2eddfe8e7c735d63e7e46f08843351134ab6b45425e9649c77afc8ecf65c97ddd8bd682644a335efb9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfb764dde3f84f4e749eb0887672cdffcb484187f36865b64e59ef1852d0c698e75280b105fc6016029a98310ac282603cf19f29eda968047da5a1977b41bc609592d1e51b7896a1a4f12923f863b18f3240e3320c2e35fcdb0f2056947a0c660aa0403f900c338e731d7f21c2cec20d0f6bde05ae455f8b47782066fea03bba1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd94b68854b8973bc2ac4f5e8e39cf36b964202c9d47ba6ecf9b3874cf8112946837f46d3cb22972ba02574a3fe07f3c07400763a7c506d0b5580dab40e114bab9bd25291719585ebd3b6e50255cc8be6b6e1e73b65122da0a5c51b8d2cbaca00e0f02232083a369888d60cb52e73edb54973314e3ae0aef0f9575db3482ec603;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h987d6601e44b77f5853901b32868861b43c4096c22edc97e9adbc5b4e203cfb3f2bf0a2ea7a6baab471d66688638f080008d6591489eb10d0944062de920021a385b4d49a30fbdde777986cd2b14b5da85d46fcafd0f5b51ca57e49253f0c5b2ba931bad26c7227c59debb85b75a13be234ad337a95580b933467b1375ba50e0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf2e9fe30c48de4d1ce26e8050c9de5c549b5d3437efa3b6035c8ab0953e9057d1954ac07f638f3cfd33e8ae7b49b7b96d0b53dc6730764d214470dd8c71bda3376fdce172a02e31d9c114291e9fe878280d9917e3e7941faa16cbb84e7272a10d2c0a510cddf8d8b1a183662dbdc30ee1876f34c7dfb3eb689adba81e3846d86;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83fc5c05a32fd248e2e62d992b84412d97993a62e2cc5b10f1c2990bbb9181c77b89535379dcf274c8cf9c8685b20bab2c0d0b91266d7ab8a09e042e3625d7eb137a0e495acd1527509e33a1610298152f2d60fb51180258ad7900b282bb2a090703965412bf49ee8c98e1646f12a845d05a4ee5ca5367046d9d00e16b36caa0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf06817dcebcfc12dbb06a7d29f3dd5a65c62137c2f24bd0f321ca1e823580ebe578d7c76fbc02245521f7274efec47b46f3ad1cbf2c472740d240e71bd22cc33f04739a0d9122aeb6d42b8636542d847ddafc6b0639927f6a9631fc01f2d5fcf3e26ded183f075a47c2a71d3bcd4587038d0405bb9c0cdb4de54d84fac3699c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h544fa0f2a11cfd78728f5535bb1b18798c65021561ae52e8401b8822e5686e126a6075c7a7cb6354d4a95ced0e89c2eeb74051265f212c55c7ed298eb39ec0345e7aded31049e6ed307e8fc67151b616c29e873673d95dfe85a9b4099ee90fc63b3d08c9c0b7dd0edc8398e5a27736e149894762b2aeabab1963933cac186eff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd272fdc9425daf59479a8eaf01388ab5d6130a8e8fc2c33d43525a3b6602a4ea6fdcacf492b452dfac28d2f78cd4080a19666cba7e7b1b1b15cf30beb027ff00e995d508a9976b296cb72ca71e94398998d2dc2a81612e00137d423976c1565bfb3dd893fd4a0d37d09b542b075f46d6f14e7009c7a75581180dc7ce44b94628;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha775457287d67112b308bbe86286bb363ad158b7ce4c6c7599d1b4abcd44ce1c464ecf1214d7d707bacdaa9dc0fac019a4ee406ed70e9cd5ce563fe497b2377af7a173af03fc8d3562e1fbe08e0c58a1cb2fad75dacc6be22cfdd849907322411db3f7642612391df31994a28384514bb08d5f37240a127932873de105381713;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h219b0daf03302a791ff97954abfee7a9a24daec451334d5afa33e837361a3ca56a806c9b2ac48f23f1320968a72f654b99d2a9c14e9b790e01fc5e9b9d9114881e8bc6a4cfbb11fef14914f4a7acff1fdaf777c3f25ad2d67e46ddc014933a9ed33700aaefaf5c82f0ea0ffc376174953aaf7a0a6c2840e1a4263453013b14a5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfaabaedbf4c8e9936f877dbc84c51017d68cfeff5227eccc71f7ba0056e069e273cdd15a051bbd71fec21bef966a96effca5119f2124f8bbce32d7acaf039e81d65dd3efd0baaf3594d49442581716f5106fa273c0e1c9512509c775797a797b5e074d8ea3dec17223a76120a9913c8827e7619745174da82370700d34eb9deb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d32764f63bad169942917851da03b0aa22f00de5aa629225311cdb710ba08ed997dc471b6be0b6cff4c9f37404801857e4418f0c0fa67d0cdf9484b115bd5b4e369447ced7e5ac299249f8b0e5807d17ec7ef3ce44af1c6f0232af8a59a900aa19b26bfe2a40cd7b4699a7517e0562b1c9b94c1124eed54d7bb91d5f87a34eb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hccb44b1a6b20c382ee8007ecf55dd008953fafb90763b7d99ecb3a7f03ad3a1d202751a39daf196712b828d4eccb37b617045456dbd8c56cee2649ae0c6847e01d1055825d960ecb01314ce0dffc2f54bac30e6a5d76cf2fc73230b121f07b505993beeea746cb5c856affcc87ff546892ce6460fa6aa1b1a5b4fd481531338b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdcd0293deef43a5eece7a3f21a49c3f9461e9181c50e1c6ffebe94d9a7a0e3d24f82a52e219ca6e8a1edce904f7aa642deb0b1fe62e826ffc9099346b20fdeb0087a0c7448c83e4b9af66adc9136489b0cf89e2de8b86bde6c638f3a873ac938bc4d986ff9a3086a51af62db02e95f03af265ce6669ae7b4a891db47f253590d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he37cbdfd75194c33c4ba09972209601954a452ec571ae9af51ebe5fef8245bc9287b2f8064a64d3478e296382452ca1f93a0d6900d083cfd542aeb4f3bcf6c6c41484f64dd5a16f5d5e7e71d96f4b0041a0fe070dce948ebb9f53800dcb497fe47709b65ab28dd2c6919edce13533a2bd78c146f50032b657b93068ce4903648;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h44958d8eef3ba910ec0973795f6b3bb3ebbacca39a431d23e33c841b247855f9f1f4893a26b920699813bfbf36b40ca9cd01e5670252ea27b9a1c435fbe9c097dde403c30cbf5e717260b616003c52bf7c1dca27ad8d73a4c887d57e49645822e386a67954d30e7d30467c095e651965343dc3d0de5ad014fe503a0be531a640;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4608789cbe70411a35a003c7695f3ff93b84212ff15c370b3328f1cdf135478dd593bb5d0bd1443d47f21c6a62968cbe49cfdcffe1365fdb21081452d4b6880f61549f7072f0e2e12b581cc26fe6e8e322119aed78703e440b158e8cf63ee085240836503d15e2fa950143057c83e532c3441ad8b9f752a1e437b470cd4bd4fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b8a8dc7b52ec8922cbf5bfc153b9700ef153f7e3c77bc412119e250c24f12cfd6b4ac3f4de994429ba71ee229aa57c19d12fc1671b01bd52cee8f623456810eb1146c6cfc9067c391d4dce16f9c88986ee621ce01e81942a04d94c80f3af53687c4947e8284d270e3e8378d6ba563b7bc59ccb8e457ce3149b2a9fa4c1dcedc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b0eca63657d1b46963e50935a9510f3d71adc04e721f58f2c85ce78da971957add0168034c14e06cd63f0dcd3af74260ab8ef8506a1aed3d1f832750045e304c5a0a7fa55ab17cf16c1a72afc52a9709ec1af988a05d418d83b5e93e2e30f3db17d480541671ef4f67cb7cf87e39642a3b763dca7f87a16f4615c6c23e70cb6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78dddda9fbf57241713236052e4779576d65a0e31c50a4c19ea96b9954570390f3d7e5d0568522bf8ded39e17a77c04505004ded3de76ff9d3e26afcf7ab2fb1a0a1ec3ecad1c8768142ff7b91d0ace9dce0111e19a96d3f2010768a0fa273c15920ac57c6ef76c37b9ac7c7c2891ef5f6dd745f04d5f237c9853c47ffa7dd54;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a020f3d9ebb53b260b0b13cbef5b14589a8d47db5445203ddf2778d449e492189dbaeaeed6ec17f8b4ca551befef4d83b7612f02eea8a0fc6f670ec680d37bd09404bba3218f4a7086a6b06d9d0f69bf94b698be5e25a5c0ce1319eb503c421ad648f83d3f4652462a6dc5857237784b12ec541106f5c97a4a3526a43e1b72a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40d5417b699ba4127ae45670fe77f567cdaffa87de5d297c19bb677e89ef68abbb7b9a5e1ccfbbde9b8929b8cefbf879940ad38cff338992eb83749393fc8ad36fbe83ac0f212465e1911143f7e9f3b9326bf21574a8feb1f5c30027ba6c7b740a6a68469b8be4e2f326a0a17f31e62a45590013838b59e311b82f20bcac082e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52f1497e133a5fd083a5e191e68c321cc52eb17c8a28798d70b13210c4ca277c37991cb6b0eaa9ec8e3b8585ca3601131ffb1bf14391ba4329ebcba49b4161354c78fa0aa426777f262ad8768f678e8eb3a1a3b2eddce19432c0610704c55b4b1e00ce851e76cf9120c0b88562336d3465f3e37b115655e7486a816ee8de972f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c587f2d7e5ee33288571a351826580c9c88023cf2dd00f5b65a6c606ae28212240d232f40479e5a6f1b78ec8d8197e3abcee23e1c038605552f5c5053c9e5c422927329d9401915f88cb0e705287f99f76443ec32e4dbdbb275c2429039f67c05bf0ff073ce52525a8c12755475fd75e34789420fae605646580355f9315dfc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1639079a351c04d082e7d3aa88b52c43c2f2bb4ee4203c66b483fcae7839ce10a4d319df8e7c2792c622a700d04a1bcf8daaa6151c73faf9d37715bd18318ad4140c8103eab8657cc4047db4f382a1388adf444baa92b475b1c6b56e8f39b714e8ae2088548868a0f02899c5feaf957c6b189f4224522b04ca0a0c4154882ce6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e14f3f43835c3a2ed7ff21e308c2295d627bd6f1b446329b92a74dc8a44d5f0c15a0667f2df4ab94fa1554f9a330ee991b3d98801a72fd95acbc070b887e02488017214c3662c738e7487a2800ea68c0cba349d6077f9cad5f7a5c1d3ff2da5f79084c439471da738436fc5ecd4b93e69e67a9f03fff6f03e92b6805fc133af;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c6e298f73061470cb0676c496da00c4c5daec8f0632b37cd93e379ebdcbdc00b6f49515e4be7e924ce0386f845f914b65e0475ac3dd9150a67a6e72040cba2ca78c01527975fa811a524261dbb7e97cddb560492538908e7c2e1aede47eb52cdb6622836550a2bede7d6d878c0220d8f4c97730c232f7fff9767e9a0be158ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2aa30ece1f562d5dcef63f69f1da22a91ea38d149ce1f5943b4340e91712f028656838bf22a4ee995223fa37bf1ba815ecb56c650baec064db9c5d10cab2e512ab67ecc7412ac1e53d0522be2d4414a40a307210e528bd4d3c00780a6d1c7c7a3b58d5dcc5111fb59d9aca4cb50f16640da1b9dc3cd6555d15161d3d381163a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf66e70991bf9775165f5f2acb3a85b616c267be0405dca1e11f480f41b5a8074fb6e955862dc7d12c536557925dfc0baff013da56b08ce5c2912d5ab41311793e2261c24d5f7fbe41bec398ca08b6e90d28f9233d0e4fb86d6fe3778a004b7e4e85fb190021e977925152d37acbf6b68568bd573f3901f6d6eb0b048ea67ee97;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7df73af5214719ce3cefd295b5aee348e97b409af4940fab1720512a9aad13e410d56b0d5bf755e40578384267253229c04c771fc30c9ace802b0b823cec4b68dc6a2c7e5413eaa247d70d41faf196410675f8dddb070b9a5405280cea309c0167267164120e68fb458c1f8a90b3bdb992809b1f39a39813ee230e1c1221e4e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9fdd25904e0233907fb5d529ee110d6a4c71c12b95c5aff845dd1fe3fd3d6843f9193b31467a3ff84d9402890695abc2250dceaa03412a6c7f5b83853ca02ec41f795ae4a53df8219fb5fc9bdf41663505937b0bf3232cc00c8d4b0446a152634be9a98484d55f78dd87c3d395496f416549f08f15f0305c040be4bd1bd89469;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8dd4309dcedc991cce30fb2a3b155ff5013d58788cf359fbdc74e2692dc71881204b2eca8ef3e858292ddd0c8ce3d9a830b3cd4928fe60a78e70b9e2a477b2857d93c9dbe5338a7bd887d8f34984b516f0efb70ae4398f761be414c0e1d4988ff7f01df40af96421bdc5515201ae43eade1c501dd75c04244ce3ad65d3e9c22;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h241d2c4c78d2beb39b8f98fa8f08f5005f5a52a653c1ccaf5e286eeca5e44ccd116a2b64db1e11ac3fba69f7ec990f9cf4cda76861176f1f7225a9944503e2f83dbd95917c24e073c13a2f996ec8f80c06cdb18f9712c5cc2072b160907c4cb2d94e2ba3b50c1f270557019ec79fba322c596c5e8ba0b129d0aa5897cd212144;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hefe5c311301aad14f3c4a25fa7946e2259486dc0542bd49608c238786407230ce0f73326b3e36a9a27bbc8a6d8339d51dbea08403abd0e27e7758f2355ba2e1a9e4ba12e33b7edce2b0d3e35e42578b37d0cf9a867fa2407bfee73938033889cb8dc68ad1e761fdca78ab9c2e247293549b81e5b40f2d73c9359c22575eef19c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81513edcf7311b5fc0cb3b01e73c7749e728ec392bbe5dede71467117489258e6b789fe6b8e92a12a0157bea7209fa1298836a08c5343d8743c9f80bde154763ef718913d3666aeee40a651cc7ae70555e14e37002196243bde8826ea03c870a0ab1bfd03dbef91f82e08a3052c9a2c02646e52969804b3dd72323d8fc419937;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h780394e8412a31da7f3905d2c1959ac7c67eebf659af30652e9976c6c5ab9b7f00c5ff5c2b7007338435534f086da573d7216bb648f185f727526b576bfcc1c95b472c0e87a30083864cda5a10d9428770b10ef54865b2a0c7a9a4b5af0fbe3b9f25dec5370306d3f09d9e0d3b5ca4d02e21c2e98d9be061e2d5e0f32b63d576;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6be78a9d8d79a53719ca9842d8cf33447ccd4c7889348cca47c88dc52372260a623043b959e69fc3ad033ed39bdb6df3f1aec5779c8298ac88c715a40445d1690b4d20d6d257e529c4b2f4cf841bdc5deff5cd4a06964402122a4f6f5cf41e87ccc71fed8130b02f23599a8ec425abba755c70dc381e8c8548945e7351df49d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h279004d4488410388bc693947b8d6233c2ac86d1fd0ce59ab905d1f18931ce55ee9283272a4f9c30455260f985ee473f6953023250375ca8de1bfb0c6213814c1d971acc59729adec7805f1cc9e30782a9a81d9e22fa04585a7d7697fc0e9e3a7874f9386a638af248144e27c2458011f533e165865ae7899154147da58dc373;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8b0960fe80e4e5684c4306e6e8fd7f4b1f23b97e3a844a9395146f1a0aaf49d433b59e0fb314f61ddf9599e2089425f8c0889042709213e4c03676a7626aeb36c480239888d6ef1c9e9de72f8c73112a93c61a25908300f800efe8697ff1a8466c71dc8487c1306c29fc2f51e651099f734b0b3b21bc4fb0ba23bc4e1658958;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed683b83d7600f3a751485ac9617e0fae302eacded5ef20d26a0758504add748a36e9d466becc794367411a0548e536654d1c3f3c785313b91f7539809b8377d9d40227ae8ae3e1f4e2b66db905c8370fbf2ef4d41f2348d3440c4d842dc71ff0b7e1744075a0c6d7439c1190e92015b0c8e340253668cfecb6b081043f8b2f1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'had9410f8d84892a91bfa7fcd71b542135cbc6fa63b230c05c02f9a9097901067538be925f02d7304d179fdc7f9fc6d02380d9e3ace21997b1f136b315f7d44e9138d25f08d62b51405040ac6c1e096b180cb89ebea0b87b9a73cc2e36f9800c81450d3e01b344e17a7e9410432aa60541c5d3e68fafb2bf855263178e1c0caa8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba7c413ba67aafad15532d93862ece3da75965f45a027744fa34fd6e05c902ff246a0c07f10023a694b8a16e19abcd9f99cc06cbc3ece29faeca577548b8f4e684a0204adc784e1f04e175ac5c69ed1e7e1f86e9944cfb9297829c8025e61dfa382000b17190490a032ae18d3b97e7cbbc1a716894127cdf4e2bf86b5d9e2de8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61a38bd1d1997759a35420deed56539c97be7f9b30420b37087e62741bcf1ab3cfa7391801db3726e188c585bb4b5c44de614f1a9a76b3396a9c853e26de55a8f8b00ec268b95b65284933c19e8429860a23f58014c5992be1d26223b11f0510c52a5aa39c311cc2441d4ab7eb1162c92d230faf7d912678662d7230958d5673;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf731dbac9ec25d69d6562eac23abea3e9534706b2e6c5576e17c11ef3af3cff05ef994bbf24dacbabb1e2eabe5af82dfff6e2458771e216cfb2df5b01d9e96ddd7f04bddfa41549da6cd24cd5a6a7f251ed53d284dfd6b6486a53f336000949631d6e4a1245abf491e56f52f2910059b6bc9c48cea6cfe9658a703f544519c07;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8a5e0d4eaec1d0c1ec07a9078dbb5d98fcdd06782cfd05a7c016ecc53b38131a2bb9530efc4ce8f38bc1205c8ef535d826905a30672256181e02401c22b489e1ae346ed9f8b76cbd403813c335d912df8330013b442386698fd2337028ad32c431a43325e44eb46f4071240e58208aabb299b10504015b4e5b21bd729d33b4a7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc0d0e2a5b21a524c8f419a834b52eb0aa6da0f4dc35e02c65f4df393d4fa0deecce8d470a75aaace2a55352ba4020b39189cab249b8c232de52dbdd22920c9697d8e611cba44c26c6326a8df391f6ef7a7cf31235a4dc1a86b26bd4be1312731ef617c31b9eec1229bc9ddd24894cf5bb58b27c9c9dd44fbb606418dbc58f816;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca0af4946dde0fd782d58772ac964cafdb7c6dd7f3d41da71238ebe7e61394993753b2e7486b12634b8d63315425be0f006061a6aced0d4dca886a3700b68e361568d7042691ef0a6ddbfe5f374b998350d5e07d709fdc5eaafedf7681ff05ce8002a80891214406b5d986b92c1305dfde53b6a4f064d5a932c2d50b9e8da5c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h830b7233c49d994a3c3d51d50210f5854c63d2adfd400c10b7e8c8c3fd44b615e0547ccfb81a211f65f767b1fa51bd339092095045cd9a7e638986ef352be3289ace5e4f557ef175e37fec465094db2d153ad1987b2b94e11cf678687fbd852b640cf747fb80c0097b6c8a994a624138a7ce0aac9b6e99572818a75f805a5618;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30fda5bc944539aee3e204b125b8f678bec4601ce4b6e9011bd677158d1095b42958307f78036f752304bd3f19292ee3ea34202613a3fcbbc3f5b77c92b8edb9875c61ae27ddd58e6d219332b7a4047ce3485b9ca7ed3560a1c9c5770088d2f1126c1581d731d207b17d41ab13ba15fab4f05370c69fb68d22015f64cf03cfb4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19c368b6bae2bb51622f08d7cf2f3223140447869d702600c1c3503e720e9bbc6c00ed874cb7f70c92a11473134629193b87f964d4f92de3391e0f2b3013aea7478075e5effa590ae4382e62456c2acfc58c4734692e7b0d95ba5e25b42e6bf9c0586ab1969a0ccc8b9944f33810a5ac2e855a5d7cecff16f1bb9b99fb5b1900;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h637464903ea6b0d283e6842c333c5ace8dc7e32c654a539fd8b4785d97e66c964664b014195389bc549b1d2112883839d968a8d73581ab35dcbcad5f8201b6be6a8023ff69dc89f8ba444ff3dcf7ccb46ee2085ed650ec79af00e02b0b636b19d5392eed3b0352e4b272171f68d66f6876631fd555b305e21eec50ed01bb72f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfdaae908b9d63a71770bfaf939a801b5482710713e7ce78fb9a122bb0e3d063ba1fbdaf19d82ac325e96be7d608937d7a2d6adc47e344581bab8229b26d7c33e9250fa5d36dc888ba01e44c6df15bfca0559c1608f4ad83d4c29fb1feb7d49aa68ad186e10a189a8f9dfe6ec982d04a8d424224a461bfc3f75bbcb47f0dd16bb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3977a7e941e7f8eeefb555407fda2056a02bea398f9ad48fdff54bcdf731a47fe37fdd2f71e44330bfa9b1fba0c28a712045ef6b16b6541302d11acc0a547707355b398deb42ad597ccfcc6fd34f5241d569fbd0c22a5bbf6ddabd826892d894553a458d0eda1187537e5a68beb44565b609c3ecd6fd6ffbe12c93a288367b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c0893ac3788970e2da191bdd92e989ecc247c487ef34c0f2700f1470b715f09090f581345bbdb03e4d651b3819f0105eb8456b51b5df2453e3ba01bbd5ad829dd50e584c1823fbe7d55bb5c8ee9fcb549d6ee6cc9a7c3641bc6277afca8b7eca33f58af1ea46e4e2e21f50b9065ac8a18020d55be6d3773f8e322b4750e465a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf587d6a56ab4fee29fc3d1a4d8f883776b64ce29ce9d3cd1a9339d7b810373c838c5b3d850ad73f8e4b4a8b851e30a5804d66062cd8a49022f665079a732d5815895d78851fd25172a5b875f06951b2fef9731bb7825c68363c01f7f41f373e5bb6304943f9770af500a5bd8fa63add074356b4f07b98e7eae2d69ebf6a00111;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30315b3f3267c2b309bb2668dbb6e4a9d5c12316406aede85f247aba47bc443cd606d649fc10a2b5865a23622c907a14d4d39e03a98c080740dfd25c06e71556511f79a0ff5aa67c8d41368433869360ebf6612e4ce70d94eedd0ab20b73948daa3d53b1885eaf3e7306d84b2608616d717d4ba51307903e958add031d9118bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8cab0bec1630fa138e813a6d18005fe49ad3754e912489f6b401376ece99195692eb8707941563a6c554090fd70df5f61742edf74889c3eb3685e6b52ebbac5382731341f86338a67750074b3bd4097c97373e0ae083786e38416a45e3b210cb4b6d4cd6330e796cb07490a312f8205726bc156bc1205f41583db0d7e2e50753;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2144e83f6afdba0af8376d54764714ae2597b7e348926916bc0281edfb68746ef2e4712ba7d432374e98497dc9cf313630987492f3ef2f6e1549a2c2701ba24a3ffe58ac29877bdfbca142b679f4bff2636149cff6ce8a0eaffade1894923fe260c39b84e6aa684673a621c7d9e1c2a1efb0f1e52d459802109da72f467b1c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf7dfcddf27d1fc8df80ce3d70f34d9f3b45175b681c008880e86adfc8dd1915d1838ac06cbe6233af941124314f6877280d150106c3900f17c84770c2ca8b021ed94d63b4cc8ea5ea5b2b67a8bd95790eec3193666286fa4eeb17c2055d51200356902c19ed64756f6d5ecde2aae349b6aca7b39ca1d7dd359c1404186dc9e7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd173f27c62bfcd247ec6a51cb33a22906199a611277bb0c8cdb2391009d46e0f3a320caa4b08e56a0afd3adceb81d99bafda7a86d52b1fcf3785a4a3d0eabfe0efd55e54f9b332c7c3276d489e11e248f53cb310c76c45aa9f82a18dfb8f163ef756e3448095f4d4d456c6f1aef7887a272aa10a20d15112e6d0305497b9497f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7a0ba7101b039222d5a2f903c1284fb9020d60ffbea5b6eb27f8a87d050bbc50a082ffc166b4f3f178b77fcb5bd2ff55f078b050a6e7f942da160f372b591c479ee512c73092d125f39e37e1f3ab5612e55da9c62c7589f3ba329c5bcfdf9e48e548beaabf4770b2bafdf3e87515dd163e9b18504aa1711b33449ac96c66b76;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2448fc9e525aa936c48936421b0ec09476061c626faa06ce78538ad32e99d996624f4dc18c5c0fa0d49f47ebe7417751d092d18d2586b409123d6b145ebfbf14fd31e9a1dc36bb42e0ef7dfd5e26df93edb444c8f5ddaec94d5c6b0f7798444c8d01fef07f8d710765c5dbff445a1987b193aecba2c3977944b3d2c79c5322f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h546dd9112900ec17bb8fd5996e7409b7a98fc84d0d24ddb706d419257c3f8cbf955dac097e68b3c68115cfd733325f5891dd51e2b9fb12d31375a58511cf83ff07f3f2555c6db2e8734f060fcb7d68f12c12e42d9e05700782d0e3a86558e196bc355f04e4e7df70483388ffd8b46d29da6fc54b15122ffed642eb5129623525;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c7453ed65d4c598f0977915f440677088b2ef5705419feeb0ee01a81fdc0c60ddb8914ec4b5f4ad002c5949859888c559cd3fc226bbb922ef4f8727503e536f06ce50ba548778c194be7fdcb5aa1d7de4c7815bf675ef82e551f538d18a07ecd7fefa1157ba94ced74a5a0bdf02e2d9ccc99d4391bbc9f5d0026e22cf90831e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a397d88f76922b45fc710fac0f05fc70dd9b192139d292127cee9e21698a68520ff19d09068053705bfee32888b9c5525530ad4d4288358648a35f1778ef48ab89f6facd3cf0b72e36f83c3fa2baff59ddb317847789a8052719d8ebba1b65088920d46ddb11c843e957b3f5f0c5082d0c1a46e1b9b7046d188f67ab2a31539;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27d880845c4470e0f683c58864a7b1555a1020e49f0e3d9241928b36ed85077dfc81d80b2f5194cd2d994fb9483aaf2b1d391fa678ef6c157b6f06e756eceae722bb2fc56804baef5d9ab07b41927cedc9c0c78622552746ced959a972708d525d6bc592628040f71e0f25e9ac02f551768a8a4643876f58ff2360f1bc76fcdd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82f51a990d6d1d09c3e18ee7b9bed7534a2d5a6376ac6d524e4cd38ab33014028731959a3abadf22462f6a092189875f683d15e5b74266a5024ae28a4e41c714b07b1ce0b23be05acafb037f10fdccd5cda86955fc0c8f0d8ce0af401b45f13a6a81b06fa155b316e8ce6e61408ac827710fe86cf661e1bd48d0dbaa60b20fc5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h77535a3052262c55239e904e2b070a1118b754cdbf1d1cbf7a8bc811022a22c840849aa0ae2d6205eb325d265776606368a468a4b7243f988db44655e9c4e74af4c47992f37c846143c075f1e53338d27025777ab767b125be238a91e474d3c3e9cafb3151ad4062af2e1e65488fdec54520faf098b05c91d496cd7076ea305d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6fb6a4cfdb8ba6de89a3522917336278094f4ac6ae9e00c26e0ac66ec70ace66db14ef799f07ed5178d8e5cba1bc3466381f5d2b62ec30dd071bef47e138d40eff2ad43b6c5e2e7100156acc08df7bdf45ba6444e42934691f2197102db4197b86bad73cadb956efb8e66d859a8dc55940f474713850a3e09ba8eebfd6eb8b91;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he0f73ec652fa005dae7b9c20aa73f38f751507fe0d1a6765a75d834bd9497746bdb0f62e1f9d9311855534c262b1d9213b6b5c6dffa7c6ea6f44cd6a037e1aff205d5340362ecb0e1a18b5d3a6de078d141edf8aafb7bc6052ba3907455bc5226ca3cd4a63e44c77fbc57370cd594f0c4837cd74ba1247eb884bb231fde27c38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h402175566ee31edc637dcc675202644faca6a7fc673dbed23a7ded4b6696dc52190c09c12c3a5fc86e36fa722cee64956c28814e6201855d1245116036eb7f95b40b26b2eb05c00da9b6a5fa05a7658b55ddd0e74c7e9dba9c75158a0eae7a7f0dc41ec608b42f00045612e9620281f456854000c21f9dfd21b63005ababff24;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89636abfb9654fb52a9ed3cd39c950f858d0b31958f67dcbfb136946f006bc4fa5c0ff1cb2155b5330205d8e299a22cbc1c280eb19479b927e26dd3db67b111118a9677523ced8dc549f5d7bdcb5e4a37f27e5c1707c00dd53474e86d26f87ce30009ad2e467a35e5a7f208ec8533f6c65e999885c5566a0acae6056e01eed38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda224ef9dd53a0ca653d13085d2bcd1efb20bfb34e0c29ba7b4b3a85fcf69f6f7cfcb55102c4b2dffac32e2b06bed4b644c4c01e2f1407c851639e1ddb8f72def9f9cca3ed45527c462cae62df0c3fa74d67d771f8f2508679ab4f6a14493a5576531a51869b2abda1c617963b4348a12d8796fb62e79300e34c7b9d96a09338;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c654bab3cf0e03fe553cda3f3409a78ce03209a0db7e025adc881f252c5098c63047bdb3654f90cfc76ea481498e40ada13c1a8cac946c7f0678ab6ca5929be23a1a4865a53813c863d548d3949a0b3c9339944b2e61ffc786a7392e1f4799cbcdc2d797f213af4b21bc60cc57d6368381b1d596913c94b55f5439dc08a348b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73151c361a773f7ee7056cae07bbd7b949b3f212ea80bde178d5ddfff396312a7923fc6400c736ed9e9e703ae85d0b920a714af1b48efafb6f919d3a251a5148f22744fd29f9646b2e4d8ccded0083a6e4a306a241c38d85569fcbd5c03bbaa33cbdca76f94bb6d5ce70eff29c626a45d626aee6553782a7be8d66d2a98feff2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he7c0c1949dae9f84c19002a1d2fd0ce04f26ddacb2a0631d1462dbe19eea4297b9d3e1c8426604673e0d91961fc5e4fe675207eb82386873026fce3b9097d02bac1378352d5ea0ebea74e869951df943817359832bee4ce95fa534dc850046461ce6941cc186841eb3ddc98b4f43ad5008eea5a47b6a910fea890effe447c54e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b1dcb679abc00ed48c8a963990faf1b6b158e5850c5a966cea8db69955c9188f9cb7f4391249ecda722bd49c4fb3c67a51ba63589bb77c566176980c1e78368af6adc1d427607cf7e9e1a16c53c395a4ac3c53779814586c3deecc49af6b5d3462d20d1088419cfafc519dbbe22de4a4a416d7f8ab1c533ecb8fc184384f4b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9bf8630a9c28160e9100ae54e169b270c5b5edaf619575f0b7b9c4ddeaaae57a5bdc71223a2bd6f694b4529654712cc2a918d5e56d243e56251918a8a40ae04bb6de0a2b99544128ae42fc7a8f2c609b5d0b653b3b28a4592bb73236059c72576ae013ddedb0609c37eb4936c9212943ae86447eddf1a05c46d4d822795e7813;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d9fc9ab21afe309fc8150d2f8b38b21dbf189d2c5e863be1fd1ace28d21a9165853cbcb2d23f466544d5e0bf6443bb1d3cf66febd534ebf0f02e33d83ff636ef9d03968099716f607188b36562e61a46f9772e91ebba931adc6e22e96f62f428a336dfb77975babd0fd89d20ae6fed6506bc8a277e7b4ec2353e4004bf3e402;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9402332a3a630254b30d60765d711af3a380e43554e1b9f97b7521627768d5c68f393ac95575d51c53934b3c95853edc296982daefc202beb2ed1186b7f96afb894df67b4a8c1783be60216e6905b5a193b4dcd3fddb9f422c47948980358add05394257f4060071788947be3196bb4e57b91d1529e6069bf23d06063a5d8d17;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20e95c4d86a1f19e547ee118f403a43d01206ed4c923a3ab122cf34e44e5312de81de90fdfd67b58c02ef80c1c56a539b0230fd0aee09d018bfeb234dd889f187155d360d9fac48e79eb81fa4bdc85ab5cbad0e0c03b7ddf9e64198d50b49b31941bb59bcc2fc059d9967c7c19aff0f83169007bd33b6de083be6cccc7b2c519;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h240ec32db50677a64cbb7f7e7326c97e8cead9ce5e58b3b3b2c5647e9f47367e4c3ff1c4e3469e6dff1518ecb8541c76842b469baf01cdf222a4054138e00e7acf4e2059ea1a07c22dfe1530ed537a0690765916126995b6810ad365d55731773dd973a018dc10bc69162f7582f0d06b0fdda1125c7cc7164c5e1d2b93971bf9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf8bdbb42d769104b7ac89fffea8a8799c9716c29487e3d4c89dd4bbb5b14a86aaad57824260fbdee5bfb2c8d379605d53f732a15edfd6a3f3dbf2af9d1dc3e9c226b12a8770fb68d5900d51b7b3ea590e8cb495deefb682e56ccdc25f1fd2da3273c9f8695d51850e4e8d6955cff049fd2de38650cf980f33fbec5b554cf6ffb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88df8b39a899a0b16a3c3c0b2c1c34a4ea3b04cd0af2fb01ecc19c071940856d7b2d5c4ff70f83e625849941460d85f2952fddbea83c01b6abe0a35f2038e75d166b7c381cefe3d6cbbbd8ba37b63b723542bd53b338c45c165705ff59531172bd7e2c2c251916dc9d578bd55f91f2a39c665a5164ebc58ba6f3d86b680c15e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7cd5b238641ef425093b4bdf3de18a1fd8ea799707d13725ec8a7a602cf48f94207135ab663ff7b61ec962c851473bf5558c08983f49cfe9282317871f92066501a27ffc8e7e962e4f848082eb6f16054be3e6d68ec957b768b5dcccf84bd4b3a9389d068706e5b73d114fc8b304d62c06bbf2e4d375a4a4db40e2db6d047b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd1c0286aaae4c744ac72793cd9ed5dc0236c79b7f811f87c4cc78678ae715e499e04014e345c1a68f4e355efcd46a9c79f31db0c5e712b0f3783c5fa7ae3d62507be4ced989dc4e5f05a63975e1033ad6cdae78cf6989f8cd7b4b4c999b851e73a5e64bad3e348825fc4850a9d705c096bd5408a813b6154a4cd04ea58e54bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf02ac650d26d84867ecf95fd7d66652ee9666bc80372878bb92a1c6e72a4d3e16d237ee065753c284dabfc90e294d43df535ac179d8c5b0b2fc449bbff5723af8b033252a50b9a754425f4a51ec9844c40eaa8a3f0ca0b0bb2643878f6ce9d6423cfe83804fec0d455ffa7dfa07b6ba8c49a696be0a29b6fd89798f485606252;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hff410919f9d82ba5a715a526f9ae00d22ef416c9f96deb97c541e87568bcc8c47ebcf18d2318764b4cd360eb882100b816425862e0138e172eebf3881078560b1960fc1210ef570bc04afe4eed8075c01c53dbf30646980481f33f5e3330617572819940945612ebaeb8f9124a689d55583f70913bc9d3cc80909e048c73a7c5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbcbb8b7e2ea6137635fba6abd10cca4ade97033a641f2e0a0510d8b4e923b0bbde5277e6dd391e49e165a0231cec92c1e77b2662f2dc27b7ecef8fb180d15051bf831d44b90d5f2ac5ea72a698372d94796a85936be2687f68de44a35849c99972b10f31ab578c95383fd31d9181bf3b07b6162edd2c3777de8a3ba92d2d9473;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc854f8dd5f79f408e42fb3be1e3e7baea092f669c36444a205560485f42984c52384d37c87cb3a90194a8beff2f9cbde83555d90f999ea7dbc20b3d52e14aeca67e4d6c4c0decaf64ebd472b0c74adeec1da9b09aa5fa4c6f411f35df8d994621daba7369b192a74f8e225fe76e092db7386cf76c2ff61aed237160440fbdd94;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heab03ba90eadce5339b159151a5d2fd67c1740a68a3997a0f6d9cd39bd1744414a29c0de6c988b7484be23903710b6f39ff64263c02442a9b79cc322d5bc2c610a0899b454af5b07ecf301b41e2584a9ea20917000a7187b6905fbc33672cb56ddfb6ae53b8d0226736ce3cc81bb7cfbce04e3edb98c0ec5deb9d427c0574c87;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b5710539a3bd0e3364528889eb7ed90e54fe14bb6e718d8a8d41c15ed9ee91b597e09650530bf60d1a0c30bb691cd8c6ea4be2dd7916ab41e8741d1f985f393d0af255ab86780e8f55ca932c3676daf71d105c8e7d5834f49dfea5960c74f71d638af500ba7835d6db5631747c2e9736eaa1ba15568b00a89d16aca21f4909d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbcf51f5f4f9f113d0869fa185d7e88a8b080197c56c5624dc23bc23ef175cdf30ab4b9ba161f166b17940edf533fa72a1873057d4082becdc9b49a5e8f5b14b1bf7343272131f3787415c3a0a985bab62169c54d54a10c88ec9a1ac86f18fa96b4615529d891a7e248d173932134849cfb86ab84764cbd9c34d3164684c448e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h67338c44a91d0583e975160c8ed58f0171376f5bb3962ec92973f78804705a2609f74903307103350547b126a1fc85ee87431be8befd4a83b64f8eb3fb8be873e9fcb0b2b265071b9240c6b9d4b3558b24bbaf562ec76b9b3f06b0eb2e9e84341cbc275c6ed5c13b30e2077b3f2dfa47eebfc551ed88e91ce3e575a7995211d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4b8291a00c6fcce5308bc77fb507254d0098302f74d150890072e13d998eda40a965c337f1af1fcb3db93bb5fa9abde1ad9427b4390a3ea70baa4457a3c2410fa24e7c595fd0d7faeac4aaa576d36c45e3c7e7fccefd7c7945fc6257e16c560f177d208961f1e6a05f36c8ba47c3579292df2fea5cc87512b1a72ff2d8d4edb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h641c7c4b4294803ee8719347be7b97db1821f4b848de1fdae34f9256252b941e253e35288a267ff7e19f8bac4adefb45be1fc89852616fc5a07b4c3fe6555df4f1d30f73a04055908403085d1fa5acac88e6852f75f2ce1424ceb84fd72299ef175a7b14eb4e4c386ac5acbd47b60f8ec49a7c86da1f94157e691b45cbaa88d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f0beae344d66c0c67a23655b768cb1f92379387ed663f23fbac12e5cfc37ee553915145ad7f771c0ded7988ffc87af9555b7b6ceb610dcc81828cf8a54e5a02f71dd4c0a5952c0087d622636da9b60122d221f31233b39c50ab6addc7da184e136359a79af528bd4a0e8ada5b8098658185c6eaeae8a09fa13bcdedcecfe135;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h128fb7eca386e9562809d055b9e1a429914f6da6723d12b7f814fb303d09f7f0d66c203bf485acdf585497a9b8549f2c255ed0f9511ce749148e293e9e0e5aee8b2c3bdb99ad349792922c54718e0ec24cf8f04f5a5fa69d784e56c0f75e4fe7dbb5c6fff9a2dfe88b79a302120a4940f7f9b4c8c83dec034d541e9c11efd6ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58571b281ce7fd59dea7717473b99914c1338af19ca748c14ff0c003ddf5ab950093e3e0a28596eb96f186bc667053a849ec276d2b7116605e1cb73fa48fdbce764f8b219ad448510ac6b4a6674b710be9e1c1eea08e22378d04e39e23f3f4040c48b6e2d6d5396a1563b556a8acccd8d50368faf90345c004921ecf531f3d5b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7684b22d97f607e7c285dc4c602bde4836a757f02cd17cabe45f9a5a60b692f87d7cfbe5b3fa9fc3ed1b61cfa39682929725d1871c3202795ed0919fb912fa615481d6ddc5f2a8f22a31427ef0050ad4b0e698d082813871423603a2a68f05ec89cebc302b43e7a6a1640c7af52748794cb892c27ec14222ed35c7ad2b0b0083;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac1b7debd088408520ef81a1127ccf213ee5acdd76bf41d2d3031d310bdfe5f66f8776de28d728578ec199cd36e39c1cf854eb820be9aac78a4341e6e8fce5b01782d5689f05111c9ed4b951263cec9c883474117459752b9b5b5b655a87a92118d9bc84606526bb789970594f5c10f51f27b585d5d255f6fabbf7e26308bfcc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c810aba9837a7e915f6df9a28c55691ecb45a215f2fee99bda51d8722f5f82818ddef5bca98302196bb7f48bb0b3bb9ddd38f129158ad24e7cf489e5a1325760c657788fe5613053d0a2dbdacaaae55df5f014711686c1fdb366b50afddcd25ce5fe7e66535887cb48d80b82a99e33418139e55c40795d8e71308b7a51d4dfa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he191b279b60188986a68de80f02f7976960a9034e376031b0c1d4a3983d51f8d33f0139dd0f3d0eab45f0052f1ea98df8543b082b7cd065f0cc28b4a30f67357daddc41e9c12fa8abd1e5792cde4ee5a416bc9c914bf86f47f7208b3c1844efff8411beea98f29c9502ad9965e9e7dabb4449035174ec3a216ec6b1c7b22807a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h99048e206e8258ddf160b4fde760ce990afb8da4e32607e5d65593912ee7a495e75f6501ffe65641b03c4c5524ae8085abc7f266637dac7c844a3dcedb78b40815bc1309c7c8cbb0ad1f5721d9c4b2decb95e26ca164da592407dedcad613fcf4af1ed95b730edd92efb415554771c57312ccdeff798adb9b3eda9bd3f2c6123;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6fb6cb8b3db6cd313983e414db747762b9e75437833310a9e8453eb4279b3d469544d720825e0601c368e4a07c6e5778d5bb5f7932c2e5056fba0cba8893af913dbe06ca8f412ca55b0a0261d6a76f34ea2bcc87d9a5b95e65b842b9715ccbccb9b7a32aebf36c896fc50fa8f358aba0a09225257f4c870b5489fc92af9968ab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d1cd089baeebba13159792b5bc57d6075b94bd816a8bcf3cb6888a32ff3c7b35251b8bb070fbe9699175abe9369ed672527dfded634fa72b839e3b356e81a2d5e48fa0528cca391a9082594221ed7346f18b45f47f6251ff19d6a755cfc6f5f6a8df1afe5f140df18425f30ec9441f36a35fc64419427e714767d48079aa655;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5240405c82b6a7b1477b0ff9093e1678855d862cf93e1e8d397c0aa9717538158ad7362f1de6b8f8a60fdb476b69a897a2f37ea1a40aee6e63f503083cca80cfc7058f3929dca6d33ee57790039e4ff7a902d4c9d73c5b8dfbdec7188a2f526b42a588d8519e29197b4ba15fe4668cf50a7aea94b10bfda8d9fd97af1c0219f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4537ec105db6a310bb03c368d3ecdeec9ea953ce6a51474339a38eb5eff6fc04d1de6de339f9242b9d712ba277120e8b0668be0bc9067e5674ab86c4be2367c0bc78fc53e3e8684bed38235aa0f7811e1981e23eb2f4f4b6d7f9c63792437417f5d49e2f3d3090036b9fdd26d4ceb2598c0587690f74fc31873abf129bfd1027;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h92b7ceefd44acf3bd7aa6397767a8ae4e1f1f9d2b76059f570c742f2ae3ae1f2172b3dec01ecdf0d1973a1d5479ad2c2e25354cbc88c2a10e25f7d20f4a03f2fcb1fba6116ea6a11dae1a303384e47d90114238821c5a72380c6b6747e5a71ab4a1169a4cb2ece05ffb4b0fe9b83183cb48559b401664d6ca88377fa225d53b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h419ade8c2f656c794215bb1c69731bbb1a37f7d430277c2350b7d77ee3da3853f5386eaf3b59787b6d52405b3684e2d3880edb87ebb09f5590d81c04a546c8f680037cd5ff248621b3b448454236ff2ce0bb32600d1a71dff5964c7801057fde5838f495eda9dacb3d4a2cef611477108cbdeedb01f4ea71b78d780d7f9e0a88;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd64cbe48eb57945f373cb3bf294346ad019560c291e4d9f1fb523b523dbef6087881ff528bc01ab39eaaa6ae53e98646a2550cef9a6b536eea7b120fa55e4237b18a37cbc1942d95fe567d90e7d1a790458035093697070e293d8746ab1db964b6e7b2fb5c50e52848b6dd3dab3e1aba0271ad021c09e35f4a1b874e5617a2c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf41c802a3a66e8d43fd82b4443bafd7902a982dbdf9ab61d78bc51b9f1450166cd4d215b9b44d4fb417e12e25cca9f96e88256904834fc1cef756af91508a7d7178e8ae3174b02aba3618d291b9c1d06324172427aa6b035d18d783002c7fbe12b070f119811d3c7180e0a74883351baf3b76c3cad6008e1d90fa92e203c7066;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53ecdcb9461ba3cfbf89c30a07ce7f12f559946161cd628ee8bd0b73090a4715c673670e571714af7ebb33d84c22a74c987fea6b19fa5ae437f568e1664e4577b10241062b6fa5db4b7ee3e5d837e9755b3194180fb5a7eaa3f92a18b9caffc847206a9e20b581820d92c48186259d26b6815c8de4e25d7a015631a764ccb31;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7be7dfd38bf9696d23a81975fa2216eedc07b133e0194b982819116927e29562546a57b951e7e38b7c53469c82ea7450c0f446b9bd267daa1539866a2416e776236f8d0f0ce51cd290528f84954153bc8e80b9b5f4743f17a422ce49ac7afc0aa6cee27ac0d0332f7a50367fd6180179b9dc17ca7c0473ccb0331eaa487af8e7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89df2ce538345a42522ea1ae9652bdf65a3eda117a008ce3c8312bcda0ea7dfb198928b4a40ddcc3b5283c8782a77a87c4cb66429396e004d721948114a044349b90da9feccaecb9f22d33055e59ebd08365370217632d125c0cb0634fef755de06a49c772031847b2b9cd9f32a20dbcdb27847ae36d5b6277f8afe5f36d8c1f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc7c971159a4179f266bcea64c4918261695d16f883c2fb2e698bbbe2ee0319001b5718ef2a53abd50a7e1dd811944861338fc0daf51e1d92f697d2eb8490b09e471efa3d24c4cf02d5362bfd238771ab5ab8aa9cb02c04b88ec6af39535626b8d553aac0a9963df9e1c940aada0cb9f099b02e14ab32ec1a07fbfbadd9d2c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h714acb55940f18b04adb4092874fb26167825a289b6058c419d0199c887767c0ecde3826f9ee2725864910dc7c6a2d2688c5e0c54c477346e97c0a7788b54588a3df05689f3699ec2df1c97c9ac9021f95eb42fe842b0b5572fb5a0164e23e480495e84c738ef471f0818f501c234c483efa56bf925bb2fbf97b9d692e5696cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h634458bec8430ccbcc58fc8fc3ef6ad770096595fdbc47917518ee1ff4c4abfc1ba1b365df716669978a08109f60b3fa5aad440d67b7bb8a82f29299ebdab31b7c8f37b91f5fa04b231f8aa49c2425fef9a2b9f40803f7559159a04284b85ad19bced9cd74fd2c572179e1ac0fa2eb50d71d8f13feafab947a466708952c4886;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h833e4b1e3ffdf15f9d56ca75f402050f7e5b68aaccdecffdd69dbf4f34f752358069587c3559eef06047763368f875f0b73144b09f06797392e7d943068c2d69faf8ca48859c44846c2c4eac0d2e54b876d084c6074f994877dfebc3b0bd80d654932d81ba61e04fa18d9ca5909190d1786fe2e37c41997a42bc2a454a35a4d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa1ed067c9e5276cf3ca54037c27468aa61269014b73eedd690f6db94a527719ce23b27b4b22c898b5d8f424ec3078fc1a9c267511beeea693f7dd8c775485dee8bc8763b3d067f7204129a8150d6de41c30dff1b92764751a087dcc483fc3fb405a012a52e7f7b60be7a465df5b355fb4bc07a69ebcf1a1a150c77f32678d6d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd341114bd87df75eb7000e14e44896aaf370d7ffe1aa8e3345b5ffdd1406bea1c214310c0eaefaa920819943f423595ffc721c832e3e7c412271acdcef39d62a49b6dcc32d9dfacf97b6a8165ae85dd96c3bf850bd6ad1ee145f0d7c7162f836792927e4cbd16007c2518cb7c9109f814fa9c980b7ae958f1bf131a4205541e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7bf3e9e89a455d0b4695e2a261d2c125ea637882978c71b62cd82b1e84d91fbef7471142fa1467955ea030bf5798e041cd501b214c4884d9ec1980d50b9400de22225b4b6593049f4117d740e93ae68469e5926b2219ec75e9e0037ce04eeb3c66471ca3b4af9b4f6e01e434fafbd3635f6ab8b78bf85b0dd1fc24465be7a8e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9cb9dbf98ab8888210788c923aad3aa9dd56094aee3fc84b2275a45efe128f8c6e1eeb9dc1b7751cce7291fe082ea059d224fa1a0426cefaa40604c5721910f192770061a814dc0b2441d99173c73914e36514a41bd84ed9e06410f8bb549e6f900744578ba00761074820dc95d34e651d3e68c74ec0a38fb3d3ffbdb6e590cb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf5be37fd85c95ca0afb2369198a48ffa910464d41a85714c6a17e304dfccf2457d02e9b76493a9e0d47c4f0622087739cc303e10cfd18f33132d72b40f0d505b32b695329bd81cc66ade9e7ab69110ffc598cb2e97208904add32aa99b9810089fb6ab75112743275f317fb3942938f60cd52b5e9f6081363e0c4039e6893a7c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he78804b94ddb20fc2079e4ca35a1ccde6c28c9af213c2da06f81a56f7b4c158118572477b57f5c70bb987aae5bfd29aed019e7f2fbf84f0570c42b1abd36a4956cc6b5a0492b999ed5b61a8cf9fb1e4e5f277944b62d2fd1f77da61c3989987188d0269ed64f21aca11154b6442cb15ebe77174af0b1555f8f79d371791fd683;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4afb9dabf3b198d12798f1059f9e9adba2333093197fed52192110f6e69b3569c6304ac1fa5f38ffce212274e9d983fb6ef70f3bb1abf7ca9adb91434eaa47a725be238460ceaee801abb4f31731bc6abdd8e4fc86b1fa6f228cb42bd7c61699b67da96827442cb3f5af9bf9cb8a39606f77ce58c5ab39d19419f02643d30296;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c3b02b3e9ed9f05a93e373b7ed0feb27147f08feb2f426134bff95a48816ebb386416e92c37c72da1716ccf1b0016d0d9ce2866a3a861ebd838c403a1074a35ebb38bf019f1a0965d8c1ad085e54c665619004656c5e7fce95e5419c7e0e44191f28976891df2b5b7a8504d282b0a09f11aa71f1d1e014c2a13495f9b677f0f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1196c57c6af09cbe300f3bd5c934ecb21b824d22c7150af07695dc14be2f8808a7c30ea67e3364a92466ed2f75c6248d3dbeae3fab7ac307b2574eee68876fe7a7622db4ac96a5ce393d5a2251cfe4efc12116441d3a8b7c8c8d771c7e5cc7f09b83519e7815cde9de9c3d79f5131dacc2cd42768334ca2540fe84abe202394b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha225b38c89316eb869153d244986bc2ec86ead845d41aed0c61af22d36dca710f0a58d68059ce2522680e5bb35f841adc5c7ee0c9711064e4016e0d1f55c194ac26a906765acc7e2a2241c3b7bb98d1e8eaa9a4d336b347a0471d3504e11af26d38e55256098f41e70c0c3e09504be0454bbec64c9617cd28c3d08846278981f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h21a40007f45dd805ad87be8209a8eef7f776fdb8e25e73600dcbd3a9f9e0ba0c718b257f0df3e378b7dd297d4094ba25dde5d00d3ce7a530ffbb163b0d723260485af730c0715bd14f11f1801cedeaba8a54d29166f33f6f3cb747686f5bcaaac7485e2f3122aadca54c2cb564c37aeb5d420370a2d69d90fac16e6c5d184889;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f5ab527839f079c4c10b871209c4a80d837602d733d8b5466711994452777598e0f1ec560fc6786f735f340a31a405ee68d66ba658ea4332ed8a1debddecd204f763835e1c40e8f9184f625bb28100f1556a7da870afacabf9b7523a0a478ccfd6e8c68e9023c6d255151a0e1fe6bd8c4f840d922c47e066311dc0c7b038f2e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee82e5510a5633fb8e255a3377ec5f45059e788049376079bd5a5d3318f5ee82e5885c7a2871322110db0260693db9e71c33b58667f2f18246fb4c94f1612b1cb51484835799f7d5c49a03e467ea265cf732a059ccbc999e1f713ffbbc4683e1bfed834ab3ba0b147c9513b5597f521be90e457b38fd3386c671347cf2b27ad6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5ab37bd04e0e04344b63f7cab44d8b65af8a7d4caddd8d808c773694948ef437492c505ec38b064f175743f537d60f5f7d5d8c3f52edd8a5fbd71c15dedf270e84b09e7308004665ceddd1f779f526bb01990a01431560f5efafe3040fc2f20f554acf6841f27af53f4acfba467ba97f824c82e3ba4ac62034dfa7711fbeceb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ae4cc160e82a002072ea9b1b2cda7d68ad7ecb658351993d08f16b123f8e02a656890135d397b01a03cb7d2f338f10baec8a6a519a2bb36b99f55e9ee99d4bad2efd766339652051ba68f6d8fb0c36747b1ddb6e10dfbff57c9ab8e2a40b5ad2d28238b3b9dcab8ed039be71fef382af32df32d9287cd2a0a01219c30eb101e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee2527c95f79984b8bad9223a6390f0eb87705e58358deb06e1e96d8fcbb6a973dffc7ff601fa1fbed735184a1874a4eaedfced42d22fe9dbd7a6178855f3cf5eeb06ab0f6d8dede2dcdb44ac2314999334de73a738c0387c135796d76347bddf511f34c28438d077e158b8cb35c931517288c1498d08a3860a783fa81ed86f7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75ebe8ba6003393e84beb237bf772f44717baf66888a1a793156d4dea017bfc2138077ca9e4e52be837f491ed98c5f28725b476bfab37d3e6c9a19ae64ffd7f31c05cedf812d52b8499cebb9a2e3d26a5d75e0f3752e3aad50fd40148436f5a599373caf5c81ab4e38485430808e87782123d9375f40ebca1e86d6aad7dd95ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8660c0ca4f1f96f3c5895552041f0b0f68476b66c7ac6984550692c1c3a9d9e447765b2cae3b61cb9ad45b4a954ce76fa043332b2f9caf408ed0046007d894bbd7c63e301cbff7ffc6966e2a47cd0d9002a267ae82140b85a84dc92f071eb2d29324ef7f21b0ed608afe96fecf998887cb93926c6f7080ed1ccb3019ea31236;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98239257f63dbc03f75d650b407ba2b3e736c6abb11a089ac9c9c9964328e4cde9ced637803c87b592e9f159f68c101b7d18ce873d5bfed54ec32ab35cdb2d9a62f8dac9ef76419b727cb72a4949fea1768b5ee90084dd31c7c6074b1d6e71c711fd9b5f743a9c39fade821eb89f6ccee2a175b38139938219ac051b2561c563;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h110daad5996df71cde7e028fec1b6381eed5f67080fe39629ec0ac5a376b8cacdc54498c8ecd2d0fb4480cd51864c0a1a244f373a28d458dc822f2024644c70955a4f4a20c09d67ba495eafea86a2992581f896441c679e595cddc75f453994f5edc6e58c068b0ae2da110debde6c993cb051af646dfd31f4c24b7efa0faeac1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc20aaf5c11bf26232bdd4687cd3040f006ca58b06db4a129adb386cd1a4f60edf68b849577af4c393383fd7eb732e698f275321ed9328af2ce59089a5e0e4c6141880c28f6d45a2bf783a74b064cf811402241a18876eaa3f9652417ddbcad0c537c330b9db661922763709cfa6c1ce2ed8eb5ab486c012043b1846f203f93b6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ae3c1ca4bc2d80aac2538e98cc5ee4116403502a24910acca47be9a12ef1bb094a3e5768b28d3440a8132c6b470eadd4d4b8d50316166026c63e8d9663e33fc852b9f167f571dea7263b711a87cfa8bec01f38e76f6c1951959ce0992b6a33e1bc99198f4a0abcc422fd2619dfc1250401366eccb0b3a152042b35bb6b63e09;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3873cd545244f5f007ffd5dc8f5f66aa3fe49f6dec1f91d0a3bdcddcaa414e6494c449adfa18c529a0126d07430bafb21b8587cd099450cf6b6034675d62cd418feead425d11ab187b81ed30271417c449b999e88ad1a229aecc0ed04695434ab61d2aac73aab959dfc6967bed02f595dc811080ce17b1109e08a262a0f9f63;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5711720e94abd47d789b12e4a4e9d982e0f106538f3d1f7441b07b8717e2461febdccadce683bda7d1e3b771d8ad11f1466b42ae6a5583d5af0ecae417f4a99b832b87eb92fea07f3eb498f0c449d988218817f5ca60f71d65523d61b16259ed3e6121a4efa37bdc4cf90513a30ecf4485f0ad05141f50e1e474e1a1bb99cdf8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8587abe100efc3dba1d9b39758b55573bdaddfcda0a37d3d8137b857d58bd8fc006c302d87f2594cd82806f628fb9096cb8a48eb299f7194b5b0260a4a10910a27f7841705b35ab69161e5fd680ae84bfbc688fe5432a88c4220ed7bdcb812621c2db0ef45912a6e8670fe1fa63b9d4c259ba8f6ea31490a97b4e0c8ba397ec9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe6fa6ee5c912d636dd88ed6458d53d3df4a6b31b1084f89af445ffff37310d3dc75e829921f73d6a0c3013f66bfcf9f8010627163a15df60b9d3c3834cad6ada64a4170bc3ff042aa80507e5859da3523fa579424b311501911b20970fe4c21d71d78e2d6929413afcf990e64e456cd937462a9ff973e495208c5b924cfebe9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b4079015640e2bbf851dff653956d1410bc59dd305bb47fe67e8d5f1f34ee57f593aeca692d7fe19ee7d3eb606932fea49b954a9bf7317d89f267c154f8997261804b2256fafb9cc04742c73b5e1cb255692ffb34c0978b856486620338bb5f3f4712d057bcd32aceb176fdd4414a5e265958061d53938b255fe0bcfabfb254;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h198a839d8969309677aad4f2b93319859bbfe490d8019d85a9f2ab3159d215300d4ba1b288c47e945a6fd51387578492ad8b522e4cdd1778a835d5807497dc878b579b799d1734924c2126dd047150b4d8ff81c45a27fe1d062158215c6cf53cf551e0520dcb63b7da60a47f920ca2aafc16b548b37d9394109a0eb91af21fa7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he12b3663b466b584d6707a4f506a987b9d2aad838abf0f11c152943e5754e474edfc455bb25cca26610e5394ce611937ef81ad15c16b5f0fd6d583da07677cd2f198f0028ec68c1d71654100abe517353425743f802fef448231b26498ab169a63190869f15e688a9c764af16b76e8b02f0c0b629422e814c48256e67b2f4517;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb4b3bd9ad125d8e8cd920dbf5f66ee55f2f48c9bb37f9bb03fc7d8378d9e6566405213c8930c83f1a847e3b092e147acb6307a98c727a36d159352e06c83fb549d1665ec35751be6179c2789d451d7855ce6c628b4db5a4f8650f8abdff82f0e41dca2541ad144f5ef3ff1e10caa3828e6f909caa7eeeae3349584b276c41047;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h834bdd147be64439a62feb1f73b3b4a9047fed5cdc9fa816ee34adb0e9e8202593aa28d6767377cd2925922667807fb6cc43fb8be44e6d0ac5bb24aa40b51f80b5671172aee9f33d15abe9c94ee950c4edde75ff5aa9a169157883b755e4a51336d572466ddb60086dc664f851eb9a880c0180c7de41b6cd10395aefa999d13b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6193e19f4a5651c8eba05c19bba6cb3d8bc784d5936df8b532cf9e4520e7c3a6a6d00fa36c14e1be2d37250a454e6d7605702bcea1b4e11c328097202aa53cb29b8e3595304821c9670d453a4b917cedcf040c88121cd85eb6f8581b23d239ba95844c1e43ff4bc68425bc02e30c4e7da24d118a58750b8ac179ff305fe58123;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e4ed01f11a9d4e3ffaa9e2455ca7d23be6fe966f03d7f1fbf9c4b334e7d019261d3e3e0006e4d698d9e0c724b9ea25a6461eba1a58270c92650f9795389385f1b62d02983a5c20e5e03dbe33c3c9e3b546190782da26f3cb1b5ab90b717a73819b44c5bb4f549281b9507199bec9dc5ca01725f9850ce810e115e5b683c6ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3cbf2726fcb7e19d9bbc86901a2e365ffd54314820c9c1ccf6dfb0b94b91711b4b8dbce2e1639fdac3462127f7323ede4d1f14ebd9a6480ea3380e30f1371da03f006e7b2a815ce66ae50d70779b21c86235c4b36162db58cc60d16b0819ad93bdfd9e21b58664bc06cf65cfc28381a434299162e9c29730fc5bdf60dd2b9b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h232ea18c9b006325f74b9722410f36520db4afd7ed52421c75af94f7b49cadd26c32408215f02cceef57ee30d53d6b76164b705321bfc2b5e3e9fc0559d167f968b1dbad508bb1b928199b96b8c24d99704e91bf8dc69f2eb7aedfa4c5f25df581bc4dfafe02a1eb137dc3831306078ab013e19fc8c254a022c0b09e78cb3f5f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ac5122ae50bb80d3aec755de0395abeac2a951d4e35a615f78cfb546273a1bccd3a0df2494165613a3f8a02d6afa663c76c55ca84e0bc42aa6d3898e86ab45507a625f9086cc132eaf7b24ebd7a14cece3c8213cc53353d665ed3091afbad75e309da83a9cb4bf888807b2f19773f538db0f45f4e34efc4b8a18ca567d721b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e2d7abcae92b42d309bce7a89f383b2d70b954b56dfb0e7860a8f0741b46baaf32c8aa3b5d4e3c16259dd9b549477a6de1ab32addcd47c51075a93b9d6567367b10628d2821af1247b84855673083ebdb304032ed727b7866ee654d35b65269d2ea559661cb351e68554c8818d45ec5a12f794a1e83967342741e61977517a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51697107052f07851499b0da2337ac133dfd92861f5f8dc755f58fd38a00811bf89794665e459bdeefa50156aa52661bb4c02c286dddfd723f1eca8164391c88d06537be004034a1112fc60ae4bfc5ea895210aef99a3b9f403046fea1816158decc9ed715a63e29d44d0bd80daf24049ea67ef878f0a2ad1734b838ac73b92;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he47eac3a3897728b40a38e8cefb506df622e648810579289c1bc752587c5db9b3b9611afc30db502da725449ac473ea43e94d2cd3f8d167216c66ad8b4ff5e3d2c76f0930893e2a7fc8d26f0472e13375c683c1b8b16ac8fcd6308a91251cfe101a729be45fe89ce1f356a2d3fb53c9658127771b79457ae9c6a8699bdac3cf0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d435dd17235dd2aaa56c26714eb03091f21d61d1674abe37c7d3959a49f0adebf4d852135cf0aa5531a4e7a832f8442a73d80c407504eec92d416e88ed668002651a285fb9303af5bc27dc167095d500bc0d9ac9899c409eee49ea5b704ceb13b877fd24b2863c9940a2c6f1fe100260158dbaf51afd95483c0ef31708acad0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hebc1becc0ee6df799f68906206a80ee3b04b15951713465e80eb67e4a772eaa410ede406fddf44c0b2bc0b240a13c9c2aa52241039e26cf92714fb73f9e39fdcfd5c6dab9f127f9b6bcf3f8a4fba0ca6a1bbf92ab80d0f859345b6cf27d4523948ec23faed19d1225f52c9f29aed46cda5d8a26880310fe00e7bc1c1d53fc9a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he96ace5979daae1a07447049ab0086f116e910aaa9d5b17840ccf474c6c3ba351e33c8d9644cf86b4d387410e1d0880986878229f414556706eecb89b59bd36137a17195e08427f85d72d91c523265ded8f50941d4b2db47753366e67d00a31c2ba252cbbcf0ab16120dcffd622a46421e47931178ea19c82615577dbd01420c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97033abbe3ac026baeeaa99840a05a08b0ff4a8e7a9cce36f6b2cc5504f544671cf8febbcf86c4753c03a537b5102208bacfb93d350ab43137a40eac6b3f8c31794c6873c95faaca8ba9d8c62af354b199ef0233e56d8035bf059de64ecdb22c5fb7b2426d8956dadcf987e49d0ecc0a50101cb850f8139a214f07eb0c45e261;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6f9800748facec24efc18a3605aa862817dd837de09634079afa66dd41c6ca9e5257d3d2671946d7c47210b330012f505e12e04032a44f6f1728cc50cc5980c3819f927fd2ebe687783d27f0024b348987a0e1c14a42482ec58807002ab1d974456e4fd2b76865e8f82da08840919ccc4689129f8bc87929f2ea6e35adf6ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3f565b5cd20628e838092f69b215344bcf0e91c6ff380de5e1c8acc9c609effc21b8d36c56979728eaa00184468b805bdd28cff8dc24fdde32c016cf3ff96c59bcb470c1dfe1f261265f4fa7b9433681a01def548e08c8aa0e17dff580b758923dbbb86b33d3761389c2c295bbb9479c3d4fda62e508be746260e329e52d7ba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53201c7a09cf82ca3750dff888ee7bb35973355d936bdc0f38fa21988780fbb5df7d4c55b5aefcf6c9f4f8dc78836a7ba17ca95f3273b2df23802b0cdb7f4dc4413e0781ee743cacfe532a5d4023d2a88d4a262d86e5d785e89546d7b2eb52b733deec2c67528af89721b2c8b6b5639eff438db09076b2bb1a025978bf3e5b37;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha00e090af612b609f8907895ea137d7ba7474c0d14b85bd6daf8fdce2b06caed1614e233a87f8fb6592f1338f7372f985a3fb27576ef858960894f81625abd802c95089879a800cb30e977af5f2ec0ebafb2345aef8242cfb6dea510d8ed39ffb81d7224b1e9b6c50a2e9b049f105dc76b3444d39907daea603a392c7f66574f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h363d482536ffec86af412553de70fc5d6f7e994fff8c6c2603c98ee37e79b1084922ce589400f810de801cb37b72d0174a363cc705f3a9dd06a98755b6d0b5958fbd60e58cc6ccea6d1f5591b4aea853f3d08dda2b06c3e1545bd3245e41a2611320302e14f12d614b13a6ca239492d099ce4445b3ed4b8379627216d6ba95bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c3bdb7ad78c548e26bf04a6fe25a259ebbab2375ed96e6f6b0e28638866aabb64b2c964dca352fc8a2e3a2e075e2d5febc43387e338cd3d064da5428c5fcc5c7dc518cfd4b0ba013afbc60fa8140c44eb35245113a3cb35a7dde59433a28ab366bc7478f4f1ff8a0ad57e5dde4c134d1ffa5821d4e24a3f0cc0df73bde675b3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7aa4d28d7f4a79fd8389bd11d0fa267f677c652e02385f18a526c604533b09de02771592d319f9160371317d139cd7f281a4c0e417f0a419a0a14f8f097cb91d8c21d77c900ac7aafd4adb248aa4a87481fe390c95cfc685f23235ee94ea3fc2da2597a073072c740f1495403573e9e62cc637fb7b0741cfa01456d4f905833;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70101e26deec9f90905a93abf9e77448c6d0229e34899c584986d918c725f95757acc74176a25d8c67177b7b6398e0918b720fc5277e93deee4d9e58e29b27dec8706932c50b8841fa03a1424b94257551d13e6f21fed98c893dc2709ebde1c12375c1637e222b9eaa25304db563a90eeeb5970274651b385452c6ef10a4c3f7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha025045a69e223aa924707815f12750d8ba231ba86369be0da0b83a1d1c64ff8ad2e6380f0edec9c1ae683830e71ff98c0f9b0f9f8a61cfaad9a0a3912768525732d56f71f8a5929363a6f7fef735b705ec5a9c22528f098fb4ab712bdb48a663ebbff6f11d4bbd8b77df9cf054d1af303d2c6c19c728416a89901c3ac976b36;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h433e61235a958152cf185ee8738fa49fcde4cb51599504384a8332d9b0fdec6bdb55a953e0eda648d1768c5e391d6440b7b30d7fe6b1f8e5e4a37106fe054ad5ca61d999eb054196d71eb11ff495290d7a5c6631d4ee07ef903787ad6bf64d97ab92ccd1e6874475d30773fa705be8f4e7e5148dee871222efd9a7f97ed2758f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6db7a1327fc9ca10e09ef8c41400cbb622633aa98dd52bab8342421d0349e5f95f43d81ce8db012866b7215c2d3fe0d8bd9705abe20913328f9f710d36a536e86b4d4ad20e17e2ceedf8e6d70d238c925a1db24099778ab6da41670527fa6ff57fa07e5133e17c944a587c37c15d50c82ca8461bf930f26b2afea31d8d0b10fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cc7586674ecaa634b8fd4a8bc30b36ec80cfa14721772569ffa46397dbb2b17b4310af63b61fdd524922395ef06aaa11acf0afe1b710a6ebd8ce5991008aeb0f8b7c6513225e9cb7de2730128b4f801985e56a7a21fb9649edf760a5b3e03a54a796504ec85be931b00373b63b7977dfcd1070f930244b253cc6b4e7c61eb17;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2bf2198a57bbae46196b38e84ecf1cf1c96ea1509caffa38006375f4d58a6530d60fb7939c13b8af2c028072488e6638edf4103f57b6405a052323b79928dd95c9ec7bdc68ce74163e34709b9b67b3ed803496bfad3cc81609541fda33935128c6374d92f4852bf94c4edb3f8e382603a4709d4773b90fa62c810372ec4db48f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15d6e5d28b536b2a6ca7080810d77181db46cd0cc150eee3785f8a594c9605fac2e0d29b06937708f0130cd71d4f2d9dbec93545a170d116fe132af299812049bc517cecfb2a412e8c59da439031ccbe34e37569116ccb5683432884c753ca8bb5f81d10f6b2f4fee9437ffcb4bea5eb432271db7a12c7bdc3fd5cc364cc224e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdeb2fa62495efe727c1bfa3bc0d33e290b744f8116afc5899615eae91d2eac059d5ec2f7ae171f7fd0acefed77b274579860595b5fcb7a11f6b8e20829c1641585a724b84d74be74809a89744ab2057c47cd04d7ba4e4bf9a86791a92593b6a2a9054db43e93efdde09c127537242152d68506f5b38b863ead93edf9c7ca65b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69b6052ef1009065176b39f9353403fd2d1d81ac2c2b7839d90510ddde535a38082801d14ea97aa913ca2039f1f3a02f1b9c91d32044f8efebed7c4d77c4ec5a0f574ac584b28244f97cf0e4d2dd7dbf3ee3ebd349cb5b2d024c1eafa714c84da0c4294b51a77bc12ffb28bc9c24d770c1f64bfe021b4fc0b06b46d229ddbe79;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h375c10a2980553c65bdc7c0a60a6b240bc757d5de78782155a23cc734254a8b8712fd68bfe79c72fecdc0bd806bd6955c397edd1ca49d91fa24461f56f1b54c276d58e488dd8103f569fe66a1a2f7ca071e87a845f3bdee3fde9afdfe7ab13e795d013049f44e37a6fb0c25b9e9a62f815e39bfb7b90222400a4b351f01b2110;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6da862afe02e74dcc20a3b6e792c2c8057f0e2f1a338f7854cb7666a8b4c97f123064fabd2d8273f6465bf909defe3f3b4f4acb5d589c164e13836af58e05eb41eefb078e96478adc1cb80170188183c7a15af42d6c1955010abebf310e0ec8f07595f99437495b01ec866549cb8573298f0ad4587cffda18cdbb1239f41226c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h69e01aed37598e06287b9e85c9e6f2f417e2397d840f533dab2ea082a4c224d1aebd900415c15bdfd49fd1cb78785ab793ca015b83e938f015acba9a17cca948703483c231f936d6b1683e99701f7e87fae3ae114019a74fb70e9fe51b11e7a1bdf528ccd21dd748ba44e0756145659a4c1f7820a4d61c442136bc74b0c33ee5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha302c3c8e7c2c2769a682c78438938bf1a9af10ab0a4127daaf46e2f7e7b5bf566b8261d5b29015fb382ff13f697ca5ce19d78130403b00ccca04292752ce45a10a437faae7e22b9585d141d8e8c3fe8fbf1ffac0dc6f5357992f64bae9ad1c3c0a417e146b29646e1ce1e8c7f21ed857228616cb3d9372113e518ab9a60b627;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h171300322b42dd2572ef6e8074f0f54228ddc405796085c438e790bfd9d3bcf7feb297f2bc367d09aad4a3063a4324e613da9b602c13df55a6251f6233703109e791aa0dd87619d9a89c1f04d2bc133796e1f46eb15b09e0fc105d3bb5f077226d752769d1a833154391b06db9c9fe5e021782d1780d1e9317f44d8a2ab783cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h280be74a22898a8c8f1b8206abed96b53803f6b7b569d45939de630ba081cdca87bfffa79f8972e0f92f88fa3f55865e49a5900b56845474651d73be1df30870f244f83899a7b574b24caecd4cb4a6c7ce6ae94aab17a32adc11282381016acd5fcc04a40aec72fe3762ad06638a2fb33985cbe15b9df9af3d5c03a76c8d28b9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3ced75dad346e5326c46d3ca54a7308f8d689ff9d7acf83bac1ed94fc0e6b4248a1cf3cceabd1177cf3b52d5a8a78a413dbdc5d15861472c17ca1661f07b32f4ab9c8efdf72dba4f5354af746f95a6f1392b0f7f574edf61b7f53f1499c95676d353c1f9eac6871a411b6f32d46afa926e42bf527ecf5c7dc89220697d767462;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h59d09b9d9f8cf5731e17eb92576d09c976028fa95532e830a1ebea2261498f44cd58c31de127c15ab5fe23044b9cfd92facfb5d6479f90a48db54230e4c59f1aa14eacab90eb2010c78ed5c124dee367d77911ff7c5685bc1daceea886c870dc16f3159919a28ba148300f35801caf078975b87e4d95bcf4e8c88e84812b862e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b68beb2fc132b95cae1df24866be9a92bb9e6af113ad9bf54db30b510ae5b8317c805b34040f3ef97ae8af0e3589d8f1a003596a4b7c6a58d0db04781daa4b74d587acab2dc7445f03651980d8353a34a5d634629c79924fbeaee69dbe4708c0e7af9bb3a7ecdf94246496fb6b5a65b7d1e7e961249f50c479e7d4f5981d4e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b16797fb97c004075c92bc06d191ae3d39e2886baecc78e73fb3a6eeaa87088588ed44a5c2ef26a9224161d2c5254910dbb271fe7982a6004de1b223b65acab2fdfdeacf6560580dfbe5fd1acf60ea3a5487cc07c42f59ece4c8c979dbd85ef18ef35d62d6d2d23d9f8eec6e7a78f322fc09eebf57c165ced37be3760030c60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h89046ba0222fef2a646f1067f897ff64f34c4040eadc96c3cc1edadab77118f60ce13cf5078a24ebf957ec43cbaf05d2ff3e42291c550ac942949ba707919b41ebe2bd7c49ce5243d33bcd9f8f7ead24339cff14fee52d37a866f4f975f923e5236f9cf3c088f3948a0cb9341136de6c27542b0ba1bae264270c8766e8c71ea4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4070b23f958b9a36119226c3062aca0a03a7bc47175f65c326ba845acca122cf675f6d310e423e28f0509d81137293dfacb4b41858142d1f268f4608263b79f7d126a624e5ad2beb3e825aefc275c2809c8ac107aa3ad44b4189cb185d898944ffb4fe423ff6b5e06ddce6a4c984211c887214c649dc8e4f72f6c0891f02e469;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4878f9006343702a480f02b6f05bd0888540cd8188cb20eb899a5bb7d7a2dab37ab234aead0495dd0aa9825345b743090f18f127c7e2f51d1d99d4741d5cf85a26a7bc906cef2634910a37008dc9d36bb248fd9b7bd6294e1293e865aa04eab9f303f7a0391b8058812bbad70b9b503663671f271c29d2a9e1899426b7162569;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6f87c1184acfb95cdb3e1f54b3b9657221e6a4b276ccd583576932db38ea0c727fe1a62dedab5c1d41e3bc3574b10364afe3968b736e34a5880fe090197f3eeab98544c2c0e5899610c31d87b08eef97d0e84da1598bf4c102ebd575b7d13be47c01c749b6aed33b8b2b4db4c0d665e4a347c13db7ec7f7727df059ea8c47b04;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h308d1909e2ed6e248e7cf11a680b4b8335d777a1782e4f5c4561c5889ca29d371d8607d2cd8fac956a1ab07ba47c1770702f710bcdc4747b901f068f489ab028d8d6b70c216343c194c7dcbb617b2c755dcb6b476cb5446cff3781a3063b6f58193d5f888f0a9cea9cf6f5384f850f630d3dba37f1355fc86d44e4c3d7440dd7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c44b1017bfa6761c6a89a06c0fab5f21c24cf01cc25c192143e0282e8cc95009b1acc1bc0eb020283968d3a021dacc10481799aeeabcba3a1e27b28fe6ae85e363cf9df03b3bf94db9f3d9ed64f3ac3c35bb73b6ff52d8f8992dd536f663b81095cfe31fa933606bb0f74c55ee3985fa0150806c06a8e46f5e5320aed6d46a1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6089f6dd9ba0e63f0166b3befb9958afeada49ea7ee39f9085558c32a5c7d9820af01aaf580f92def065faf607f794671b8de91545b7f4b00b7b2a9a1f7c302ba19689df6341bc211c576a92fb5d39bfe4c12691f0f20451fa8a4b0eecc0e93023f95ac1c107153f4d6a33de9439b2de138c09e86f4323d85d7211e4febfd00;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h135750acaf79d5c92482142c7b6331ec6e180d72e8be2af66707561c611de8f0bba5c3d50a7de9005b8b7f11b5ccd0a4a56ef6793ee994f4091e5f52a377d90e2990cca74e7c59a5a0fb81af6fa650ba941058affc3a43871cd1a53c2535b19743990f6e5e842e8eff7389fe6cd7e5b99d42743214b728ad2075efdff421c629;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee8787f7799798e92780cc61c5c474bc77df96a26a5dd720c265eb0f91943ca070505a015524a96904d1d777e816e521f25676abbf4a2e54de2ea9a1e6d46d126c4ccf10a19ea5a35c68c78daf563e57d9cb7c79369a6b6d9e6697cd0461d65f1db898ec2396a303219151178f26c9e1ed58af23f85e3a0824dd614e46beadd9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'habec68d6ebb1c76975d9ade0ed7f9228b6fa302be5d286b209c0047c419a0be2ebe1a775158001ea281b8ce222c7a8ec973d7ccb57a305bcdcd0ac5a335f0d6712763cfb34dc52ab06934d8e0848ee242c8bebd8c2f3ea8b47792506494755c248933aaeed7cc2ebd0fc8e4f68f935f20907d180105870d574413fbd1154d3e7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc27149efe6f7ae28bc6256325ce090ba90b91bf14a9f420777b90f21394d5de9d3ca31654c27b8543a7421f4c9f16a7d1a651d5cfe840579a865eed286de5281dfc9c30d2bd985c8e1c83cc1428403f31f7e091b7c0564158b981cf7985d9f43c46fa958b6d56d99ef4369eb559533b134ac81d30442f617990dbbf054aea366;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h104e6cc941415c9cecb1340aad9fb9b09fad3fd56560c204f204a84b666445de3883ff1edb8d99f3cbd918aba0b05b3238367e34d11a6343bd8e23e41dfea675215774f9a489fb055e5a4c529e60d45595257a6587a320f4aeefed42fa5c222227d673b25399f3d1f2179810aeedd5dede257955d134c50fc1c3efe0ae81fe6c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc337294d5334574f90267a7eba623d841b7b07e6bf6f0c2143c46c4722d0624e86415ae4ec103e9bd9ee26898a65393b51fb06a6f3388ff11f16f56ba274fb28e8996efa5d2075db7ad6cb321a7b55f3eeed1dc3ffebc264f291204906649d1741f82d62034f11a3b34f963c4244ac45d9824f311b3339492d0ee8bcdf1a101;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbcc5d7430a7034ea7b04b2ae10fe3745e654721ea90db2a9445a122f89aa07ab1919c37c8f07cf950cc211909a7389e19221600dda8744f1161014b4ce5b0b4d963976a502681dd0f3b5415fc8e3d82e2a185135b6057d8348540408affabf1cbdae1fde790382bbe17352263dbfdb1296e99a3c165dd85907290c03298500ff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h539c109b20bc3fe068ac9aae8433fb8fb2b489a8d4871bc43ef61d085f4a1c75e9b30ec6e76dd707b5a57a045215fe94d23b7ae9aeca54eee0c0de9649c6d1ae06fdcccfb29a1954fd8ce978aa276b65e0d09eb518b30ac1253fc4e6aebf245367c2c54a22d4f6f5ea7a1c86b6a586940e6aec134b43cba5cf06798459716d2a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h159da55f9a2f415a09e2c8dbac99083990a2939f59b1388b958c82b0cf5fe03cb17a61306513628a67af7ad087b3199b0b886e925c4ed7c9924e8dbf158aa15b132575cd354d647f4bc39e430101dda36ab7783ae47b8ff43168f2224ebd35ea275b348df04b599d09d1efe3642afcb1a19334ebb2e7849f176723dfe793454f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h58ab69160c05cccaa96bdab9c3dae3fe3d3e0a26289e282ab84ebbe8e9b6ba5b99bad8a6cbbe3c98ea62265f09e7e179a486c0a4b92df303c9009aa863d96e349e3b4f5977409de22c211e465ef8c051a466fdd2a5cf8173c5f77502e7edd1b1f60ba5e73d8c00f8d2578a03ce7e866adc0996dee5e5ecdbe3065ff14237cc71;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbaf5213aa1df39ab51adf4592c91293c76fb35bfd3d6926551698062fd17b0415c5573b85d26c4b63d2d4e1b415acbbfa76d298935d0a715d74cb3783dfdfde406adad7ad0ce62b94e9840348e5359856d691babb86820a675da5576a0e745241059ba58a63f1d9fbcbd0ee31a70909d0e341e864ed10838e3aa30feefd0cd96;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2da85aece469b7bcbcac52e23d05f3dcbda6214f65da279198728e14105ffc5cdea12c15d7797d3abe789d6cbbd8089186ffb714efc4726afd24e1a9c322b0bb48d1fa61d0a2c8b400244b041fb275028118c4d4d55a0842ce701ad0f6ff630114bfa6dd2d5525acabaaf3b2ceea8145b14d0330fa816dbc9d724f76ec8f9250;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a2fa4ee5130651ab7e2ee7cad85738fe7c65377556916ee80a04b9f87038c06266f1598b0e66685c2e27e295c40574af0b041a7392cccb7e04394333cd24bc8787f47b357bdceec0d5b6857918585aa61ec8582a4d2c9feea6ac08671b328edcbf567b162a547db237084f9975ad34aaaa548092a6f7257a8fc7394b8cd25ca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba0fd3000cf63a8c44e98369f1e332c79e6b0cab77b6b66bb4509344c5d5d8a919d9fdf4d9cfe0c354b7088b552ddcacc5b061f6cb9d9720dc35ecb3d10d4bb8bd34f3b1a79c46328b3c1ca9bdf798e883f91b3284d69af2ab9e63b98bc99505f16fe02efe095409c85d583e9b95185ddc090f5436a74db9623c9eb7cbb50d89;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7241c7dc34a239b6c608fb433bdbca7277b7edb9fa313ec6da0784f605812a917c391eb80b962f42b20e28736a08b8dab2f2707e4bbb5ce283429c63599db98ae2ecf66511f217826e6e30406c062cf43873b3c506c69a01ca787f44aba3a8eb2ba3ec338d71c20db36b59e1a43a81af3ab10ff2baf64b05e948045e80303388;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h48e0997a08bb12be65aebb249ce88e42023352503cd2ad900d1baf35efa1f372219607e61ab5f1ec5111122fb576c23b999f94791f457b0e043b6ecf9b5119393d99d1ef45f37ea80947eaea1911ca157ebc521f2ac38f961aefbfe3be0b7ec22b09236b6c80536b9a5df2c5ec967d558c876377be75771bd31f115fabb7de46;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b25091f6b55c8fe9249f7663fa24a6b8f09c5108e74b66f47a3ba5d1f8768a319fed0d8acedabd3c2c5d69d01277775b7decc73dccc0bdae65a37750759c84aa2b85b8b77f8795ed520719430ace114c9a6bd3a78e1d56a9c67acfd8f5c634736f5ed284deb811fd9ed3c834d0e3f1c8bae64ba2168a616ed21c1a80b06a86e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40be70621bc97777fc63228fcb59ee816277f663877e9c31e853fcb3a46a8c1c16c3e3c7315e78b649745ed497f9469d2422287606875b424c55d51c511965b1edfbb366e94112110ff151f7e21bb3cc11ee835fb42a24f01f84a56f97b73f3a4bc0cf8586f8be53f91acce35c8a35e5f0fa04a34225f50f950ef8fe6136664b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha13ad5eede1d4b62b32606786d12bb674adf59da45b82a4b0021e17c98a8cb12210ac6238e26a891b9ae09c0fcd2fd5497013ab80cf829cccee6f7030b037fe6c558db45362d04188647021b0376d1c79b81870585521cd4dea0afa4d701908a5589c092e940d99ae3d70681bb41c8e562d159d80c6f97cbf083e5e941ab0c9f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e60df9e7bf1cd8e6f07e6fbfbfb23744a72379a1e9def81a0c1dc701cf48dc0f92a33fc15d60705d937e2d5ae22079d5d64325d667145d2e4579dc4c273e36ac4b7eaf6a3401ca162eedc921c18efce2e150d45407bcd2b605fb303a1598b44789235a6b91ec9f2b21eeaa97ef0e3dad4371725d22decb8cb28fed6717840fd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he857984e78fd4e365f26c68ca45bd51bdbad2f6bfbf29b06ae0149937881c38d268d2ca1807c241492d1c94754fee98608043838bfd9a14e8acad7b6573e3d6eb8c6a93a4fd7d95e5e43b4815d54759e295c70c152280d90f5ee221da1aee171759c2b5c5a84afc19fdf1ee846bdd2dd128ac6b3a1e5578eaaeb02145bcc0a04;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h215ad0db3a4ea33bf7734630dfa455220492238b8fbd69186b0d837f81785b0a1d61ef5e26117274d8e5a432fad29d95f84fbc790a42958a8923b8ec8df6ad679ad33a2e788cb14d1bb2f692e204f7297dd449503c0fce8aa287b39c819da3f8697d2d5850b84abecc703ef4d98b3816742f7366b0294bbbcfb1225c29824b27;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha42aff548649f2f9e117f186f82bd44b824d9d929fb8361a0e244bdbf2c4372ed1a8cc6c3ab96ead2490c84668bbceef8f1bf53b760dc5fb9c35e303a1dfc394b70d5d56ed7f15541c1b5f1f5e63bcbd714c5f96e024940cab13a7344b277f65fa7a18a03d038475683cd2aea8f16febd8c87fce9b560e7fa0656e682c3559a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha030f087b9b73b3eed00b5330a9116308e0720f3210be7072936a7f7050fd0527235af4497b6420c84375db87f1eb630d97f20594277870b7059a6efd12b05a067aff17ef935845092df6e6234d10c3778bc66799f2f7d0036a5665683b1d6ce10bc90b6ad3908132af535f17f03246bd03f16062deefb347bd123ab00d379;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9bc0dcc7d3f0fc67eb64d1d4c20dda0dea70ac7472c030cdcb26e59191040efdc4e356c4c6b83ec88b278895f3d2856bea3bbce7b74561912706c939c0889a384a2ad476da7f9f4e07bb450b7c64544bd0cd8d5e7b4ba0a2fb05ceb14e9f897e00d9987ca5f218dfc8270e63883fd4371f0ed40082a9e32c706c6a72adbd7e06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc81fbf3e35bd7911247a3587871273661632c82dfaf1b91440c68371c5b03ba00010103a4827ef4da247b5578f6dbd138c76698452f43e3c82d4e7871b2e57e34038d6655e515a5527efcbebe660761524aff01c1673589d87292eda5e579f62ff12858271ef626c3d7199a57f0a3ee9a88eee3713c2cbde91a9ea4b3bcf121;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h11fe3d12a7162673253cf583c0780034d998240f3009583e59ab637c3b33d9cc96642e7cb307abdbe0aebf559a43ea5d348eeca15691c5acca609dec61ddea6a177f0d3d158af8d32e18ad00233c11503df33ab53f60940ba1c40e76f9c235f516195ee6c269a742e23decbf291b38f46b511d8ae7f90abb96c3f671f2dcf9d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6cfeb40a1052ab8d4e60c7bebe8afea19c8f85c59dfc48b7e5cce8ab876a5cd26e4492ef23c8bf029d6ef79073022459ca1700ae92deaef645c8c7175285296625df49373577c27330b82aae5b7458d18443121ffc05f23cb801e7d264e9c708e48fe6d03c23cc488cd3a24877ab23b03f5d66751c389ddfb20f7ef9764adc88;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haec472306a746f175b951732db6167806a5a12d96a6b4fca1dbea38b09beb4315d996f7ab66b608ef60d0429db62abbc5eab801a1cf9cbf42fa043c5ca9d47bb4213a15c91d809ffd1b946abb9af6edbe37bcff5147da10b6673c9d6cd4e8d556a5f82e17ce2e881c40a5f47a6231f86056d6e5cab7fde113f14ed74208d9651;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1063fd1a1171c8a471d71c7d291c6a32ab138f34daf6f5cd69e34ce3df899d2e7934b1c2879c4dfe2139cdd5287dbc0073e245b2a689e5963d336f40e6ce6a0c6bab30740b4f7c836aeef5e6578c898ff9945d557a580f9e7946148bb4c38ace907d1b59f5000d899d8f2fe9ddd38fa3632c28f28ceb2d6260c27d800ff7efae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6355d40357fae09ad3f17ef455bca8a7f6c256316992b3467662aeac7506aff9c340177b7c137f360cd2cd41dd531b165b8afb7fee490198fe0417b82f013cedca94e41ac637f8436e26e7abc8e82b6a5c12c8d32311600cd5c19519d5714f25c6fcfe1d2698063424dddd9336f581cd50936a55b5219471a8843f8f4a0a8d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h120225808659a9555f75250f29de4b914a19dbaedc75341c249194be6d234d8e882901c402e51e94e943dc7546738c239d7650e4fdea95c838ded13b905519195c03a0af85bb57e555bf45efb13c5a58d2c3bb68141bf3d22c7151c80b05969efb2f6114ea2d44c7dcb4b669182534ec7bce2c75e8d599a621ee6c81a9e22de3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2af4d666e3889c4f669533750bf9d7e50157d7bf0c7796097455de16ed2f9f9646780b0c5c92365f3f934140ffa7a40fa523ad2b7dd351b7b6412845bc0283d4a28443201140c8ba0a390bd359748dd8cee2e26bd2c76a35efdacdb26fd33cdd1af2be331eb7bd5b20bf14130b6693a7e61b9cc77be992c55e6a31409b3d30e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed7acb5575f369b76637085a85145d6bd574a664a6fec069fdc6a7ca44f0ac25a9bfc6d026851304a4b86d6664112d454848d43e3bfc1c6f9da7d99229abd9f354e6702a58462ea8ebfd17be1bef9df7cf2d6d52cf4a5a87d93ed990eda93412075534d92400a13ac4556cb9b57e604dcf4c52467562b96306adb6925450d807;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54135f0bbcd8d4b4c44e63933ae298fa460b20497f5d571cd8b21b33aaf1d0c522cc2a9ce1a77b0923ff9a1220fb3bbf5ff7c40407efda005ecfca911a0c09977be8a4dfb4b658c9dee2b169d3e54406eba93c050fd18c16a8ce2c4eee8699e09a2221278aae98a37ba8943269d4addd558037d93913b1f530d86ac12eba101a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf2095e812366159a6ff7546b69faa08dfea68556e15023379bb4dd4c661b51e899a80c71503a6f2034a78a837261b008711aac03f6e547ec57bef4a3abe69309366a55ea54da69426b5352670688c2748b01889124110978934fa81db292946abcb00c12c328a9ac46ed137413d5bc663408cd99513f3d256272d948cb733aa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4888af41958e95d25efe692e87a96a10927f1ca8e8176d68f5d3dd16c7d72bd1a2a18d1b146881d8bac0a79e6d78e151701c4c97c2afdc6f9ecd747b929d0556d6e759c7283ec4bc308b7309fe59760c760f538c6c2429489e6d734b1eb054f712ca8db78597c1c687c4a66d1a0f5b3b932155b14d032e5b94d6730bab48b49;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a96445257fc985f28f1ebff69c4d6a4a86be729aabc9378a47d0c1a85de1445366ba6840029779fbbd82f6b370a3276e5a53dc4302fb6c2612edf214ecedaa0fd810193e06f26fc44fd3c0076dc40e51eb8bca33f49681560f802f84faa50a73ab088ddd53fb365788bb436442e660a8801cbab198fb7ae970c501ee8afe681;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h48cbe956f7c14e5f7dadb59d57c267c93bcda05dfeef94142434aee662cef93a4a0e939f0a2f8a0c1bdefd28a772b938a9e4f243fd5d2653097e8952e32f019bdec3979c5a333a21aeb9a0d8c0489dcbec7ab9bec01ef5fc2e4bf00e2e1e5befdacf0a49b069652813e790de17be7340a3cfe189ca101df498b2497e005a0ddb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc8f7e8ecb3031b3af0c20376970f60f89169621dacf5f864642cabcc7bbb3292bea6b305e05afc82676ee803bbd2c234a585f1d8351cb9c12c550dad58df354ff7859b2c01c789b8d6fe2542809c529c22ec9563c3886ba2326b5afba01a95ddbe8df8ed1b6963b906ccfe7d9639778eca2566cb5429189526cde4420ac4a61e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb22ca75e652b4c759140567a15659893e747c727aa2138a1cc97cd264b1e128b7aec494626e62f0412e097fb7d90aacd73b6bfd0cf980948ef81c331790390b49440c1e4491bf3166c1071f0c4b07567e203186744adff86758d1e86d5a1c6b84b7ff932668da2d18dd833dcc07815bcadf1f507b84b515ac7124b3911ba5913;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffeebba91e8d0d623aec7537b97f47029fa2da898227495a33c26dc565a54b074e91c23bdaca5882b6ab269638e7d7547ee2ce59309dbee33298f0ab0a50a37a19d5818ab5221ddec12b51b603bf28195baf10f4cd4c5f54b3db2a1c78e5a4bf7d0c82761cd38dd5f1df44810f8e5f7075a93ba6aa26677769e87bd719f63b7c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hafa1a647983098106ef8efa45f6c586154df4fd5198e55e5779fc0a1b2a2d89fcd6a0f0840bc7f90778dd8b92b5a54352bdbb3efe581ebbadd461cacf2c3ae788fc62e8e9061b4b43f440192d6e7d403b04e79774a0457027663c08aada97e1010ca5c1e6f1a8d7c940f82b67e9f91c5b390257dd660c4e63f43d6ec3e31fe55;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe70ebc56ae61ddfdc38546b3b13c7e86d4bee57f873fc40a3657621d92a9ee1b5c90243af60eb763b8508b890dd26595fba52c0fa7807bbc1aefc8c501521db14ae3522971d52bd3a3aa569e29cf4b2c1090fd44cb95a5d8ab0dbcc6e92dbfeaf33af04031fa1ff4a074c1c538e923949daf3053b572d8ef7629908496aaa3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9ef43c598e89ba9eb7208d1efa50eaf1495dd187cfc9f5b471d56bf477b4da4e6bc9fc21af5c24bcd4497139b8b04a294b9b7672d65755ff288ff2f2accf1266fa91ca8b395f82d633f4ff0f17488f6dca1ab38e69152e8c37c585839f8b96dc556fdb29f3542abbadc3e4c703f61de52647962dfc3175ae3cd8d3e86469863;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35157765afa52a2d847b010d1370471908fdf854e7b60a56f44dc2a54dbe248e8a09d137db2fad08ac6af3a5c0ef27759522bd569011ae656632982af4a1ee64fac0afcdd168624a0e6969f194c7cbfa799e1b4c8e19f354c3462de6d20b9730c02068501076182e9f642e7c7d0762cf31a4504acc903d92c61c524f1b7f0d9d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha175f58caffa37db724ca8758ab3bc763cdada50a84631af90fd078ba98b41484a6bd57ffcd8b27fa429aea1b14cd6abe6689e9b6a1a6de85b18f1f66fd9a14a4ce564c1926606878802ba5da5cc85eee12b0965001347e427489400ed9bd6f427db164fa9fb165874c28e2f1e49d422f2239e248aa4b158876253162ce7f4e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfbb834200f721b436bae1080d27cd1fd7da64b6d7eb72d236832b1df3514ab6072d51e0db8fc15b3f13646289e6631b00c60e66261d3f7fc18d7fa2e215cfd63c472bc61187a2dbfb90ada01f360f39185bc08fd9e27f5da67f1c7f0f85f84d86e85a813cd431112b22e34075dc5ef35232d1b06e3df38a5c461354dc6e7f96b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe4a3a4e0597b1ee2dd76308b066fc2c518b302c0cf8129eaf09a98602cd0e205c1e46d0052350acdecaa103d872ebf20e8b953ae1efe2ca8554b20f90769f3c3c9c5dd971f0a75f189a2f1c908b440750ec33879a0a48e2a267a93a49b58ce5018a939e6841c28e5e14fd5ec1b8ce17be10dfea24a28407a4db95421473c753;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf427dc1bddbda1d0ab2d7277ba9da7f80efb10dca8d549854baf481c5f80cc607e1aa2388fb6a8be6dc280f9f2e61b0cc453027f05ff10ed7a23044f5e4923296e28e36e4f1c5bc66871d76220b7fb26ab757842796aba9e604a1fe909696c35ee1ff820043c6cb9a359df8dcbdbf3e70b1fb3d2e8e02cdf522660a10939c5bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb658e518f038e21fa0197c54fc7d9bdaee9b8465d26a27487b1cda080c072be8d70ed81acd2974eccce4134ee6b81f69b1d57c377a664e0d5f6af60447271413fed34e3dedae85dd2e7bb75911bf2d59a0e5f63e0151f2ecf9465c40d5401c37da7eba071bcbfd7f04a1c4ad2248f381140cf1ed39c94631daf01fccf54b3a8d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3957a7cca4e891bdb297cea7bec754297d2bbdb3740c1ca3245713dda18ce9f3bc8832e693b41e9dcae6b5fef79bd4024b9c9c755271f331dc2e21b55ee5f0bd38f20fdf3e9d4debd1452c22c7c8588258cbe66218656f4cf5155b79cc367f846155becb6eea74b63d42cf824a2662a4f8a9dcc7bf1f5e80db719b5933537a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3644c289a7752b4eb2969ac1b09c172ae453f0c1de26c823e074576f6b8a07db29c22840f25a8c85897117e3b50dc4d0718c7bdf13856b0b0ada1f05331bb9dbf0bf173198e16a6e8f427b1c8294c3eef965c69878ad7284d268f4fe02cb41914527e9935d0a1874f10caa92e7438235117d768dbfe3693a82d157aa9a00ea4c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1be8553b22cf4c840c57e54ba37645384215fc5da488b776ed106ef1a8484b5cc6b574348ac412e6816c6e055b0feb7b7cd44e538218db940d46604d9cf70d3364f07236d0bbf27f4c370ddf5519bea660097d7a98922b53e57963f73f31ad6e4444e96a76a2c5f6220f70223e1c70ea20d10ef2ad177fe619a089b2599a8708;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h23c5b1c937f53d3a1bc313b2855a0666341a43892d74aadc71016e26af778b470eb75cdc2a884ac32fdf89e7757357f876302f6fb904aa1dd1fbffe2e0343fb39d4acb964dc6a788039fc50a3e9f7d5dce1bf4b91eb4e0a402d16e25661910cd346da55fd84a5968f09c6fc73a437111fa6d0b410a25634a0841f7e9809470c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h282f4f21b03095a1030db7519ef838998a4b8dd373093afa287708b07b8a800459d0cf1dd3119e731c822f407ef5413404d3979e1998fe1dcb9366c49724c334c165cb2350b786b77185fdc8f27a3125b6e23358c8de8420b2ab2cdad92d32a51fed40264b7277d33b8b7894ef8d12d0c3b62552fd70c7fadc95ec667623792a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0434a98887cc2b33936e9d521330dfcc7147ff77a5c74d75d76879834db1c7ce51f7ed4c0762253f85609f7966192f5591332dbede437e9514dd7c89fa77b4ba44d2383027b4c6836821acf1c48abfb11fdde261ead887f8facbe8fd3a0f17c0fbc40509393659ad30db04d0b629b1b1c2ce576b31919b8c06124a2ac227216;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7fa30aab218530d19eb8b360f2671ce3b9d375dfc745885e1746299ed02023997c67a94e48fe8b010c906a822ed5a597657dd6d359436e49c63d48d3ff31e1cafeb5647a1674fadedda72ac95d7055a2b22a49c67b7ac80b527e4c46d1d5b2563eb81881707f3246c9e021cfda8ce28ab73ec629e03cada0c8306257f80a827f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef738635e1bfffc4db459efa05650dd0784f7935e59174dc7452c6bf11a796f4eb5ffd0dbfbddc35d058b5c34764df8c7fe3f73d8116b99ded7c7173c4a4efc5210fa25134ecb4a4b654410d1bfbce2300e1858535249688fecdbec9be1446c85aa9039b30f209eb50baa08146dd7fb236c595da3e5c8321eaab6f4dd6cda7fc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1049bd1c40eb83c15bf471392ed30275093bda5e83f305d0bdccb7c0bfb085beddcde1cf0dd6a8f4733c43c7c0ad6f588669ff1c791aa4e160ff076690feedbd679f7cf2b57dab09c5be4780f343c7a2d0caa7682d10245cfc733b8a13e228dbe70b52a2a4b2e9e2738da93dc3eee77bc0c0d26a30706e8028f34a8f09338de7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb6fb089b5355fde2ddd15b3ea8406ddfc6cbc18a8f21131afbdcd2781ee26aa6867139bfdad4369a08a3f419996e4f6f1c9519b4ef9f0b46045e450b6d6d51f15259e8b5d8d600847fdc8c522551b9157df9dddbf982b3bdef52ed0047d0a4384f7fa3084ce85ca071b1acb48d0c68ad12536e3f5d58195455fe2b22efc8443d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52c1c48965db3519c6ca0b9a0e6553727c068f6d7a7e5d498a9cabd34a754cf185eee22da9beda449d03ca4630a571f730b4c32a507812500c78fe4983c6ee23e393836408124cdab3c59e61b50e1ea91bff03726b30bfd13c9b3180f0103b5734a961515992cf07796cecd021c16c086b8abf59f01a5a8621330750f907585;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hac82c211c87969bd092c2a42e5532bb58f3e135284a7084e1b2c228d01438db7ab837e3ee3d23e508a13932486dacc8c8820b592d859ccdb259d03fd99a9b67094a4f74c4a23858bdd2c1244076f49ae06ed44dac8321b02d31ef684f87f9c13a86fc90ddd27269bc5a82dd33aff872b3bcb06709405d348a89b64ba326786c5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb2cdc9e9330b913d79f6c9ae32018b2ccb5e99c45579403069447f109bb93bc79876db2fae3c160d9d90d2ddefb02244e686eef94720f3d51de8c4d9f6e7b77059ea0af895a49a34f8d8f4f2f2531514784f1b01ca20a5cdbbb193534ffcc092ffcfced56f25e330e5b71cd8bd840bf53921ee704d4a2fa71885a3e0ef5f003;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d21df6e29ef58de75ca21be0caf24d2f6420f1a6fc370e61201d75f8422545aeeb1eb082745ab51d9e3d21ef461e1db435d6f90996f17044a53c85bc925d9f881c3365e9574cd93d91ef5ec633fe832487265d2eac59f6e3fcb0b98303b18b1e6d684365c2a1b78b037a185a73735e26b836c79ec2c33f3545421f183a8a889;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he23af1ba77024ece8ec54c3be602d40cfe492872faccfab69a5b4dfef2420987d5da249db3e5f002e54ca626b40f64532e065839e07fbaa1fadbaafdc9e2856f167ae837031cca712a57001c4fc9d59b1d8047a0d480e19036f70934be33206f751e6cd06f149daac7fcc5be3ea56302de7f11291579c1e616e1e6d255ab188;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h637e4072bd5fce8355f06f2754775b60afe8a6657059d63a91d2acbe2658fe4901a992a2128a1156747051382dc8a659e58b02afad483d69b50413d0b0873ae79c7b765fb7a8d2a0e222e2da66ccea485d80b2f39e798006826ae805fe6488137fc090beeb5efe0b0d970787d257c085ff5f70321b6a4471da676108e08fd1e4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4566bcfa3406059509c7a0421e582bcc5e304afea19b884fd44f95cd08d5750ab901e4f0996c71f10cdd4d6cf4e861bb17128acb24e0368229f17eb7ec1f0a5c204d27f3ab303d481a2ead1e3eefd008a2b1170ea88fb7b1340633fdd596781009691d8389ee7fb1f149985b5b95b6dd0af341d3660dc69b90d060e0d4889708;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19b0253921a8d3574193ac42b0e185db9d710968300abff1b4bdd0908088d21d1dc4ef8eb974dd1fbd93aadf081fff3037572eeed41687c66a7cb7111a9aabbd172c1d2803363f862c782a0fd434d0c4ba61caa099f0259aeaa3dd7aae4d7a31083de7bd837fe44e8e16c3da99c01aaa9ae2d0cadedf3e0f8276ae4b1b8f274f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10edcbfcf718afff5ff123d9211c1952abeb2eba8dbc7e6f13d23789a190bb0480b5883537d717bfaa9931ad6fa5fcc8c7da839830b3fe26aa8dc881f6bba73049d18cd488d848eaa087120b10e136aa065a01638b4a71a31957226df4f64db82bd8089ee7384a71886291fbba8f812b62a0cc5d1a821e680743d53056488f82;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h126e52ebd39b044965547d0882ee62496aed121477a4f5e597a081d49bb50271d10e371cd386cea68cc81ea22cb933a7c5c9e2fb473daa5f56368f8fc7c8e19935d9b5febf3d78a44ff98cf1ec1086efd48ebb7f1ad67ada9af4fde61a9607216d556940983ed0543525ac72356711db3f4b57e9f18c72d524cb642e40f21f8f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5dca0a84bc6cd81d97435e20e5705016c11d0c3ad8d3e4a281a64ca0ae9c3477c79b64a1698e1a05e9c92a1db35c21cb4dedca59f18a2df53f23c0ece9438327adab51c3ff81721ae27efb07b288c57f307661ffa92e22295f2367ee6e1d5f70b45953adb437d4779dd8fe9a5b828a990dcbc45cf6d22e39cb58122c45f89e89;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h556ff22c0e4528f68b4c0d3dff607ddcf0ec7cb519f785fd735261d18ea3857b7173a3229cab55795ff79e33f3bb538957f4a83fefc45c106dc646d4ff383e6a99394fa2cf47ccaffc1d4a57d72b13636ce8f06a0a6406960a4e7dc3068c84a3793e413b49e072e33e3535722de89e55ebd059fd31098d73bffad04aea94a0ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h529a3149375731ae205636e006840bffd4f306934940ca01b970f0f299e3f607a09b0fd7aa6d87e43fe2e96c1fb089b3dfe0ff8081650156d0039e39d4bdc6115925048d201978ad699b14685dfacc0555750d7cf5de2f6fe43a3c3090a0ebc50ab6433944a47b8b22703991862bf92069320545234c5fb03e9d6657c2b11429;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hee6efd78aa893c7638c71599a99877bdfd8971cac0d5e58b2ad85aaf86782715f7df2856132c01b4197fa1c030dfb79833bd4516a4def9220fc65bf8812a22de8e1a0a0bff026876558e2eacc8782ef81c3d3abcc64b18f1b1a9156b9bbfd737faf86a12ec9bc70712045b72c297346eea0029d7b1cef3083948783c76187587;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f506b9794099c0985116aafbd648815ac7b7482b32415a94503bb4e15a4609e5bce1edfff0aaf365df14d9faa0a5c721aa4bec75ae6487a0de42f3237ddfea6714153c19eb6de23822aaf330fc06898a763a6dc8c93066452ab30643c245f987a07e242b067aa883c876963e90806e73244986a6fbd86929939724f9d66ba44;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1969bda1c8d54126eba4f41005ef72f4f5a75c5d215a629fc2ed2c40b044ffd142f7063c9a93b9ca0b113ff038f5a07ea06dc9c22c7e97aa7e3d5b59f96ad73c537af511195512fdaae2cc1bc9e7e3e497c6b4f05688814bb2928fe93f1114a393a680da19fc76910422b2ffd4978cae0c70040d03cd30eeaf749a2c79fe82b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h988cb05f1bbe7c31facdf790e39cc4f77d75d13d94262c1772f8e407f06823d59d993f93fb7fbc76bf7fe12f2d447f16ee2d36e2fb2b339be8ef8d9d5c672f701037299dd947911785daf4ac9e573c0b2e2c7603f06a10b3a134e7284fccc552d47c7268e1ba48d6bc1b409de77985040c7c33a1ea8ec82d66e1ab824bdd9996;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97a3a4ab60c9b7a6a0f2fb8a3b566c711db7d1fc4259bd7297abd87ed7eae02c8b00c7835d78f826cfd5d7be07cbe1ef0043a0630614c05cf9e83e4bf2a7cb1572d49c04310bfb500274704335675234044bf0fdbc985224a5306a51cb97cb83c8eb4582151868cf17e818ced7abb6aaf75a5dad648ac47e60acb379b885d619;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h572f22dc3b2ea3f0ddb48f9fcbade34735b9596c9c5043fe20958811195dfbb3f6f0e1d828f591901e4f0cfa1a8106a6b31aaf65559413c22cb681e2037bc18aec7b369677ad1fe30d7cf2208451b06b12aa56302475cb8a62cc03d49c5e454125fa52f2538006d9496e308068f8d8c9b8eefdc0d462186a930c776065769267;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h945ae7a96c42a5399881024268c33d5c3e0d4b5f45eb2ffcbb697ef5a76c93a8bad1c340c03132dfe487e808b77ad0a4dc927e8f9ecbf1ef321e415ea00117eb9dfc7f5a996e8f2b4d1d4ea7a63013f293caa0ada7c1349334fe3b9754507461b45e26d2f39e855bdb36dfa887fb67b23e705e800907c626ebd48bb204e1bd9e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a5a45f5c94b525ed20c3ff7b3cf473ef6fad82c2f7b28a2d60146b8ba72f9dabc2193e10a87294fe84ab84b24719697294d2a1b0f4d44c2c0b0443931e72dcb5fcc21b42220e7372862b4e89b685dc0b928dfbf81664421d9d6706e528f3eb34b836fa5e8dc14f07a7039c8fde39f428a96b76d3b4af5939718caabe6ebd9ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0a58ce4b84142d106bd84724cb4bafac36decc18a69875debb1b9d268a326dabad641825251ed8223757852f1b85ca9a99e40924dfa16873c377e8937837e0db2040d8e0afc5c5b7eb8580faf0dfabc7c1be266a74ec1bfc00d8b4728a9ef71e05789548672fd9aebdfa03d1f32115f0a022f4025bf4efb8e0a588781e3ab57;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3af6fa697074e2b31b5baf99a2bfdd71af90986eb2fac65feb85726fa60a977b7a0fabeeb3a36ea7f1668da467f03e0415e772b7f76a805f76ab9bf0fd52d9bb7747686b85951363bb8694d03954bc29a636bdf715749788b6ebcad835ae4af5301c4872df355b902892817ebf1c11af27cecd49403a94da5026182b2268c9e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc319ed12a83d3d4a600678ba7504aad1ffa1cdf5126425d9f55deb07a723a7b08bbc080004cab3b77b3327e31dae490573e3af51e59b9a14c3357679b7d6b8ec54b7dd2f0613014b2fb363186c831e6a1a8883ae2ad63714bd7fa89116bef99c486b31c812850dcd10f2fad709ac919437bc5775d67d798fdc2aad8b0c57e874;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hadf9b4df20e954304a0bf0698c24a233ca27299e0e3c01e30aec0ea5fcc7cfb22008535942ecbfc42b9c5b06cccbe67a06bde14dd9be948fd70d515b9844095a2e34d2d86d42f2ac1b21b8bd18c3b433166abe377dfeab480011833107ca5638b5d02fa98100ff83b4cd6d354b765fa0b5101d6912b6af50d4ad7fef56cb91a5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20fa3fd69cefab95f02b15cfb099ec8f6b4148c1acc6d52b4a6fbb60cb038a8479fddf2699bc6e7353f4c176bc6724a6277bb33c62128302b8b015c05c5d8ce09a0ddcfc51f9ec59b8f3bb8e88edd236271d30cc333c2fe652544a84a8137591f36f83596f73e3bfad13b5c0c3e13f3e3b4d2f1cb3c62491a9503fadbf58c2d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h51af3218822e6a9b7588f1cc9119570e77755e883a704ae332ed01d0a9b6c31a1bbff0cb19cd775043f93894fb9b2ad8e0b0fb91538e741dc68c9ff1d1c498d33cb9ae162597f68fa237778c33df16f41102cb61812cb47f3306798cfc3b20758696ca48f03291b35f0c99a0c216e82879aa061a5dde976007353fab0ece1833;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h81abc6ed43f7d16446bbd9ff2c94298aa992e3fbaed97f536d98a0951d4b29297aaffa8cdd77a177eb8646e3e8989482497c0d7785449273103a5bded920e8e35cb9093849b5426508abd4e19d7a79285c913cb90a97bc336208b89a0c808c252856ef7c4961b87b2ea8966d8da3c2fbf0ab608cc6ee2f6d78a1786a840353d9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1837be7a9dd52814bffa348c106f114bcdd83b82589a94e09b120c69cfe00a258ab012368f9a5268987e6e268c1d483443d37f379dd2005311c1b62bf96396e3a26a1469093afd8255b0fffdde84d14f7a7fc969598c55d3fe7ca4aa6f94e03f1af19a24353bb989121002e1e4a41a694c02bf4099c3966f0a33c204306196c8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h96fa0cf7e0c0068b0139c4b6168de4f72507d35075b284f3482c7b5c8bc3530ab1b46988a26e32d5b69097287a78aefb0f73a7830aae420c517828015bd6884e112862ff8eb37ad158dfb898534e5a1293e53876bf4da0451b8fe97a6aa9ba89040be98f602543911df7c6c7024f642e8bc21d8f699f36507b1ea352855fd2a8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b4e7e6db8921eb44f992825c21108e388ad7f2d40813d245a39956937af30472ba22c35ba55f3eb9676b8e52b3acba22a621d3d254071e71446979b42693e54f84a89bd49610e5bf08ce58cd0c5d00f897ccbc56406defe950ea7c17864dce9846af7b568dce9a2e55d463ae07be1223b8b139d783be7947c1351a876d98b23;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf0b3e97c62f0b0b0c9608e2263a020271dfb83c53853abe881643587b45893fb0cc792f64d744bde2f9c04960e91e272f32ee95af7db68bea60679e0be199c31c8191f03124ab7f4446754064cb49c9860eaa58664f092f0b07ebf1d4355603e98bd0f97f9c70a6592164c8676d42e194d4013ac23f9b932eae162bdf9ce69e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb3e080308c8beaddeeed055fcb104ae9c5f814df8eed4402f9e861850616f7488b5201c6f7333f43392d39a77ee4933bb59c4652d928196b1ed21778123d8b88a193ca3f36823577db1f659c235036c993759ec56877892e17cfb8a8080e1c43ebb162889c8bf48218baffdd572fc9eaabc5677809abc7caec028e6b52defaad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h96ccad572a5ed4e0185101b9aeab8e8a20173c8bf2ce3915265d5d082391e946823eb9d3e6d2e50723e131225875099887aba2d81ce759c3d7ec8ccc25d91aa68e2f8e0dce197fca177a69c2e28668e7ffcde5cc3c3257b6e7fc555a86953596429171a0efaabf12b0f4e6db0f43ae1e2100499fa7f71fbeada2a8ad7d9861b3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb04aba38e5914c2cad85364ed29a84710e95433989c531b42b4ed15840f965f1bd785baecd8efd8113b97a7ddf33b8a129a4e5c36fafda0cd3d6f786f48f37c190783f19e02a3370734c487be179dd3cd1f3b12f8326d630aa0f9c7371dbe9b2fc052b0fc3f6c09a9adb877560a4547ea99b26a37c5edfc4b62f84d1b8af166c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e702bf1d86eecd50941730e36613959db26b54543d8c8ea810cedebb97652781ec872614137d2acec215ab66a7fc36454c55182a78c1f1a5f7b3701e78b00f8b9994aa2829dc1f4d67a03cccadf09f090b8f52bc9875d2274c08391631aea6cba72e935b227a15d8d2c758b0f7ddc33c00257e8ca8000535c45caf0d7893e70;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc15687792fbd959a6f03fd3b21961fa22eb8d48028b494386f44c9a7a0671c634961a7150f9636d78e08a3ea6c830b4405e87eca96c307f86c88f6eada78981f16eb0fa72698cd288d73f2d3458e8d8197778b98b1d0ecc07e2b245f465c0c686cc2e63c870491e5cfa4c8f8c669a80faf383c067d99069b82fd2b1856d0423f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb639226428be5c995399c710233ebc3bbf92ec9351bbacca85ffa29f7cb228477e35a9d06c12f87bc24aabcd3b5d8b088925aacf4dc3288ada1a963fb457816a6e76a50379ffba8e225bacd4a73af4686ae92b34f4bd2ea5a14f6b1916e9f7f32a5c03dff7c5846b746ae38d9c4161ad20f5c9311d6777a8d47390ee20e8bcf5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa8edcfc6ef5b3bbd165cefee5dc3e6eebe46424337022533fce217a4ff5ce98cf91648293a5e30a1fb7e179dd4a420c48a695e822991a165d9ffa6c52774af98188484ff239d2c182c4968efbacac69cce1cb60f59c5b4135e3f4ea397d4d90ef9be5338c340b54a555295b31d10da3a43d1759cc6e7099ead01385517a7bed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd893f1017642dbd78af57cac6b525325e0943d9051500112515a6f9b047262c385fb9d469de5ab19f3d782db9e0648930b75ef7c68f3c6523b9409cab823fd18120450e5cf00bada8ff4a1f55b6e3cabed43795c87c6d1a5a763998faea2d8de48b72e11420ed3fbb641b9d3af369805e91fc056c5f85ec77d7a5359e339d804;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15dd7098186dc261e3f6f55eba472b71122d597dec34ba989f94050b5af777450118742979141f16c5f9e5b48c2b9f6afd7464c0f1efc0dafc1a7a571acbe7a2fa509506a94b8efd0d1fe8ac00cd79fdacac292dda778191ac42dcc920eee8c76d851bbbce445e971325e3f187861162fe494115dddaee028af0e4b7864cc541;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb4019422e676899bd24bebcdc5f8578ec8a8d5c61564a41257eb719c111fb0216d44e7db56b017fc712e7d337e2debdfa308fd34e318e5e344cc78e465652be0c57b52aa30cd02793de9308b3ccc51a7d13260687d862bf5d0093bf7151ca9c6e35478294289764789523e090f54a27b4466dc5d65fe2f58aa0c90e137098b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd3cb1a256c46b20d61d371dec8a9928f1c700a501d68d6255c16e068ceacbab680491ab76c930bed90994e3463496ec1a683b490ab162d85d21e261908f56bad0e612788c3e3bcf8868dbcd8595cf78ff6ee8e266eb9fab6bd434da0a6339335e8727ac73752121f21398c54b57402fcc93f503c94884543af9c1d35d3146d62;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc69989a3843c5fba9691ae5a31df07618083173ce684ace98a1ac9689774acf278048645c99fc48778a414dd3de88fc195709db1fb1029dcaaad2111de77a9c869d8f34f78dbfd7b7030dd7b449a5e04ec2daa11cfa108b905dbd1f8b512e2d170a0c5d7fcb6fd9f5881aa9323e43303a2b1af2aa4667333e7bad6d790ebbaeb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3afba4283781cd543fd0081e6aea79a0fdb05122d982c02e28f572aece7711ac2b013b6fb83ceba85ff621f025d79ff42b96ecf18f472d26277797b56a7a4637b322c1abe10e1c3a626395a846e202c76a5833748b151985d54592a968127d010654fb20cf72ab83fbbfd277b321ac5278e60dcc687e5e4a89f18768d9cb9664;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h38896c1bc416927003be779b6971a5a1a8014d32c122cb3bb635e36d4c033fc224aadc559455d86e036324cbcc549d61fcef6085d7c6113c0668070b6fd31c64e0884c6a4b33d96877576049388b5b5f60a48d9dbba95642399ba02f2f48512659263854eb35b2514e867ab0f341988c01fb400f561188df38d79c46765c789;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe13f9a78c2c5d6e6e79c68a5899e66b227dbcab057eb7dc09cd67155aadc30804478d41b08568b2f133950eb45fa4eac9458baa97e1b2ec79dbcb62440d7820e7e39b0731d6e1b66561458067f6ece494908e4d0c733d1f4cc1d210e5d56c141b5dd7b9e44740cb44a0d8d76909e9e4a8f059509524b74b00e1693398e74841;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6bf9a270fffbb9f5d2cbe2c7e85cd9eb9fcb8d02ef31fc47458cb9cb75ae09c0f97d783f06ee7845a46cabedf4ae24240040845c7a14702871f6ba9e7c52c6780d10131adcc380bc2402f62f0be29fe5d3788427d8b07d07f65271cd07a728c85ac30e9618827f14738fcc4f0e5450502ae99ed0fac35e2f5cce42533f8e0279;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd453639325fe721ab22bbdb3f93cd00101299caa38a1827bd5d665ef04fe78167543f3e836bc493f3585b5718a81096fe1e62af84786c9fc7f0fca55bdfc7c80fbd295824b4a7dc76a4360dc8eb747b963631b4cb2cea8fbefe05192d7df19024d34aad164f52d0a04bcdf991983f0ba71987541812a5dd0966e473bf3a776fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5c815c53cb323dddc806c8a63d960c8b6dc38a74053e23064833c42e92146fe5060fc79cc0d595ee11c2bc7c5c978daffc5d0074e5d35965a86189413ec877a0f4225d7db1e1f58d8feb7054a2ac3004759e46999d3d1cc555c3aefb5dbcc96efa5fd6a3dc2bdbc58f0993f7dc2205cc919d139251d867609908fa6b8e4821f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha6e8609db5558e726a89ca270fbaac5fd297c5fea5d9689f03f24c0681c3f5f42ef05e585b0d7f91adfbfa05a40703563009957232da16a9d3f96376bd7905d4f2aee5885621c5dae548e5bf85d4d383850fd69ddfa4a2e4b4087fb4668ad0e55da2dfc80ad337fa06010e5228cab9f450c14488ae3321977b1a2159e21e83b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h49e6fbe70308bb4390ac5fff2bba821980b5046c73e3a5774c48f7af6a0a090b3773b7f89265216a61739482763d431fab3dafd5a7216cb11ddf10095b8c797048f4b98c3c43ba1cd5119099404add29263fcd3fe37bcd3bedd49b86eb4a8b959b8fee17684cb6314c27954d5cf24e193635794070584c8cb0b6a1b0b5786a57;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2647b71a4980dc67ae86c16e970d3bb0cdc841a8b08765e3b07869b7ab32594a4e78233945224d6809061d2c77202cb6b6b6c14c64b2661c8349f0e59b7ac6ff6f3a70561c4333228c58025f6c9d5b35c26641ddd02ae747d7e493bddb53a222c437cfe03fd76d54b05b4a4faa910a67aed1c5c0ee5e3a010cf5a2cdf41a8375;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd073587f5509368e77c5f1742b658e7b67c8133b4066171c1ba973519542a79e53add280c54cc6fd83a7f835b0f69c77fd3a01916544d22c5aa0dfcd7ee9456b70489b6a2830da1da298a53288a2c06823abcaedf8ed197ac53cc80901b8c9ca924ed1af70d6a442887ef742b32180567d84b846f6b3f8636d5e2bc861e13fd5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b32a24c6cb3d010bbf790fdaa1ea5df1ea1e88f75699ab48b1ee7f87364539f613fafab6a70a236c5ae3332e6af8d45222fddc222b40be4640853fb155737e096f344ea689cba5158c821b4b8924dfb6e70346001ac954b32f503266d20c50ae6dbd7007340d839c3c53df8812a3269fdf3781b83a65510f2ff2986abee2ab0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b2f8f94bfd5e64b01f3bf2dfbb9b5628f62ed44ec9ab51d2907ed747a00976adc9b172aaa5e5c54c60a6c6bf0c80e1c02293ed60172824e5c1f4b9050d946007cd11610c35121062da4f57b8d5a94e140fbf384c5ca544847f09be7527e636657ff59f81cb8ac1ac75dc9a90eb635c2d28265e770964d829e769601909159d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4eb75317d24c914a837e8f385e166b29c155b3b1a657ca810418e798a247cb8da85fe40918353ff4b1a778c356e7bc82e81d55bb40e1b0f5ba564395aa1ed18b10640d84d856ff16d05eb2443bde24cb514e5079df38916d12e7dccef40afd455c9d4f2d80cfac3882296567ebc7c28508653ddb81f1f9391e75eddbf4e113f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53e40205c8bfd11c7a8da012781c89cefc75d3367ebd433adead0b4f65dcd4068ac2a97a2d604b5e568a3ea3735313dee5e1325041e50005ee09e5340af907ce4b051935b96df1c14f2cd451ea39ab757c4bc2d8e9b41f4edc6797e2ce0f38094657a264e06b0da1cc419ec07b89530ccd63d85f08f9cb100544c3fda37bfc6a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50b9c3021b4628541e6ddb1ef0768731487a8917ecdaed229e1eb63d7533a37b59d497414fbf308af874c33d959debb92299e9167c6d68283c642a32d8dc1900b8c0b4db2ff6ee760958055578f5d808814145b9d0c7fb360cc7a8e0f4310961aca7e355c93df9eb5d521eecad4c382ed902b8b77e0ed1840002b415dec226f7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b70b5a5e196bc131eaac6298ea9bcd04844a80978a6d3676ffc0e75a9ecb90c682df77fc08939045436ee483d6ae20d39ba6ba2b1463272e24a6ba3d70f189321c35d0423fe507500cf30094f13fd209e585f3640ad967c4cc96b9123c575e2060a038ae2d8c71ecc32414ef2ca30003b93842c0e1ada4bb75dcca8e1786f67;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2cf829b44d82f1e69db7e0522f0463ad8d874b557e41598ca6be50329c35575f73b1a339b4976d343fcc95398e70c215a76689be1432a8c36cc433600d63c7240b83eb33484f59817ffaec06b884e09bdba122da5dae64ae3eb49fa9f407e9ba0369d585c522dabe19d71927d9430ac7a037f5944d863bb983f8710c6d434ecf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc2e2f54f31eaefa10714d2fd11124ff3dc117832fa9da8712f303e4bf6b24851af4ae9ff7999e58fb99e7069c7530421f685ef676cf00d394765788485414f65e92c9e0a0d4889e764b8f7c1728d5318f37da2659c923e0621e7784ced52b99adb94082ae3b309646839604d7c973e2b41fc94534502c48a612ce29ad9f00d62;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22637beb27f44a6fb608ea4ee46151b2ff7f383624bc46e087ae183515e4a251685a873985e1607f80c23e3466e1a829851187f30435e7e9708f7288f2b182a478f76ee87922dd43793e32eb85d47e734eadb09ae6b5147f3a612563a4aec62d561b3932ab9dfd0aeb8152f90d8073792bda4f6b833b3d093cc3aaca4ec6513;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he36dd4e8294ccf5e2dac4c11b5c072a9c446bf4926453dbe30b8c2f3e189b22e84564e6c12f0b39d1bcbaefcd20c568437493106e616f77dcf248dd45fd4d932e5dd587b1c89c58cc5679d71998d6c51caec98244a46e2c803a040e2acaa8188ab5b61b859cdc7fabcbfb514595e465242cac4f3755d05fa8c61fc262dcddfcc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94b0a69259bc2b9c71e3f7f5332caa5752c83ea91361788d6c00eb0bb51a209f7e7f1212228f40b7fc859fb935bdafe9a7670f14254e2b10fe02c332765d25fb94bb6b07b87f2cbe2cadeb77b728de18bdaad44791470beed713115b04bfa6e5ea65b986f358a2412821fd37e57f9383bbcb4357411381ee67319556770d0710;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7dbd18fc48f6ece32a22f8ddc1ebae5a909a9b26904ff752c24aacadb69815fe9f31ab67bcae1f8d43c33630d6e7c85976b5ee1789d09573b011bb2b56e51c64b818ed2629676d141cbc1d58617c403cf4ea72461957ed5c0bf32b4304343a204fb259b50cf0315d057d9a3e74b14ff39fbc81d2b5d4870da7ea5994d79b4a7c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h526aef8376afd3a55b7fc65db719c673f4fe715368019b1c8788da4733162cd54eb05652c73238814829d9d751bf6f64338222fe590bcc06ad92baacad9c17380abbe9d1617d21b4968f4f9fe2e9f24e64378d2858b2b551723eaeb3620b3cecadeb01d75330d92b106c3ef5e9055fd9ac28ea8f7af8bf106a89f45229681a27;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a9d7cbdfb9dfa56d1fda6359a5570cf9441945a0c77384a4621b208716009dab45368db9f83cf1eff550bdb9556957b60b5145bb77c4f1960592b80fedd4c1b8b343e522bbca3f43464397c608b05f5aca01c61861ee798e17302ee6cf8d373633fe904707836a18ae18f2f50626c7999f11bd93e6a2740485d7a84a0ad5ede;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b18043aed08622d729659990c1bf4d2b490255ec9444e7b260fa75231bf544d90701feef6a441cb93c3428dbaaf9782d0949bb3d6e80141fe75dcee269edc5bd73816f788828acdfce3c4cb69d40edfa54e96cb95a74e4da3f4ec011adae7a29486701b6dd7ffd91db32751ca021614da6016918a95fb8aeb32a055ba2bf93c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h79f9c30301ea6355730cb9b57f9a05836256e8a7c62acad1d1b7549409fe33997dec001c9a6e6fe4acd410af710f88c33c6fb6179d8400c435b0ba87c97a48823414ff26ca596a092f7aad24ebf4a6c2693eb0aa91cdac042a9654d9d2c990d1992353148f6f4fa758204fad47748a5df47bfde5aaf66694e5f5122cd5f21a1b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hed7b71ae16175a8bbaed0d6315b12c7b237da876cc34db766b23170ae74d09c99a4a52d1edd22d0f90b86414cddbbd59e8fd9730feea56c35353e93cb44effad4f61d729b652c5cbe5547fe1ba3e76e854c643ac2f04d3f5d63a9c1e91989d4891b16dd8b81a4c1efa5f6cae158ed9671adcc805a6a64f11de5c6db3c126ab19;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfd79bbc135b1f3a775e8b35ce6f5a3481af509f86bd9996aac3e3998a8ba39e6cbd72d7e72219c92f4b0956c9f0f77478bbd11785d335c24b791eeba2b54ac7fbc74ace44fed78c894e5af1191c30967fff9f699866575af68357f007f817e250f9db406d6ababf5e6d72be4da4c04e5cfd3e487af08439134100aeab15e13c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d2e4dc9a6967b34f9d7760733d81e25a6a03c175e48d56cbf060796863d933a0b7846adfa422370f89a26eb1582bb93138e1e74ea18474787cc6919191c7c72e8618952f34fa6a949c7fbd30b8105b66d32a3a890b80ab4e95fe356eb24463698144d6bda3d8568e4142e5db3feac693eb3ff3bb8460d86888ea7f561ff82d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h340af7283ed2b9334059fd82cd2c7e1cbac4fbb913bb8d4a45f71340de138352004d50e6df420ab0c51673021519237dc947d5f7b2bf0d1079695ca43d680bf142586e5c5813113c5a0aa1a8cef2a5e06ced002b576c6391ef67c859f41c3d61f6394d1e03946ed43fd0fa9067519ce17e58e8b19851bb947a00795e62161124;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5fc03b15776ab46c1ea81f51382758298e5c35f9a810f00ce852504e9dc24ce585db279a11ae2a577849877a4786a271feb7bcd376e7b97f2138a754023ba21ee1eeb0d2f603bba40f3d71624975b637e611c93913d7520c3f8be59d6ca0f58a4c8a8c6897ba0d8b45c83399926f9b79079ca6c734e056eacec19784925e891b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15ab4cd86bd0777dd1efd6b7ff1aabfec9b6e1a20d8b30cdc3df12d142dc80179ef3a94e6cabcd639f37d31f6592d15fc6647cd8f1b85ab36291e5604b9acfa58fac71f786a197cc6d3cf6b89870eca2f41f43b527e40f29094ea0b3242642e6d3b21f8b3a53b11549b97ff449e2941b59e1c0e3a567839e830c759406959497;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha0b639dc2cc7e6273f1420746bcf5a8a2872457e605068d00edf2e0218d87249e9d717494f919db6c9a2addb695b6c3faab88a4a6d8e600fa9d58599840baade8e5e78f7ccf6a38c10f77717199e6bbe1fe5d581e475893ff925a19ff0566918ca187000b3ea7bb36f8927857b25bf1fea6dd24a7e924a456f490c389bc2734e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b262807eb077c388921c324c9be6afc6686d17db6f82f5300ada615a98315dbf6af7e9d9dcfceae0ae9b916950a8cbda29bc0256a3886855d3199def54a8453bb5ab0ea4ad4b96d9c23daf2eda22482f14b4b2bc3c637fd941a887c35cfa8e1184831254b8647c16d25d6473cab120fe6aa5995587314b07516a22992332f4d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haeabc851adbf8ac687b66f929af5dd435e5ac265514d2a951ec2abcd073bf4e981f1d2969a30a2a77fa5f83f017eec2f9947e73b2ae150c7e28080cd7896883f1732d1ddf390b9c391f7d9be6e1e3c21bf312831d10bee3f8d5eb4d44e3a6fc4c267d4f2b293a0420fef7e0be6b8a1200bcd39f6695978b8d42a54f75bd09c31;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6abf76191d03dbd2126364585ff2aebf9a11a83f60f3ea13eac4415ec84d613b12ce1db5a804804e489a86966509548779be8b41979a17353a66592b40f48bbfede5362ccf296f54e17fb2850bcf0e1ee398436a76936926ab3df7c35c131c0260fd1c333c724941e05843e9cf2f0cf2aeed11b0683384fd8ba22fcbbec7157d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hce3c24d2c564ccdaf5d58742d203cacb5dbaca1afefce167036be7aaa1cb05d89b9656b1b775d897dc97fb4b4ed773c2997581578093db90ff3ec59bb84e853f032967e8a62f7b8cba1b6cc7959285577deccc64df2a634e3eb011d1cd7253b656d8f1d553065d540c97c8ed8092fe9e9046fa81cbb68fde5a5bdb4f5f14b596;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3cd80c54580eedf5d57f7a1e9356a36df186e4f52db7d25402e9378206b7fb35903d4693358218dcbac5db7779dcb804a5fd9c178f8047d69641f74313d17f2265e17e51aa3a2d84e9f9d10d3c89135660f0e00f35a8b16ac1bd00ea80cfe44776cc139e6f64c10ae99deee8beaab2cc23984e9083d3f3e66152704dcaab9629;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd9bfb875a0a369a29ca3d3fe60d89cd226f2873d280a41693ec70124c1c6eddba794ab085811001f68400490d0aa969e45790b1ea77ec407789ec9e8d72060fd504b08f3f9c68bd9953b80316f374cac7172bb326802d5c20cd3b858b4b189ac71c4a83e6acc46bb118298aafc4f64d5d711a8f8aebff533d10808e58cef05a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h791bd6ff58238d76e491fe04ac587b6930340399c8d2da0579a0dc93bdd3ae1b310d58291da6bb4504bc3fba4cfc44b7397b2b4084af976e6aa813f44de399c8faeb6d7cdfe163dabd88bb9711443ac716be18b23f61dc9443ad47a6d6cbf12cfeb3fcd205873775d750bb9d17e90587bdd88b4732cb9daa4c5b70c840ac9515;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he56226ebccafdc2a0df2fc254b1908a56bcdebcecbaaa9afa42139e4a380032451ace23305b49b655f30b73a14415c9a07f83c11204448b7fa40482f71cfac08e3fc259e4075629f86352dcf6364f5169f933b0084bfa8188ca713fe67bf184b57315a0beff393537bd28ff851c38998f2a15b73d73943c72118c8de6044516d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he691957817468bd070841c2ddd8c2a6002b8a310b73159f036c30472cd87e7b2344b2a4b95f15197708f874587f4e1c7f7b13f03efa968e63f183faa4693dd437e97309e6832a3253198424a3692a9aeea308709e7bff1796b14e2a3fcc2a8232480389ba4d96bda898e8b263780d027796b597672a0dd23e8d318407d3f2df3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c005897dc42c9c1e4809b1ea3732ec42a0baf64216a8c26861ffbd086341b946a84b725464b8b936da44ec8a4feb1b799ff55650e65004bc0e64fc58d128968aede8c5c91bca48c3aa283941a49c6902c2a6330e25c005d0d317699948461a0c8025b4754315463e9b9576ad0988257f00ff8dce4f1f4c4a2b5d7513f61ac0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a1e709c6d058c5ee2c54d05f016c5350e9548ae343b510494c954ba34728b03142e8b0729ab984d8de1e80eeaa11693d8c81bf49385b809b2b05a0a6764c327f82abfde9b87d7b8372600c94b5d1242ce495b435b15f51698090e1cf48a6708a4ca15a3517298b38862a8a4bd1565278ac3b8fd1b8ef5a8cb4d042ce593d4ae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h969667713ed6241e41428b4e7200d783bbefacb1470ec0c425cac90d5338d3ce741ad0c021e49d657406fc1feb86f4926490d883bbc453cc743dac452e7166630a6dc54925c50e7aee3720ce32274c242be14c2e538ceabfe2dbf283cb7bd98d6eac679bf36760100b9a3ceb3e7e7ef4838028be86f9973e08673f9588dddcd3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8867176c85505075dc682b145b68e59cdc7463046f8087369f5b7af713b9f7791f41347a5dedbad8b4ffa3f57770a9afd43e73c4714ceba530457e26df5b7485705982dfe4ab1221e031cda674943ea54edd9bd83d332fe8d94fb84977b97730a059fc075b2d26cbf22fc464b14b07b824e6a5ea024b6b78af8f0b517ff862b8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b472c7fa8280ba435b16a7e6ee10057ace6228bfa8d6447267232145eef0800fcbe1bd4a09c24e12875b6fe2638bcfb427c19008480cec0ad5f9b238a84b97ca69daac781c916bf33c1c3a7d49bc5a28b6700f99f2b8c7656ec74801e94020ee92bfb26d26b7ad469dfe0dc5059ce908d7001aa50335ac6c341b8d348d6e4bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94a3e43a1ef683eeb7f270964f4851013f7090be368bf48647d19fb74cabe263e1718cd67b8e767328788b8cb0ca5b4ebb04391a811de900b894d46e6d6ff038e7a9d1cc49c75be552d11812a066eeb3389fe2fa68e069f9c05c0c6009e0114e1b25fc8c01138c40cae96b2828157b07d46045c3a0ff3647fac8c45d2700597b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1d7bc99e08dffabe374021b50512337f4d8ac6deb1e58567fccf6f154ff525286760b420eed4e99a8d57282cb6fa80bdcc70903aaaf6c7f6c6c6d0390c0fa2c396854e2bbc432322e50ff28602e0c6d0c5e64bbca3ce8420ca347ba473ffb5fa56d2712a8ab61f754d4e093341d342abcfc6459164d1211827ab16b2fb9a3759;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb03da3b5621cfd6fdf16c34f6cf8e0a1d9a72a65a5d14c593d1c79af2c0f31e289fbde13ae0207c4760aa7ded2d18d4e71b3411885a2b972fa87d69ff907f7e7321122d4a275f40c3ebcd826ab3e0ff598155ee2cb397ee88ff0f9f463af0b19190ecbde05d9dbe564546354269eee5d09536fae08713cfc6f054581eb31c7b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b25b520f0ecaf831fe43a00e480f6ed7941855522b53c3d52d2fb6a8006d1899c5970189b9fb10d77b023f44af4dc4e248c8e753dcc53f0fd5bed8a7357513646be2beb2f21b4b8077698f082269f77742830a6da2d3907965eac6876b25618a471e06b99540a7b299faef53cd100bceb8737198f46d19eb3d05ae91ac12dd2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9ce7a8143fd909a2e0e9fac5033a410e106a33b0dd9a59ad7192ebc43f9f11b52db12736eb6bbc13cc5b447e1464dc46545a425ff38377a92f2e1aa4e58540a3e3665043c3f6c3b1957fc76297678557e63520fa9b91aa860ead3c107ad3bddd15a217fb833c070152ecc4266d30ab915fc6516b59890f59003024aabd9394;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h808b2547e57eb5a66ceac93c967e90285982882d9068ccccd55b0657e615a7efcab1a5d7de1dc3750093f6c17687a3b54c4e1d621e36cff929c48a13c06e6c3037c49c32a6eb877bc00f535c53ee282b4fcce91669e5c01998fb44580555c2d53323c85cd2a3f65dee5b9940930a6ccdfb4599f17e2e2da9043b4784f445da13;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3ed1a879ed720fb35967b2c3ac3e385531ed9e17478d839dae53dab0db727aac26e26c6ed3e1ccd76f3c33142646192df07fc8157930214369a490e78da9c9ced61ae79feb843522cf9d42ed56355b5be8d5398cac65903af2b4c0c2b1a212d1dfd39f183dcd2f962c1a1c0a494aec6f7ca0e8ccc7d213246d96c7c6a7f8a8f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7af16ed66ea8abb5e74a0c5a30cf2d598b5dddd5f857991568a70cb1bd21c198f81892f40485cc839a3547fe0df3cbad820e2fa0da58650afc43d89c071ac042f3d4c5084b2370378289e3693687246e5dfcb974c03b8f98b01bec6dfc831043e5f4b98c744d1736fcd2f74d467236e380d6af6f59f14b2cff636e5fdc2a66c2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a703100164cf70caa286c038dac874d7325fe56cbdeeede1695d82425244194f3b4acec3eff9c82c3e31060c19c12062c616d361ca16dcbeba1eea11b43de3d2ca136fc53dddaf8beab3b13830fa981c7ea7f1d7e64441da7c00db3aa03b2d9cb46e08a935a92ade1b299877ee65cd6e12b3296363d577aaa08b8aad1c24443;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h855cfb09f0470a52f53200aec4d068c953e73f0dbb6b0398f4ff6185f09ec84a64f3497c4fbbb1d1fd9172b56421ec77f30f84b1e5cc9268c24979bc0a5e2e5c95548bf5d8ef23287b1804dc5fcc5db2a810c2dd2daab552ec6727ca374625ba43491a0d9802dcca54623eef06313705431b2396a811294c2cf1e38e65193499;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4da03ba43d07f700567de6527f0ef9b70c44c76921cf2c0bcabd2d17edccf782d99223b31481a05ca6a224382c9a0ff5de2793199ce652af6e134c63301bf84185cdbf29b496c18e9b2490ce3fde6513f4e2a797e86e3fa7d3e8351a2a4b34e640129443830d503db7111b71c2aa44ea0dc505a099325221469d5f878fb6fd52;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb04de653e87ce089c97598f5473aadb9c130a08db9d50357f5f4f47845878d4866eaa16ab63f2a7034ac06975b1e0e638f75a1e396e264ee80d69dcaf03d6b5a51b054b16409ee25b182d4ff450b44fc883049b956f931b9c1e50f44785cc948f504035c34342c53260240c75cbfaf46d8c112ac82e07f4a2b0d730171fa8525;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd10069b9b7e524acfc74a08d94f6f23c42c2cedff8c39c432565ab7604534ecaf349ef5b87faa080d13e0620cebe2a42311266d8ced261eb02129167b419072cfcc699d8949d4d0636ee770cff37a410a6bb40a8f9153a7eb5b9f50d6d8953fb70af5cacc062e5b03e03569fa8656361b0d4d01c249dc52b5e553b77cec523ce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdbfe04297c15e3ecc4ae1b7da566fb701321cf35f6ab46ea6e28ac730de5f3de61592926ac355fd33a4bb18b8890c2f3b2342f7d0b5b1abc978befd0f7baa516de5dd08aacbdc6cd32d25047735e7363d0e4af2c7f7f2aeecfee50bfaa33967a8f211ac7618972b83c0db33136799104a8dafa7e80881dabf78a6961303ba9ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf0774d45fb9db522ec3413dc2ce25d6e780426dfc2ee36103b03601c811b26171defdcd48befddfcf1095f6ba20aee30c1916def994695ceed23b4758e6b32e105c9b0e63e4f1627dcf4648c7fb1aafb3d99d6fc66b642aaff87e2d5d6bc2bd2a962a02c8940c1458efc1af02ec8cc54cecf9cec77fdeef9447cf268aa411e2a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50806e3cf69f88e4edfa75ad31e389076a32c87a2dce9d13aaeaf051bacb628e772b11ef90b9fc97435b26a5c3f2f3fe42315f2d8f1f06782b568aa56c12a1f4970798b75ebd36a96a8ada9c8a81dae5aafd25ae04a946ba4dfdf51159cc5d7f2001408a3c0c12559631fa56f1f23a0ecc3fa325b4d62c30d5f35d285a165caa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he927c91198b059eb55409ffca0492d5ce121a97f2141d5a87fa16b6d8963d0bc62db722de7881f932ec803be92b53b275d4891ec45cfb0845d46f2eb946c65fa22dbea61f9005da7e4a45bcb0d883de29738c7c3df7ac38700c05327c29c19668e30dae4b5eb856d0e062b96a3a467ca4c164696873cad5fe444f0eeb5bd8e37;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2e21b3ef4bdb26c6cde5fa3176a801404abdf3c02042208df8d8477b42010ff3515f079e1ad02f501177fe267f2664e9469653e89679b50d76e1d8af3c64023e2188b072a906675b8f844e0d648d858e39f70a28b9a7bb8f023707980cd2b3d563084244e9b9ba8240ec47032c14eda3a1ef4226afa0c5cab96a3dd2acd9702;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c1554aa8737fcfbb06a5ddcf15bfb3b92b9ecc26453bbb485ad945b81f732ec4e81845d70bbe81b45d3209306a14f24b9fde3b1d9e1750b71cdb62d3da4246108c507c7c1e1f682a15a219847858d18c4bee4f80c78fa2ad115f650352f61856490935207736461974821384a4be137978c6b172711dcfb13d853d246ed6f6f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba3473b911e5c01649c9a74c3c4a5289111188cde781d119c37e444c717fff3e1f109e789353d5a5e2509b4ae4f5e474f7af34e2630ab9243040836198d8a26f3902d962a6a02d2aa1e3ee02ebccb0247654f705296c89b2e7b7a7d52b2f90fa835d42deb5be0735df48b9e9b245379cbc719e3d39250141ea34c86631571af4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h890045210d6a3ce90e531aa0727813a8dc24f2e8de8c862aaf34d1bd3395d16081b5bf9a0fb72e4a8897b3f5501d0d3b7fa3c50248aa8a1c57f133facad3572cd20bf96d588772df78db5dd41b17c18d27b9f45695ae6b8cd1bc3158eab36b37df84c061b60edc7c6b6200b3f5fe78629e77113d34f59072da3c865409f58f4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24d4f5aea4cc32bd5cdca4163c54dda5eb837bf08ff6c6dd598b357bd52c655be586f3c34b7bc42a24007b1499b97198fcea2006fe8d24b58a1b7d5e13fcedf0873a070cf54f8fe6ce012eaeb99d2e46698e7e1cc916091835d58ebefaa5491d603b15e80023c915bc9a4119a4b199c80bf8c6819b2c7886ddc8a35e86ff7d75;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52d2096a6c7d20e53cc2d45fa58231a0ecc945ab8707f4292d7f2ec942cf2773fbeed8fb4713fd0b1c33ec6d592a466028cdb74663d6598ab3ab617e5b0f17b33e1ca0c4aa50b1c6e30d2bfe0a1c3f475dbd12ef46dcda35daa60cbdef36f21a3e2ebac620887354db083d0f5035095f167aafb14b3ce12e16e2cbd69387cb18;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he88ea46c90061ce73e9e19a56f05715296829cf8c646c2119584c570f70f6e97db5ce142b8edd9d49da5c9494cf4c15afdb1a3d3dfa6b656778e023a1766ca4d13c6107bcf431f629a0419a24fd731b1b283fc51f987f98ec73b95068c27784885664fdf4d9f11539b66c20b73d4215a865e7820f8c44201334c6f0079d7af1e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1fbfe88dfe98c6f7df7ddebb54f3c7a56d69fede77b7ece68cd7b353f85a1b250dc5f9db662938185c4067f73f48bdbd8c2f92c78361340fc63e54577f139f0daef9bcd76a85d94318ab7710b10e4f0fe74fd94b1019092654be3883bb4bf575c35528f788c5c46972540a8fc300ba5a8b21bd02ea2e9c6bdd44ca4100b58540;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haeb3114f13b135b5e352067bb552a982dae472c7c609aea5fd2e7b4c1664e01bbb4b4077141f8e8f46b9fe4589d2d4ba154202434c49e9a0ebf8a5de4dc6552ed7930ae84c719971e77b9816d5acfbc7df59af65fc140c67924bda57245362fc211a26a2b9add40d13d3187c7b49e9fa4c4c4aa217e4e1d753e1cccd6c86529f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74b39086155aa0edac56d24446aa570ef8f696ee8e4b2492354a5a17f7fbb5faf3f1283d8f5af1ee99ccbf8258a3102cbb8da834f856e629565bbb3a6142483c290c7a805dc13ec278e38fbd6b99fa289989216dc1ed061f646596d366b8ed7286275008caf12b6c752171ed456bec99f4f0b3e8ccde77750c8a4de691c0ba91;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7fae3bd4e8e357df415ba5a3ec8b660b4b512c106db26792d8146aed7e7c9081f63056ff09131261d03a13222ed26d0945a5d0b0de1716ba734f6b2949c7d11b4adfd17bcaac9aa3611d3ef14f41a6d2b7a5bf1a8feff6f514d81610a657b15ab448bbef5964493638358e104dca1805859bffd355d424de7e3b35c8314faf82;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he15446acffbb83cf3c9c71ae80e0a500496a5df52969797e30729cf2742bf75b9bb68aa05431ee494080d9056212231828a0b4f162188419f0ac7da44d532315df8aea342e7485188bb348bcfe71eb67e2bc9eea54d4856f2bd8255c1950b7205d9e09d76d67b3f347459089c54da466ea92c666387c3734207114727629e5fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h56a9d7065c4620ede29dfe5ee769f73194bb91ed5b896afcbc89968ad688e4f07faef640003cc401b5b855865f966113b4defa627b9b482dee00d030aa56489e52a31fd4c38bec014f2f65bd8e6ef022546e3949f50b2f03101b3d75a5ceaf2617699b77dbec7b931f35f3ac9ae1647bd4553992821fbba6bc1c27385fc3769;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha412ca8790e6fdaee3e02f721c8d0199319fb91185bc805a97badba1052177d25891acbc710ac1faa2b9f20db7cdff1fe8fe9fd7a0d41177fa31fa181bf27c33d5bbe413dc0f1906960c13338ac4d037f85cecbd2df73ef605e9d89bd74a739022736fa8c6936a730dd295cc30280dc8ae18bcf46a64f226d5eeac721418e8e2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h178c890f83af423f351e9de7b1d7550696893bb7f773351b4c9977b5dddf5f3cde893fd1a187e230865aae776d0c27e18e2996ad8277f4f28546d89a7d7ec9be78d093085c960b3b5cf5ac70d10884a53606a6b00130324f66e43f8f9dfdf978a2b711ff4a4b2abb436456f2060196ee3d544086d3c28eb3d08049a78f322b9a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e55e43f798476820defb5186cba488f2c8a5b14fad80fbd55de32218817315a00f6c0be60b1b33a415936472e8d90a150883abb944d131e36e2ac6e58a288b4ba9fd4e2c53ce1bf67866e3be320be45ecda0851c2311a7afb9bacd40ba6a56378b7c404fe63c7d09dcc65ce1bc230c04d82b47984bb8f3da5b023a891e9d7d6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66492175c0202d79450449deb37db067cf08234df84930422ba782ee3eda890e5a6c776429b5e3308bf05ce2a543c3b106fc5ee473f07b275605846bf6ca4509cf37a6ba5f7bd7f90373ce64ebedfa5ff245c38d4e028a6dfbe44d1c34824c3dd227359d530a589b3f5f4059567ce4bce04c09e650bbd0056c053083b68b53cc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h760e530049c5996098433cf1f076ce4ad46ca0ee7a3a2265a10e231ca3d80d2d103eebf38e0669194a2aea6f6187fd2a0886a2ef617522fbdf2ad325df285f6bb0d2a6d2ab31c967a5a8f02b397672c96033ac38d7ff09af734c9ac5c51006d5ad329a5a9e282aff89279e037023bd2c52e17585eae2b018282621d64b3cb531;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e21033d14ae9b3c349341f427663a9414fd3eded24d540e8598030e092717fe4263b2fc760655c4f28285ac414b157e017c2d9f3595073104513b37c5a2ead5e355fb27ab2ff0ebe80db8cb4d45d8b2bcb3f02e01a69d0a4479f98b0514a448bf3b3ab2d590a041105de20d9ed531c21a38e0f33b930c56f4afdfcaf1aab3ce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8d4846656476a5285cb9a938e160466ae49dee4e20665857cdab6f75163935a3443ad95e328bef6f7f8a088b02a873f4e0792ee7ff444cac05e7732ac710be481441b536b1de7c1d926b43385469e16d4f65419e35c2b1ef6d83b3f6148b264aaef824b5430269b48493222a7df97e09bf08be8689d3d5f03def08bf2ef3f871;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc2291520e8a01825919ec43629208a83c5d52aae744ff6326ce7a9ebfcb678405f4e694bfc7314977a47e761d169738a12040218b086499e5c9364e86cf589123c35ce332a24f394882ad2e706f3d167cb35bcd18c4aa537afab9133311eef17babd6698829b30af3ce5d6c034989cc8a85e085b50fc71fa184e087801ef5682;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a21d138ce94f4fbe018443a70434c97e9f5d0386271c7e7a37f08e9660e3b73d12c619655c419694974334dd3b4d23b798b20aac76c96f19dd9345fd7f68d27e8cfc38523c648db57c75f590f06703c746ae46cb1c42123ec1592f15bc99fd108d0aadbbaea6e55e1e89ad8af5d9fe8fd9908c9b1083c2a21fbc1c18126958d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcfa2662ac86c6d444cb4ce77640b252b2651018262ff0698a33cffd98194b9c56862014b22ee35f09223cbd3cd5121457192751c6d2a72bba05e70b58fafd59e320d21b76e1d73de7e34eaff8562f2e92f3f5dfbff76fb118f30fafe4c74ba9d2603d99696e9cf31a81ce353948a8088775194b7ea306e12019091449c759d2f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53fe6fd2d17d2f33daa5b6ffbe183f8c743df08fdacdf98fcb563aa2a604765c19d2fd4b009cd1b5521273868f9b41d3e32946e924bb5c12b43d6d3ff306c069bbf4fd613bac6463a1cc415ab75729857106965c9ae008f86d124c6b471328b4116f24e74572024dd630fccdc10f80639c82317c8e27ba3d9e98b9cf2dfd4d61;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4710f765b76c7467e3236f605455173d74f00c886c0aac1e221b2f1301c349a9add797afc139b840deae5b2438445122363556a52e0d411a9a1baf5200a4d5735593125057b5539801d328541ea8f0b00aba81eb4bbb7e8c44a871f3576686f9d2d5aa62872ab3e5399f52425af65558780020afa1b990291528840c4226a3d6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d5f5c7bc0439d9e18323123f556384551890fcbf7d8ba950af3a72fb088e886c14a9f7c97136090caa3fafb778ad5d9d465e37e0036a03949125b45683351d17cfa1b7693101130f64c060173a79274b1e00849679f85494a364cc097260a616034bf3d0d2f3e9f49043eeef090e021cc209a82fa9668ad606f3cd9a887ab73;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf929cf2c211b1bf74289d85c533641931b9d1ca65a9bfbb02f3100c3e1d2537668c66712923ce1622793e372058b60e3e02048a1b8ee1c9e91252c90ea547f1af38b4c01f6969d2ff49e635158a83fdf1806bdb9a4cda79ff1bd2262eeac8e6f78d875a9c195607279237d0ce48101c225f21b17c62a29e3e76931019790d6a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfaabdd0bee18c65b36db28a45fb21717db0b2122ae254998bf67d0d1bafdf732c73c4b63be6de161ad468f6023d8623e4455a5eeb4ba80a9b9d662f459fc1c95c41d045c22cd35e76f975c0e2965036db08cc7a9a792cff38412703f22cbf02d36121e8293699fd605fd72f354e229308c42c2d6e7c31ecdfc70becc126fb9e7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e6b6862a43bfb39d4b58f0bc0410560d34b76370eb33d0ab117b388e0ae093caf6de405e24d9fad82c293e4b44726c7fe10df9130644543b5ccbb2b9e0f991d337ef45295533838607d2e5d2b30d85821233d9cb6c3ecab3e77df11af971a1e74de843281ab85c3d53c59225855793aa12945f1c3699c11c3a46b1c82a756c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4e61d283d2760dc4d61a30122832fd8f7465d8c68d7d61de33be605bf063009850866131072eeece155a6071d7a6d82e64ace70d3e2f40e5386de4c962e477c92e67765715966400dd72ad8fa3119bac578d4b95a004f7285ed9fffe316601cc3187a336ea0c5d700a0b0b4465164ed753d42088e1fb011af63e97dfb591645;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e79eaf78eb95ca0d11184be429a25abf9c12f19425399c8f7588df46664558966a7ccbabb459f3c823fafe830e246d128ac7a79bec0e006b557391f996c1bbfae582bc3b6ece1a6939a03d005c5e2c22d3097add80db24200695b1113e6c3ce4a302e1c1aeb6a859246e668bc67880e08660c14336acc2cf81b56660652a40e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h957c4a633124e77c377c9af2d607573b3065e55931c5c0ea610c0954243208a46c50acbc0f206c3dd3bc1a6cd2c7569cbb338ecef8ce3b301648c7750cd46dddbdd43e9be58bbc0a8567ea5e35ca8bab3603876d0cb51fd32695a148200ee4c0f0540d3107046e5955f55eaa8a0d07acec77372e168296114dc1a71d257b1144;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2ef67c21f0db76cbbdd2242f7beec29b792020da9687b69cac0b1df7855f0a8ccff8a159011df0c78fcb8e4e8c8e5b280c95f9f2aad88cb179c1ffa10ca453a9be7dccdb62f01e079e0dcf759403d2f40134b3b008e50a7223ec30444020931a7a28c0212ac7cbbab499d059d5e9b30a4ec16c25c9c1b9fcf27c8d40bd42d33;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h19fc9f2c30b5d930d6129ba5a24ceb60555d03987c046891802add6479a8031f2c9d3d4d6d4f59b69580c771ebbfeead61b45c8c68f4f11e3e8e3e0c55befc713de53e16fe2dfc01380f6a479b112cd5dac71ecfefeae0e8171312eef566167491b952a94475e68e8d988f46e09d38996a69bf43abbb3d62ca194c72284dbe20;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d8815129cf34fcc16067182024e2583ffa92916fc2c1d92a9b78a7009701c8653d417ba11b08f56c3640f103b64498cb63ae7a1e510e1f5ace70229878b039162b10a1667d9084a1f2a6655aaecaa35d03faa364f220c8336ac65dbd33b25ecec7fdbb48a7d5726c532d2bafe92eaa60a6798ade12f69bed98c4891e38abbb2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he48ddf4479baae0a81db961ef6408f2d6ddf69367b57eefdb0aa73b43e058cd8b9aebe89db68cc1c55b38b4552bc7c6f51df6d44e177329c79c0127a465ef6365a6cdb3cd17c4618cd0df691358123b7e3ce367554e459489bfc27f00b7f11bd6b322037ff37e8ea4e10bddfa7590f68c9c4e36acfcdaa49c0e81620756d5550;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7254f9ba93c8f015e0af6bef3d2cc49be409a148f793fd1dd2f6d53f29d8610e82b26e90e65fedf6564fd081ed09cd1cc7adcc1d36d1368a98b72621ef100187ded57101e31784ae26c447fe0b1bb4cd68823ec120595f33a614bd63bf3aa6f1c9e092325ef5e6bcd89cbb34f6705c42404beb2613052af2c02206f9a3c2980;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6b4e22fc9225daa6767c176524067e6d3110ca4d49c25a2fd194898f302801cd0819f8fd2292558f7e124d1a4934150ceab86d88c485a410d8631bb43c23432589462d0c1b51e1597a551232e7254cc42d8816823296ecc24088ab4faf5a85f695a03f40200e08d6ad6a3d98dbef6e915aa03a20f65acc8c5987de4c3af94a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86d9b6e66cf6c03cb2080d65b228f16d0b47b8e7a027d640a07eb8c74543467cf9e1198577b4a219fe5095216b6939bc1a21016cddb0ae37fde867221475688a330bc31ddf2034cc62b82b4f27fa9d5201752b2d273179c369400e16f00f3045dfa1d7f12fab83f66c09c71d6028b3212be133c6db473c2298f7c7198a985ec5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heba8d09cecc9cdac7ff67f06ab2e345e76840964209471470ea076712af53c5cf42a468da68ebde9f020d7faac6d9dc347ba5587206cc877c837d427b12f4e3c6d88514e927c8c0392b287d99353fc68a295471995fbe37444c32e4745ee08f68a8c863977a786efff1e9ef1b21cf99818341e2db328c3e7baa7c2290364dec5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6f75283c57bd03db2efe94391e95396e08e21fbb48b7b028a0572202f8003cd351cd5b3ea97fb12e0a68d65602b01cee8186927f8d53e9e255b0d318aec6d6aa74c984e245ffdb7b8bd5ebb9980e39a5e0231b6589831afdae159837f41e47a9fa614ca852d379380d184a675af05947f596ab181a827edb279ae4a91ff96e70;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdf6049c3651145a7655dfdaeace5b55baac262aaa78fab6e6d8e163303173fc4076eb131b8a8dc31deff474b12a4c1faa834b44f6d457a268da81c92ba5d60d54d9fffc9665963def94cdf0c921b0f99cc3b278bedc2fc3d8b2c83b975ec40003af2e688d46bf411ce1b5dc3f95177a2ccb2d05bc8d037dbea536a420f4bd333;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24811e3156cd14e0c91899193877be7647f5e460c6d3bb59264f52082b79be66319f1c4ea4b949b49834b01257a3efadec83d1ca3e5d5f304008b14c703a101d4e76eb0ccdbe7110fb57d1c02f74bb8c51ae709d34094f5095f815b4bca6f32fb45cbff37fdf03b5eb2bd20f83cdbba5f54e9aabbe5182af83cb380d57f51106;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c375005cff7aba0626d52b5a90673035d539b0dd1cd2903e72252c2a34feeadb75505878adf953543066d1bd4898f4c12c5359e4b44631d53884de3ffdadb2a34804674e60e5720461953b98323521ffbfe0fdf1d235dbb9e09723e45c244a76299d8f9bb75bf13489be0df46c9809400bfe7c540ecce73048d06575a70add4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a912717df6e299aa55e7c1cb2f5875d3550c9b9296efa1437431d83006373700ab7486f7fa1700ffb2d2bcb7467683dc5c14d8db480c62b97b4312bedaa253859233d058d08650b071c1673c467ee353c32f5b9ffeeaaf805b86c94e6d3c5487070b4153e905882f7a131a2dc19351ba78ff3b2d286f22bc72945a0c5e62c19;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h634f653014430b299f82c6e39d60d618dbbeb71db1b5b2ef8fa39d4359b50828aa65d38d543de6c8d99e0a46cd303f6c7ef5e11ebaa0c97ba900613bca9e7badcce9f40e42ba08ee250dba17ef427e3dac16192078f2ac725d7613c8a3327f09d905ab11de25559bcd176a1555a8f411fcb352c9b8ee9b21e6fa13c67c7a404e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71a833d97067d401144d66d8a33b31da0edc4ac8b300222e87799c8ec3e546a674e2a41b83036048891b9053e33e87818afd5e26b54709d3874b37d6e152bc40d4f757a282e4884ef85a559881110762c25ad8311a9a5616531a8c8071f081bfdb361cdfd0aebf4950cbbfff1c5cce5181d5d69e7a7f20df999d9f6d0d3862ab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc22d9134bcc7377a34bcaf48bad5216b130e766d30d68141be944046c06c6253f936ecaad377f209379f38c02222cd979efb0341740d87d59852c4046955058fd66b5d4ef13b8409c57126eaeb37c142cadb2e02f894ea98ea7a6e0ff07baa379af5f26712b31fea037e51e1907b593d64640e11fdbc1325c36d05fc9f92dca8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d9b528496206387d63f0c988e953d1247210fc1a51a76354c8c50157c4735a6863f6c02a2e2fdaa8df179604fca003f732ff3b1bdc9d93f9546d7059b1b5782bf7756300c997d0d3f1e1d84c982c2ebc44e354d60f75697324158043757851bf5b93451e30562f33e1f033a2633f108a998569bce7533a192d74b1204c0bdf2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27bd25d8bc1a9b1cb94f723e6a5bbbbaa1c298426bc04b10f3adf53c58360776e87a191dcc5d33d883de0e1862b3a1d3b0db42ff57c61bb6c08614b01fcede4e817e68902eded38d6c8078027dfaa2f05c28ff8aac1fc93388f6f4cf13ae0134e133b069a9c00d013882619ca9066a1af5665ce15d95da5165a61a7628e5796;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e3deff10ffce81c2732b71bf30ef4d624b2d84148af5e842abfed530ef42b95da38a9ae8e7b7a216b0c8b4be0c09d95d6a8ee4456149947c954a6ce5daec4eeb8a717b64e3eb1197a2bdfe8cefe35bc9b6419e9b016b89826b23ae41f4acc9ff8323158bc06791555c21634ce0952e22bd146c52ce9725bb83353e148441693;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78af0fbf49f16b8f6721ca21fe931ebba99c336d7e1311ea50b3e90bb5f32ce232bd207faaed1396ae8c8c1c4f39940ca9402a2d4453f2619d8f5b9378139f8145095e2af0f90839ad30ab8cb0158d313bdeb045a4dff70477126515be2caafa2d8bfd3a980009d174052a5e66a7c8d55d4308f9de95d6c3e5b05be42cd39ca5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h97c7d670d210d4eb6a330fd8526ecb12d4b307b1c172df9e207ff5f25494581bf9aa6a1584f9d822452cf532359de5399b7a4618ec79694290a6d93a36d8c0ea0f87eaa38535d971cd238b326db4c5edbe6a7b83a315dd763ff61c9b81893519ef1ac796a028af0475c363d207b5718bfef32896db1d1939cc4d09095b94f25e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he047eebcbf9ed63d852c4b0709246d1415964c7e3cf3cf291b0cc4de682a5e5164ba4926726766e1f4ef0b8f5a2329967f4551f3f47c8cbc15cc0409ff4fe7f67f09ac375438fed1a7a3a5869f0999825092006868dd801e53c7b314377e9b072d5132b5820e226e20883ca646bb8db7b802476e0c505ba94d915309773d9e76;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h75c8fa52cbaf819b5daf113d2fa62fc7e017b2492cd9e5c55374a5d75a7b0dc04b4fefb3a2de79a0bd4c67103d789bed263ec5f081b3303ab361ba316a646253b8ec00deb11726990c16b059d7ae19818673fa2271cdbd18c0d81e1411792e90d9f3f9803493c7a48ca5366467edac5ae9a2dc1d5a04ddff32aa8323d8aa1e3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h32595c4ce10edce3c08ed93c8583af6a3064270c9fcbaa68e3d2cb727258dd7cccec40f6d3f9e6a6346a1930a95bdd94167d5c524b426a791c741b24b34b677259cbdbfab693ba0b5ee26a6f01d8a33a3aac39cb327cf12e40abd7697693d0f86e7b7f9ee68f5239389e5e138c1b1cbdf8b4b8073f2dbebb3c9c0813192e4f1c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6879577eca77195f54e5fab4b3fcdb2ab4c32d692cbe8fa5e56ae5642a8664b1e3b1236119a391cd5a368c9b1594a9e3446d9c7684e584ec5419f442725f069ee41aa01bffa34440c68b2c918b88c1c144f49b2845f33f343f5f111e8d0481f4682c060d8eda7786b401b21e102875979a4e29f93cb1a9b901abf98e82f1e37;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2bc3bd685c4fabf90ec037d85086a475607378c82c331cae719a972a517949a7613fd723963db06c2901517a4d68da979557ca243bf7872e769d2dd843e0d01f58575faab12ae6eb2f64002a0e0b1bd006866ac506f1d818fc9264cd4bae8f6e40dfab7422a283eb860d8cf94a49d1e8f782b0ee19ce7e03036c3cf829ea4b61;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hafe4d8cd8bdf4516283072a7913398cf4d77b43b65c2b920e5ea879d53fa512fa6e3f0612e60f89b521e504cba04974f88e9710795c43e03656d643df2f1406d99e7a64a853bb52d4aedf56e6dc9ede15fef73dc5ff56b81de27c867725f2fe39d5e521f8f8c045a531dd8dbad889ba1e248e3f5698cd7ccc580ec604575492c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb0cb6f96aa58f42d4a73d7ba65496af504d7eddfe7395e68921022eb9b9922803d475181a24dcaaf69c2ae7fbba60a7bb167afe671e8752d07b06eee97bc9280a0c7d8e9fbd52cae0db0b7b70dcca8dfe68ac058f0926e0218517011db0eea4219a18f151d0548c67a86bd7991fab8903aa5db058c217cdc4e78f6801b370df1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd466153e70f4de0d124ffe20947ed8246619d0568eaace885f27ea47379b5aca0c4d2eeaf92149b6f088fbfbaa70e4b5f349521497e281bca85a66386a285caf1d25078cac41fc6fc1439afb1cb5a9cfc07a6373715a35ab92d011e367b5c4e993ec85ba7f146096775afeeb87de1e545987e6d6faa4d8a1182842dd030fd1f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h77c5c6dd285b88cb43bc9b14eb8ea84e0297fbd094e74cb1e78415c092ae135e1e6655611f5f8744fde3f8fb932d2bc0197be553ffeb9e1580599a6c08d2bff52299dd01617d06532a0edabde35a5d7878f460ce2c78c8ef7ffcc4269a4df585e01e66d1b926e35818c75f4ec74e71745e85c2dcdb783018652fb68f571b3914;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haff6f570376cb2c91b49957688831375eaacdfe526b19ab56d2f5bd7a1a8182148cf909c28ff6b6d188d652129064a5d0ab3dfb8dd2c7fbf6ad468695bcef76e5ee58624266d45baba09de96956cb86c2c170044d9751fff45a707f7d536d9fdde9d7a1037cfb0c33a0b0f48b0aadc9a69a15b6f30b8e1e51e21317dc386d0c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b0d9323bb5f27068c00c10071554d349bcddca3c0b57e473c0cf01628d4616a60c1dca6e430fdd19a992c576588cc86c1d54783881c8018a30a9fff293c92a63194934a096360bac88b4e9212df0da40b721b30e3f1abffc2d8a112a4d7b84fa83674da9aff9994e5f7d9039e3218911b553a46abf314cf97a69fbdb04eb940;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h708729c1ca968b05543e41195ee22621287f353a90c8fc2de6d6b93e123398cd7d020a730468bf56ea7e3a64123409d16a108cadbe10dc441a4b40475f5f19718563cb0fdec104c6a1cddc7c3c0e9ee308b5f9bd72a53d628dc1b8902ffa95ef59f33e09a381e68b505bceae9ff67345ab1bfd9b6c8a9555d94cd274e090acf5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40cb3e7f3535b23dce3b7cf485e00053358ea8297fa3cc2a2fe7cd98e8fe6f54dcecc84419ebde004424c93ec478bfd894f2013d126f1b502f4f177a73918c796b918b585cef495d0a359f357ad84973eac56bff7aef14622925c2d03f84406252b47d41d1dc2ab5e94c7e2dccae823f960735e8c40aaf88b9eb17859143ec85;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h867d40d46783dc332e15c8c340d96cee382329738590ed971ba212152799d29891d299d6095971577a8143ea3149d5a1b5c6a251c9bce2dab833b625e6040d8b1e7e5d16809f115d3a16769cf81b66035df90d3df9e3b46ffa34d72f71f4b263f188ca403dd333bc708105cc69f995fcc202616398bf92683131860d6a13c4af;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h93a168a7adac808ff900c70691a75d2e3fb43939af6f3ded2b9eeb9a8b6184d431277c7a61bc9f7a067712bed57d9b1b36af0ef0e7f17977153468afa2ae6bdfb4acb4864f45ef48a32a0aa3107edf5267c1b228d85bcae963a70c75c9f45d97753d4fc86dced358260a73cac8710afc8e474fb3319d40e9d39ec5f3a22ba4f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haf664571862a2b378c77ebbc1f85ce92db0aa50367fbf05fc37f4b49f7e4dce11dd11a1550a394ec27c60b62ec9dfbc5e87488a262e75be5e0b62d18f8ac835ac9c66a9a3d3f0b5428c3aa0e6322a3715cd376b4b608f56087899eaaa7b7440c2f24c991f1a006e246a702843d92ac3a19aebd865add7fb535a69a3d9508d8e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha453567250a2d482e810fe17c89d7f7ae678fb82a07c0f6b89811483ce7290df95ca4681939df00cce15aa416b1ceedce447db6a0be0a7993acabaf2725ec9fd9ef40bc5dbf35ec0723551655fbfff118a57b005e095f26156ee5af7935c8feacf19a1d6feda4697c8b2ebd9248444c762ba85bbe042b8242154c19688c66e3e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1f644ef0bb6967a314a4fb87aab4a53b74b767075019dfdebda1d3f7e00f9551a2fa37a6120fddce4f10483ef54aab37ff65f49e9f3f74afec66c3da05f057a56e21ebdde975835037fbfb0ea8c16e92d68c27073e3b6eb19bbeb42fedf8d81fda5238745ecc2c07c96473a17e6905499c04a9b7012d84b83b06ba86a888967;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7e66541c4156518145d66735534b993014aa04b40106aebab2a2ba7dca4d802a470a1783526a4aa908d6ed0c960e97e9dc85540a650643ee43306319c239992e2239a951e40a0a0a9068d09b1918c639c6bcc738b60604eea8d49744c2836cc1d7a09b9351a4fe2a56e2400009dd498c21c0ea96ea6b6f6c7f615ba71a64040;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h130606741643f95dfe55055acffc9bd8d1f3535b26ad6816a638c0f14109a5ce819a24b5451a853a0804cfb06b0fc7ad3b50756a3755e67d14d76ad131b85fc1e860db30cf365676b8c8eb9d3baacfab29c3f2657a2cdd89540064ac7943817b5f826480e97c542f19d7cadc1cd7a558e60e25817ac0d01ec289b532b14ddfe7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2565403014f3bd269461d9d90b2e843975c1ee3c5830158db109d7081202817c7dd1f47c25b1a2169102474c09fb58691922f557258ca3cfba4c9a1319fbb336561a07b7c436d0a28bae9912445a157dc0537b8016110449c294e4b44a4599ff2406aedc66f8cf5a3ea554c8754497e766141032982cea60f5648af988c46234;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h71b9ada4a54ec9d2e5581340fb81abe784922f6fd5a1d4b44211b508d78a90f47398cd004c92a469d8135ddfe334be64e2705f473a82ee570fa0c403c5cb9992c933caf59a642d2013fb288fc4c0dd091d4874b529299d315783b020d98c14daf6fafe0668a5cf5609874fe57edcabb90467c737aa25c44bb2fdddfa5335486f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5dc0944c14f84748784098b539c918f589bd4c774c7b5913da9e32962b53ab197e34f2fa7a74a8b0501f8f287aa69d039bcb67cbd72aafd5e2ae2517fd50d3b3fd155812af79a014644d3a8a7ad7d1c802268166d02e8fb4ebd033de09106a4645caf63f589f3b9718eaaf405c74880cdfa1f0a30e475afdec8c0b9fb51bfc19;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0064b1ad7c5ddc19dd63b6e64ca5f71aa69bbb18d8f187f40f94c66087aabc51a6d32adc82a764aa24c23fc893b1ef885226b75396bd2e5cfbc861a580f345936f5f201e180ecacd4b0351424c587584b1ec6d8b7d8c32abdbbdf3de9845d240be7de720f69afad79b1b08fc8e259b9ea18952aff892c6c9d3b8aa129c0f93e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8151ddbde31baedfacdc952c5e7d46ebed3e2a0131a0e0bab621cec9775e444ed20cdd60757a2e3cd673d981075ac0821aaae177a8af113cd5f740836e0f2341195e2c25feb82046ea17bbae0453fd84dd4b3d0c2c8c650a8015e81e159833f82368a65ec7580ceb660a05ec4bfa68336ece76f40ba2a4932d538bb4b774c570;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7247d676a1dbd0a6e46f4fe908697e1921166b0cbc71626d14c5c7ff3bc6657a253214320f12cfcffcb3ca03a7fad5bd218ce02a884809700ca67034bfa50b9e0eb1b9b391dce306411c00eba1afa3fdfdb9264460b82c4a75c8f7986087a46a0807b159e450f0e92faf9b59665139b476a4f6a0c458fa7e5edd108e6296d96f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcf86ed239bec93e88d46ebb8118cf511c043c3446cd899e7448ec71c70cc40243dd15a2c3d38212dead0295eeee49b8ac36e9e40a531c378b961fa3462b9c59282e0f3e62087234301dcac65a31de24f928b7cfcaa33b564c39afb066825ff793753a253210b77910c4716a803d60fc3c987373ff86969867ce4cb957e503ef7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe5fb0a7eaa1c5978bb3cb5f9bf8d119e9b8725e86c0d89b76be51ed2d18d723f7f809bbf981800be36af3fc0718a67c5f66e8a19957e0448d9abe40b2abba4a5e88d877449c4d6b1c38751e7e06e4114876c650f6ef45d1dcddcfc62bdcb7c9d77e9411bcb07c02d007f52cf6d8426c5c6840d25b78572c47c3e872b1587441;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1efa6624510c1d41da8c58df52ddde8bcc842840d81a8eae9dc0214e50093433eb5dc00dfa8254615c0ef7cbee82d8bd8fffd31e774d74a2877947cb9c32a089088c42ea0ac494034a262384e4433f5ee244b8f7703132bcb7cf5f1d9f0821d1b2b5d273827bc66d52472090a4423900e85348324e7da944c45a3714af9c5862;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a1f519ecb8c226d06c7bd44e1fcde7b724a9c5790bb177e073faf5f3b5321aae3ad1e4006eabdcf90a7a1e77476538f7f1e321e0a15ce48a21bf0ff24c88372e6796c2731335ae0fd77719677e71c020dce0c5412a452dd8ae3dca2148a76a7db0189e46bfb16e3e5db86c46772325e2b99a9be73f863f5c662ea341662f19b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b00a5ad606e746b4803bca0ff663cf936cf2eb725aad5e4b3ebba377fb9cfbf6b0356cc5edce5d99905484404d6908c46ce07b613b13b7aa683b47dc4f735a8e02a56c88e990d314edb107642fea75c3613e54dabf3bc6e583a7738ec83b05effc95cc10462c4bddbdd5c8b81becff1f2b1657b3f15625cdd7aeb0a4db68e02;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe5fa842809b7c5ae29ab64d73e1f419a84ff7777163732eb761246fd1f099c43a2da5df13d51331c998e55d00929160019d25f3cf87f53e89ffd0d6e39642b0d00709edc69097926ca91ccd256d46089da77d90a12128ee90851d6bc5dd47ab1204700b2230bf1ae9bc429c717de2090a24ccdb2be94455da4bb80e62cec1b3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heeff238719c0ad328703d299c7b06ac984af12aab0b119454753cd902d6ba7f20b43ad320f4976e895d4d2eeec8e9b8f827401f4df73b37d02f5baa47a75daa25c6b05f3cd8fe989160d80e0e00abbd68e774f5775c433622c94ce6d6f44cb50a454e8f05b98031f612088b4d125dbf6fdb5dcd9d8f68be597109abce57a073e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcdc4bb93523beb1df982a8676fac8f162ab8f0544545ba3dae162386797080a5a15abd6858cfc52d0c8adc10bd84c315b837b16e547e9c1e2a91c5f28232a3f7da40be9f81409841416d430595c8a8ba457842a98c0df450152e94eb76a3c228368cbfa2b880f05ee7037b16c767563916c36f777b1b42d72cdff30e14c45f38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd779ea2534803e079b4630b07ed480d080f54980f103e90b06ce720030feb7a4a642f8986ce3a2e8c9636dc50580cd6cd9de6e0537e78a57c197e88c5347322cf4155f0d59ed08a4b621b41ad0d522cfa2629722dff05546697c5795dc49468874b3ea7835470252d5e7a4f09261099ce6279580172eddcf5061012d382b6da6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8c8cbfad505294643020ca655c8c763ac2295308c7f475976cb522abe507a5d415abab10bf71d177ad0d6a5c0e61af406801274298a6d5834e85e9addc728ca8c255ccf9f569288a0aadc2da17f02f8892c624c158e5832f1d8292d014f1a75fb4673b1bbdcf34dcb14b89ffa43deb99cf16a489cf72b3f579fd44a173ebc01b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8becdacf79d6cf4d40e7f2c86beaa6ad60c5cf3220b9c9f420b3e21f1216b441d4b3b635c5ba1a63a623b21db9ce6e08a83194d7c309cc2dd09a9a611382944d5446d9ff6146bc038587c848fdc6cadd4cd2725dc95e923edde536ae4744595d687d250e658679c65d699b0af78d4cdb40e6343b356ced4579134f47b643006b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc34c20afab1571adccf1bc87bbb71e1229f59c5b677fcf8ae3ccf98bb4601441771bbe0951216e3d36659ff33b81d602351d76b05a1e2bc5f180bed79e6745871caa5d1fc88c3b05abf501a1a2fdd4fdc94a50093a92af0eed92a6ac0cc42bc4d3ed76b2eefe061d3158fb52726121c1c9f6e60972d987ab910219404f02af1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbd55e1f62968d73cbfdbd2bf85a940707232251d9aefbe56523d84984685b67717becd6b3cf407f4767b41413e30a9ba9d5877c55b23a789d561f72f716149759cd78e52560ce135b481b868c73aff1b2fe4a9f1497499502e8215f91d3eddc32721d58d62428083af883a93f710f358df1a40e9c49688f1b97d17d3f5d6a0df;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1b42624953ba9035d57326ea33dabe213c3c36e325aa1b3cda731f56e021d74829b2e5e32120c76505a3176cb9e11a3f64ba0825604affb509adcb7891966f10c3bcbbe70abb83b3ca33621b92976f1c2aebd3877ef4e911c83230b1319e01be85fcfb2c4dca057af6619a38cab9736738b0e62559cec67c1ca7f1f9a8c0806;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda75ec697bf30fc10d343f7fe90e0e2bf8565addaed5d230916bd8d41d822038ef57109287203b35e41f6afadb337931ae8d04835cafbc5fa1a98e699f28ac339cbfcbe7c609d3f55e6c0046f04457a9f282bf9c890fd1fdd6f4659cda7257077a9b2aa59ef53bc16201d6bb7b032d2332b6501caabeb04951852baeca89c024;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37fcf824e83d46858dbdfde2602f15258001a2e49cf428fc8bdf84f09551a66b9c03c1d06f11209ad0eb1936853fe14f90d7cfea33c1c5b5b85191265d581f7aa03dd5332cbf1e543be8368cdcaa5561e87a644b13ada6e2508a88a45e48ca76e76ecf8babdf58773f4e0763b407d1e0b0c32798793d1e971d2249c819eff705;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e953839d8230a910629442dd8c3cdbca6dc8e3f7abfd47b9d597d2b05afaa3b954fdaea92c72ea7f76ba17e314dad345b32c9feb28ba427023539ee367aa3ac2c8d7c01550e91b68e0034b5f6fce1d426528820babc5a8983d34e8caa5cefb3bd8c4c20cc8bbc299cda97e133c66e78156966ee0151b1105950371519fb51f8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6ceb98d4800a9844da689ae9ae1a15b0193d91ede9d8f56031545286b1798d48744f14352b78700932d2337ffee86f05a45d879fa0c83c8c51f540f0b33a85c6573843f9b179e2a4d704acf501a660ca4531d1eeaac504ed4df75cb066b26cf6e935b86d91826df24e4d6dc134768294a357782630bfbe75abf42812caec4c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9706baffef3fbf04730a574947c904fa76aecdb016b5f5d3be9fac2f3cb23fa3efdf4fa13d9a1a43c24abd4d6620a3684dc7bfa704e7cd1626d2705fcade8dd53eca15322cf68fe141b466441d93655ba0314d6e6ed9db9aad46843f66477e88365723f3ccc4b923dc783a7c25a2125a4f5ad0fa049ab08fcd53ee5d0605cb4a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfc37b3403fbe2d69d5a599337a9628cd4976b21a1c83bd9dceb302a0f953e3fa7575f4216203eaf5e40a089e85cb796a00ed77b957dd708ebdeb7a8ba844d53b77a3a082908469586d221064f8a9d11873dfbc54965fc37dd47d656b09f27228297b53f76fc5a95d8728b543223d3b1e73519a4463c27247f2beabec809f79d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h515b91d57911bcb487fe99e226747af0be24fb58cef89adc9f9a4771422554cfa26214c9d26077bae80a85a1958572e78197fd15359b3a13687975baf5c6988915890752b14f113d79d6d1e8291d2ea53b75cc8f1e475d526b6d5d50ad81fea67e2a7e4872348eb3d2d20d2589232dc3d1f80aebd16f96a6de9340351c243b4f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3988d50099bfa6d3080c4240c212415d6a84331728b9b6d2d57fb237fd171fd9a127a11f046d955b75429ca859a497804c7bc03ddbf2b92374d123ed929faf82077a9376104205c41db93a1a01dc59848afa66527cc7922241aca71380b244775e6cb4eed192c858ccd3157d1ea7891d726b49ca78cf0bf36428cdb8b2186234;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74c3a1069df5b2d4f1dfe258d92550bb482a7028a4646a90488bbb768f4443054831c51c1f49a266a8fe982208674965f663f34be7cc73b942bb28bbc531e9f32a460c2ea167f915461ec8d12d79120ae751f3ccd8a54e5d313286c3e7765cda177b5488d9cbdb2983031652173af601f5da93bd4aa3979d880598dbb82445ab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb1c3a477f37c37caee7197b09d687b5c44d9c05f83578bad47ff1c930466361c88dfa561d342d4bda4c24e50ab95dd3130cf881a82fd0b77a5edcb4fe16a9506981ee6710379e0bf94ba88428cfb747730c9488aa7dde8063b6dcf38a2acf058098566fe2ab3fed2f45f45ee7868b3bf1a4675ca243edf826f77135fb1d219a9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b76f7533fb8cc04970f86bcf260fb41839434be6d41709cebd68d6367015ca716de2b5edb7bc23088bf9559f14fc0ea22bdc7d0bc69dc1e2ed5dc03a3cdb92aefc39d94e38340627e329e589fb81fd005ec8bd7aa9d0a9d9eb2f39c68ea69cc37a4d1345ebeab93dfd4a7da8d3453799aef398f783408d2eae0ea464715444d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9394065c9d0b24fb3d7fbe7a2348d70ea245e86679392aa63ce28b70d52bf4d9e1cedd4f483f48be0344622e2e82a586b79f5fd4067991a8a3c1d9f58303dd2c027f162a3d3d8bdd550bda9f8e30c164f96aa2af7e421fe6c69bb54d769b25cae90c27f70ca55186eae347f93590528910d0ca2b9a137b4bcf3f57d1bd610bb8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h776f7996b9d4d24e91a8f1b743616b22bf24de43cba9151898f1a0957928da3319ad91e8415eecf23c311e2a3d1f1466309e998131e5d186c4bd3f45b5f09047915f0fefd8b71952df57a32a6b7f1e05113b81c364806784d16c6a8374bc3761a1a3511c7642c7c5c85948eea0ca170bd7e313d5f35dd431fde5448f33e3c28b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8ed3db001f71665d2ae1a25a5c57ff255b0d73df9c3986154dedf984d125e3afaefa99b5a4b6cc0691d3deca404efa7dff2842f22c806117a76980fcbe0de0eac41493cd6194d5dcdf6eafa381ba2f62f97cbc2ace1e1c0a168bcd8c7162fd70799ec599bff88eca8eb3ae91a9344a27d9f8e93c60cde19dc4c03e927ff8d63;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc4d5a89b95103bccdf190d2a99e98a0b3d5b42699415254e8cec2d74bbad4d544225a6f3f1d5405d7d3fa1f5b1d1cead1291e15fc4eb28d6cb49dcbf83cae6a8b640b58dce582d50fda799deab09d6552307c72c8936ca9d94f57767dc30382c60313f1a2802bf2cca806aaa96573bc1a371018d98d69a6a7e86a87eec3ac099;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae2994f5ce55390b16d65770f97e3b75f117b582dea0b35aa8d7c78d7df9b86a2f42319f88ec18a6bbaa8ba0e08dc4e42a50df5473fe54ad82b421fb2750911ef858eec849105daf7a6f2f384cecce732e9d2218d6d5b79867a4a52ea88c1ade031979f7ddebe279d44da903e3896af1ebfbc6e1147f10f7a9953fd00886d080;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h42a07c3505b7b5278ef74c946722777b33260155f3d253a4c5baffbf16b11dfde9a1b5d63bc26c006108a2fbe757d128b4a38ce398f497e6d41c75db02501151195c762f5c7764f2b6d48bbf14a3e5d9295d9d2d0a36eb1a0e87c909bb37b750e808596988519691612670045cdc705be5c2000e41ff510ccb527ceda438aee3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9428eb05018a67eb3f98e0bed9dde166309f5d73642aaeb4e77ab8858ef8bebf95610956113c041dd768ccb2f8d174e71e9e0d9d4a0b2a71c7b0f6d5ac5e9bc82233b9b622753120b971baa2852cf2616a900019b358f3e4722f1a9ea2c660f76f1c1771406818bcf04936434c44c0acc5c299ec7c14680770df3cfd8add0b67;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h99c32a7210cfd259fe516f5b640df7af81aba300d0e78f78867b3606c0f1d5e236ae5ee9cdbe6ef48f9e2becae2a6cf99bd09c5e5c3560353035e1e48121d77d40c4011465dc14f51bfa6e42fda9614c1ea3d9054dbc7e85a2d2f47d6408f2ac485d22099436fd05c2be336f16a7715e4d9a00c23febbcca60312e8f849374d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc286e919ad22cf6aa35029b4e999717f176a09bc0aabeb692393d999051eaa02b0e1e04cb53716678884238025f47a528569b253192afb2c02eb9cbbc6d6892280e5df9e9ea318b57710351ee33408f2907e7d981da7b4935750dcbf33bae36b578afb743b4b42d05457c2a89430224c2879a318ab8a55b579dc38a1a6eb8ce0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7ebb3d66e2b38b35411b862fbb9d7f0f12d605cb6812c6927e4b9c628c54b013e6a92f283dfc61bdfce2694ef1b5955eeb4f771d1c21ff6eb663e99e90f891dbc7c6480c427b07ff348555dc64223fb0eae0e68ddeb8ce5e2bd445a3f5634c0a61d30a11c53877254feb2ef98a01a45e6b7ed498af57187ceb7fbdc49eb6a84;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hca18e95bb10d9b4ec43b9766399280bfdc945803b170a8374d194b0df0e8a26c97853e7190a8bc7936df606432ca043d2a6eb406549b400b29bc820edf776bcd6f72819d8a55f4461cdde2f928dbc9342ce97ce9b9f5b5f9dcd317377c154dd4babe711c26a0c189326254a2538244ae5db1c766f1908fe49ec5b79fa5d196b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf68801d06bfe761ba02a0cd8778e12eb57bdc4fbccf081ed2dce301df74910050a60896381a87bcedf848c86880af833ba40e73051a8fce08110819551ff85033a7a0a7a550375976ead4b759a5e48a95225205799c94a53f4d21ef484958c962f3c4265a3306bdbab241956fd9f20b2b41ac936ea4eca6c5841c9a996cd666d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f3d17fe02254725c54e11bec9434445be45dda3b69121d96da61279daece094f7d07ff54e4477f4845672845f66aaf61d1c5d9272274c71bc8fcd991e70556a86a8434b279b02dff07623629f8936580df4f4e590e74ee51056b301a2061428ce2955b61bfefd085a0c02920cd3a2f8f840f13de1f3ab8c5d7b49428b0c8484;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h371db74a596d4375e84fac74b58a1b6a5805dbc69c1f6779ca18f88ddf19edc926319078f8bae69690b9466b2d3c64c0b92231f299796fd4babd3d0caa1158e060b0db0c6d1c53c5ce83a4b986b6d3c727e85dde19897cbc5beef683ccab77abfac8e3bd8c22d2815b4a0e2923597973f730ab2b725287d634569991ca2eb95b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6146ee3c5d352288a7cff2500ad5835be370e2e92fc5adb0f24412de7776fc057991acbe5687c4d8bc1ab209750788fe0ae7231d8ced75e749912d562e3e388011d94df38701102e99a4479fc4612c8fc857c784f15669fc9338f2dc109b8620407066b68c92ab47f413d3909216d5f194eff0ad538659bd8e341574097fa275;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hef9ce0749a2e298ee6d344dc94e47f43223c495a0d5ac8f786fc54bf69b7b25cd1b0038dc7afea6407db2d4a56e70434ab408d9b6e37e690c9fd85433b66d40545b3650468767dbaca7efc326283e43c53341eb82f46ab628338a439b740c6609c7d58f425ec4894438437dff50c3f54d8cc11db1e64e79d3d134199948aa268;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ccf5cd28cbd60c655c26bb1d4d601128ea42e8b1355634f29c7447c0b95c36085b0ac1c00f33ba51a568d2c16d5b5c1df56a23434d6260ec408860c921f3d97cada992a4f9b3505972f956a28424dfb3a8fcd71aa730e4e6eb62ff3ef99bb0edbe787fb960cd4b101726328625ccb091dcfab5aed54ee6e31b723021f9e3b41;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3f7e87f1c1d2f187f2d56091fdcaf0e34d29e6a402ae7d5ceb805721fd40f866bd57f4fd580334201260078fbc85331057295b7458b5ce24da996ff8f9bcfccf0e1dc46d052850b7aa00193bbafa17b682e66c1d6fdb982e7bd21da3d792d2dd0d8de6cdba4dabc68703757ae46bdfead3f4ce7ed912fbfc99f29baf5fcbff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h842a0f76091853c3303b74b44cca23151c0218479784b4b35ef52d8b590cc9c6807229078b14dacccb1f5660bfb02c1ae528d9c48b2d229fc3cde86b44f451267452e3fdc3196c45eff8fc5b490d2ca59d7b68a06bd741ffb201c5a332141e4fb008a1311653f0c560f760b0f7c55414af0417887cb5ac9df4f71ee918c5f261;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4ce9ffce86642f6a08addfcdbff2f1d4423b1578476c22086ab0eb09dabb9f014497aad5cb6d34fde8aee6f5b1d9b889cd828b4dd1638afebb80908e2fc1cd477edbf514c40ac541a2a8129f52e3109bce1a4ece93c565eb6aaa63828bbb3eade7d5d5e3609ff7bc949c71ee375ca39e6b1ab29b903492cf198be21c8e39b6e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb6314841eb81b6136c9df3ee3bc4ffe45c7c665e5a2aaa8f8cc159879fae8dbf1b2d6acdbd85b364247895daa92293240f8c2674119e3af4c7261d00fa162e317fbe6c7e834d64ff0ef2bc7a8713b04fc6da8f755f4fc898cde91634d85727a802a880e5685a402f6fcdfaab4d5edd480bc4fc18ac752fd007aec4b36557d7fd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8a81f4b17d26686a63d482706df06b11bd4bd7ac82c2a257ca3192319d13950719e7335496dc547055b458ce7d4b5314d6f2eb0af3b445de620d61a7c7f35fe6d6b09d4fa5e7bfcbeb71bf77314e0f2bdaa352e4596d168cddc5b8aa59b59fc170f17e84c0d51b23888b329e75030487dc489a48063f112386a10105e3a7612;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbbc854bf2c2ae20f9562bde62e0f08f3f75c01ebd2bc907823fee8f7a74b03009142bbbb20da81681f0df09476336342738569d57c7eab852ebac6cdc810ac41a3e13128a06ed1edb0cb72b6fec8845dba98077bc231bdd93319e7ae34d68a8840a2a7889c32a5b4195fbd63c7e480a068c03dda85fefde1e41769f6c16d67b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8de09ac863d0257c9aa7b29119af1916d132ea71c9416ff29b18954be71d366bed35a7b7fcc9c2b629937c6e0990e26d08235a50debd453f4e094c4a4d3d8901d8cac0c9b5d395eeba560060418c55103cc2f76c703f5ad125b0287661558e7ebb05c2f72ed3a7bf038ad2fe159ac30721a7b3d74e56b52fccc02b3c7d4e693;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb707128c037d1103eaec366cc26ed6ed1553e26fef7629fee9dfa49f8397ce57b076278274abeb12171df00afff1dd6a80799bb0980e21da52102049ea1292efca38180d1af23b5e5cd788e1e8628e44250bbac562b0ef5827754d495453365feb7faa64b1ac4279152c8da2d21ac406a524c5c557265bdd3a5d335e3f661feb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd061041c47af1ac71862cb63ef0e48d76cf2afe398d9dee25796f4c7d8e27da2597f088093fa5000781b269a6cfbe177faf390fade9cb2b3fd05bc3d29ed0aa4c4760ae02d45206c12975b9e880181a799aeeef5c29cd9ed98cf732751ed7b3a06807d9ce7bde3ea2bbdedde876594003f461aa37adba7136e30946680a9f16b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab23f017f1103f51036d86f67dd942506131091076a9461037b2b0ffc88ab82ed99a873f7b06f6bec94372d1ae7c2fe094267fb3c27b3be96ce0fc747d87d9674f6cc800879141c62f5c7d9761c5121e670f0dc3fd81a3971a9d964704d2490fb85017ccbaad267a326a0e226078557f6121a67ec7f48c82992c2aaa100762c2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha54c6e85176fdbc9e49cc853da5aaa63a1ca9982abab923a609689b6d23212596704dc45471eb8fd2c3b8143a8a732da708de45a74e5026275150a68a8726abdf3a6f70df23bea795e82fe624ffdc64da65479f5ebe9e6088a3b5789265b7946411f0e0fe93dae3189db312a710b0edb039c996aacef489f547ec1b2c2bd9196;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haeec53d9d7cd87e8fc34f90618c9e56e10547db4b6fc46f991a424527951d8147717339b2a857d5b39765044d1c32ebbe4752e1085b5d451d132af9b6477792abda16757e5a302d0edeb2de28f07da7a7148e20b35d77b4a15672013f7784e4fbaad09b3d447a46605a33c7205c9be5afcd69246a339b4f3884244765d6f2a86;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha45af34c93344775d621b6b089ba15e26e061397f209ba3ec88b715e0ed2230b64eb992aadd769d041f59e0969506ec6a79f7c61bb6ff4b41197e607b08ca3e63ab0f5601f745ad2d64d6a2c107f8df7f8a627f3597f4952a6e99df6c9b62910c433f6dfe38f6999070c436ff9e52e33717f503c422739a5206bc7e3a2b9599;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36ebbd5f912e01188a6fb8f910b3263a6e497f7efe6bd1665cd7cd12217a52b4b5944b5603e74d89b1e65e1761215cba69b74a8e78af72d3e8d51f83f91a3cc0509fe1a279a0c25880a3422ff528080b042adc15aa7baa61ec4cec42f1304869ad41ea218eb4ab08527c49690524cd642c09bca477958d36406318cd0a98d9e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2310ec8d8bb590ac4698c6d1eba78a1cca2dbd40e4dffc267d53813cbcb963661641c8c597f07aa3a0396fdc827cffd1f9bb0db2c8a6ebb792b5ca6affeca7f3d6c9b3f5bfca55dfd8749fc8ac3a442425db1d842e46d91afac2c139e6d27174e1ce3294e28668c6867c7db84dfea97e9398e894623085d31d9d8179ada330ab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h29d4d4084e9802c1a53a3f46f0c59b8bb2df13bc1868cc75e85d5a19765e99b23307a21d1080cb9f594504baa0331631f008c438ef93d9d684a4084c445beacdaad18fd32a8126d1d972ef0e83c3ee402abd9b55a3392b99327ff669a553a262fe0262371e46707daf2498fa5709fc5b2fbceb6151e5e34e2e7cc5d51bc44727;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43125e13832a6d3186e487dc26e92a45f422aca13ea0d635fae107e802314872a053c7dbe182ef5d46c8028887ae61c1042b67372754d89607fc8af34afa3591f3c280328e80c30fe701774162bbebf373aa2e4bf139bf7706c684060a60c13eccf4afb0b0ae26b5bf3324ba1e64b777998eec48e312586fb4093553199adfa1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74fb59587c9c0ee5ef266b8d928ce3e91e674adb8b410c91867efc6618ba6a529fbfb3167969806c0183a4817e0ebfee93ef1edf4242ced9220aa6ba22e7755d24f8eb4dd11ed83ecd140339e1443715de74fa58b19c244af29bbda979ad87ab8eea63b26b97c3f6e02ceb2c07db9bc24daa2a4f17803a191b623742edeb0607;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h30e75a8bfb2b2db2ca04d62a798b5b290a05f11a2a92aa4034b5f173e97a7af76f4af977c75a3ae45a7a4cd9ea272fe302e157c1bce4a97953c373526d501a963dfdf698cbe6fdf92972d4d6af613280723980c4f319a82631532b6fd6ed92b5dcb22cd678211bad5eb6c8629d6b71f8388bee3025a13be5b1a5b20634a06f08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h85f5015ffd4f2ab5f8156beef89934f96d5274c812ceefdd797f7c102848d2067f9a2451c62116e23054dcd952992cdf845bf774e1dc0edee11df773756814d389f84f104e6fdd0b414c49354b8471ffe7f6e0aaee5c18c24589f351e38c0705864c2c0f7f40615b6b30170bfe1aee59b55d9a3267d0840cb5ccd12604003753;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa20536adc4919880daffa43ffe470df5f64db3983ac4425695315731009f479dbab5611049e8b5c5f4672786a74ba571c58aff5c19a358f3f02f601ac3863b4513094a58aecdbd5128213dff21f26c69014ebab9065e6c7111c9289a3c2588e5c9d3c320ff4ec1da3d652fe84f16eef7a0a4567632bec093d74ac7b6a5fd699;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3336bd1159ea45b1223ac91ed13c2ffe81f3eab0d4a4333181b1e025cd963d56a1efeec28185c9dd63e331a6093ab6cfdc17c9a512bdf020c9573462fedade5f1ae68e3fb604863dc11cec4e0997e9b4ad6cd42a1e3b51f977868a2fe2b79f1182fe7a0887054789228dd8924863a6c00633b7e464e427bcf14a977657aeb84a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1567104da525beb7d27357dd096d72c9fc6eed17ae14f544bfc09c49e62ef6fc447f68ae0ed3763418e87e672c12495e5ddb192d16e99fca81110b9bfe20e3f17e3f02d19fc956cd0833858674e9a26c70afbb2f0b925c6c096dc928c25fb9ed9d404f84f5c07cf2352e20433c88faef69350693252087aa3695ac966a8edc3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb53199b73751b90e655a3333f04c0e8fc90914b3619f7785078c03417362c253613090ec8367a009e3ba2f93f74f508dbf7fafc598a540b3250c223da57fa3f929e8cd7d1321f908fec10a6d500eb9eeaffb519bddf55dde0b21df6b9dc766fcf77d7457a157c2eef475955772e37a2dfefa79bad11896b41d6f05f00cb91fff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b3a46b67e7b9e97cbcbbc248ed51ab90a3a14a9ca7c8087bfcc30c2cd4cbda6633bc09557af30a0335cfad9e61410cb10c479bdbb2ed6b093831d70bc382f2ea9685fc6919fd7f9030f5d17582101e712ff26adfcca394c7be3afb1d2a573a0a02f51df9e86179c0e9c27740276045dc7aaa4bc2aa69a2a0dc275ceca1974a2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h82b3e71b673e7e7b9293249011b0102a0f37ad6e166cf8034182c046198a11e0fe4c1c7eb689ed6b855b850772079db485713fb1163b51ec36b5da362aaa6fe83e2984751d021781ed8e96689904f80bc867820be4c4b73e38038ed3cb1e150d4343ee72fd2c17251fd1ea6520200cdb0e53666c4e7d866436e8413393f89cf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd333ebd019a1842f8e0b945e3599105133d48348556f064eb416dab8841756b4d7b55aeac8cfc586a3b0fb5eb50f7ca04622299bfd9fa831ced884d90620baf1ee401ffc17f7d1b9546ba8dd20d858e32cc5c843055be7fa258e137d48c096306d00433fe30d47efab727c04e2da1f775be1a8719389478a3bc0159fe0c01c13;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha7572150186386518e515ca065d162a6dd56636e40ae4aa80137339ae2c6abfce25efec092ff0950a488ef2ece51e310970541c605ce978546529b9f7ac0334873f2506cc059010c982516d61e5765fff9529ff13e5d7677d66c1c73ce8a68d467e90a72d2500d3ba0c5fdf57de1f9499155e1105074d81f249076bbdf1d1426;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6fa61d28440396e7b0fbe51046d878061f49da97ea074fa73cdc39680bb5946d6f70d32e785939dd675b158cea3f249a0c0ee5530ae62a3c6a53f74dd5683022169f4e938f958fb7f5a95cbd22708330716b91af473a388edff9a52a9aff947452fc1594de412c7aeb189a1e1f1efe26a22b9ea18a322b1712e9648db99c0741;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h266f0c873e4c54f6ae347e522d6feb214c871127a3658886782648d4c8d89481b91acb883a9b89015ca4fda8df52b92fcbcb52323072ec1ec4b57c41c7e463bf91cf77150af06296c7c4ed7cf140d0424dd754599b3382d77a883382407ae9615690174bdf3fd98cb75d4f6aced5da3484a85011d79328756c0fc21c00d4769a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6dfd940eaeb879f7647dc33bc681d5c407e1e01eb0405b7f54cbaa9bd5ea32bf6d61c0fdda8b253b5cff3088ec1c78cf363188c53b7cf4043b3538e5f87cef73621ede60a28ec9455d3805f3a1b778b2d5b558fba159b9811564c1dad34501e7b3c187963275c39987ac7a800076ee888fbfaf0d76cb10061140bb1cf8562d3c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd94cfa950fad284aab1d629801daa0a3ce383553ac097f9dea7a2a18949c48c421a29e77a753f1fbca4b6906d5cb66cd2f1086fbc21278ae60c0ac3424b51c7185d0e143c31d8152da29453f9f042610b09ae1f39349725c1d80735e19ecbe220ea6f4abfeeeb4588debd9947c891cc699fb7bcae829c41567ed78bd2e7865ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8827b61aebd77740e861de2547c2ffc298e3547c76a5c042d9542aa73efafff0a44aa394d82e38a91d40688232114745650906da4ea3062a52700c9aaef9df985462166e184ba60bd3d5f086d92c4ec9a84affe452bc7dd7fa06d895171f21d6934c7464eb54a03151acedb73f8820db26b3ff8318130e56b5bf5a9659c96a8a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f619deae979002cba1b57f8c24f645dcdddf38e0eb295d5a9888290d0476872dad0a22f32483822fa5926d40f701e58c8550cabff219db74985b090105477ce77269e9ee75c9c89ebd9f1e6ac8e8ba4632a97200acfa84da395b806e4a0661d56b9543f7ebad3c482d4eb88f7dd66aeb531015aa7aa5b2237ccfd1dfc4839b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb28499a56188fbf2dfb36ba4544ca85ddfc11dd03fc2aa809bb171970bb2d1472a42bcbeacc45ce1a7e6e6049476c9c73a09d215c7825a98dba855e810f802bc02f4ef65ca845c401a4127edaf5e78c27a44e92eced07f8ca4df6a914e22aa73d65384b133ab3e7fe61b770785612ba11d83c6932126649047feb93e41372579;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd3eddb75ac03709ceb5872f3d16ccc199d142daddb5f0ccf541c7ff324eeff12fb153373fc63ff7e003b65b86dd3555d82832411ae04b41cc6c0a37a16ba5ffe4da903901e16aac8ba4ea86e79b589ec9ecfef494479b89179eccdca231ef78ae80b90e100b8884960e67c64266489bae2a721efbb814ad90790343181b42c17;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h99f2a311d8da3fc9af0f24264232b6e952dc072c39e5ec03d8e3f052121309896d5196686e62d7a2f5a7751f0c4dcf3824990733db8607dac42a6642856fa069fdffc4da41f70772cf45d69380dccdfd8e4b5e02e75f7d0432fe930c46b444016e36ff4c1285c584012bae821cd7da01da149d687d97f50e103d2d5c86182074;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7d09325b37237babc5fc13c65dc3e5a426b329f0df2d2908ae674e0cacbb9b91d8db2482e0386f03e4587d602efc2ee2ba16744583b24b3b7120a73bcad46d93d3bd08254e0480274d68f3032d5615c47b23dc4413d3f2e0d3f911f67f176978d628b502dc22cdcbaff6a49ba0c3593b610d676274699a730e37368add4bfd69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdb714d244678ad042738e26a41e76a6b18a7f36b9563608c6365836b76c0f146db95f9d575f0a320d46313576d2d056389d72a5eb8363830076c47ef158fa4b7ac70e396d40d1b172a0cc5713314282f6aabf680dabb562fcd292a9c34d5c34124ee27cae024248b33cb6cff70faf342bed6d844aeca59deb00823cb7bae7a40;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9fd2f30c6ab63d584ea3738ee258b81a4ac0eff963b1c2cb103f3305fbb8ff58fa96b4cedc98e8d1a0ba7cf4f45040efbac6f529d1e77e0cdcecf2c4cebc263bb1c6a8a080521a416116a070c08e8799d40800822ea94b3b0eb7ea568e63c690a42ade2f7c8b952997357da5d95b1d2d982a945ebdcd60f5dfea3af0bd1c1be4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ddac0f3c036558a429e5286660ed7d3aba5c135ee1dfa5d1b02ed37f74b708567658331448cb12edc0c66fd68d890d0aef2021230830d96caa2718caafc6239ac2e42b3116e5ccd91b0e030adff4eb28121a15e4beed9ce34fcec63dcfa675bcefe9d64a729257b53833c9b2ac45d4f40bd78ddab8c4d44fdbfc4d2827b8fa0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4220bec9f9af705501fb4e06b9ab7a8b86793707367f9066fce1c2dfb3dca5bad6cc688473b26153f22cbeaecca83f7b73b2bfd2dcd54fe9a701fb9664591ca27eacaea7ec8c6ffc0b5bb426ad4652ad3fd6ba4ddf95500f2dee35db4da21138d7cbe00573045720b14f7f510393155830647c431b0c5d3b242f8f8391192e91;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5077acfefe9f768d3602eeb9693b30110bafa88a278a34c1307dd3cd7c29feff9ac2fa87e319df2724f7fa76acb684630d2657bd60e8903e300db6ed3731a96f581d79ba7c4c309836a286a4d7462c618689080aad51d726bade40cd7e9a6acfe3e4eba6a29c759041a3d90f718290ceaf86e198fd1c8839ed1986dc5e85f478;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h66395a2bf7fda88bc63c9e0dba52e91bbbc14ef338ed41792644914160027393559e2b5d26b36e65d9bda9d7e567c5d2b339e180abd9537400f11c1a5e19ec0911997e3bfbc510fff19a3d424814c679f54a4aa59b6442e99d66632aa177846bd176ab508d244b3690cfd5c2c311f8f87a77a750dc8ebc31435bb7809a282dc8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4d1a10f5302f69335349e5575daa9d50ddceedb11ecd5af140acf58e38a193d9313c86e4679c1d44eb3a50b094e3fc3610585198974316888c180ea8f7421711ac0afe8ab62d36a7064f935896148548b8f70ad7ee3347f8ddc331b07696d40faf6d11e25226d190b26b789a3b0bed677cebebb4d701ed31691f8c22f4c0d909;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha15f38ba97caecd0e212fda72dc59806afb0579d03c9b13360d5c260666b5040d13832b779579ef15085f5369de0962bbb970fffbbdb783db0d5363d6457feb82d752ff749e8d46f199380f5cdd48c7428a4e7f040665aac7a93fe4c5e4c22fb584fd09dda1859f0196f07d00c5b0fba5bbd47750527d25268973f2ca4484707;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h50356e86c5596ca519624cb1e98d9f762e0ae6cdcf09b532cbcba491d56f0d1bd7c11e1d445615e050c0e1adaf03f1d91f31b1a0b9ed7f3ee643b1a7065c57dbe65714b3804f87080f31a87f8a05cb54fb9bee5ec23c43b6a266151e229cfadb95e89d7617e2f715da9bf8d76d8617d78c9bee29fa23089a03b1548087d15c99;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h516fda7f64a342bf38eda33d8a60be4ea737aad8f81d2e12e7b9d12cf00ca9673e323da9859b24b1e963cb7655b3135f984d71ba10de894bfc64a0a0d165808b1e7df121dd601e482f80caaa3cf5f2ce5c71cc33ee66fe55ceefcfdfdaf5fc21809d060eb99db1f5436f7db84776f22b516fa5242268093657a43bead95e1963;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6549daa8d5777d1e38986274703f10c59f0fa62d041b29d18bae850df8639e12d3e2db6a57c69d187fc05e8c72eecc134b569a1a4fee8f396c1ec78b7b7c95ec13a1802ba0c5c7a65287ac732143a1f3ee0f6c3fdd841ac1cf2c8f86500db920c37ee6f110fd44d66a84588cc0901e26594d5ea2a3d7c58613bf727755b04b80;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb038ea9077834edc6283270ce3f7e709f0dc549bb0964257798f756ee0d534c5e32ccd6f900bbc22440d4198cf129d582570a38b68cf3ac220ab3a779d4ebbbc00e862548162ca45dbab3d3e5c3e2f88dd86645097c565c14db975a8f5540f2a0df16f7ff5a5987b88d49e4afbe8e18f3cb75c0e167881a482db6822f047297e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6b4c3cb73426aaed516f40db56a5d666eb344bcfac9f2ff59c0d8aa993631d373d13a380a62fbebfbe26abf7a0c84457a9139dc3ad0ac94e6dbff5b8f90d2b05f4da8670b101afa457920a24693f0a881b3dce501fd5113d05de9ad7d4605f1cb51dd44f3e8fe57c6396a9cc5c416234854e082e97b65aa89b36ef229884ef06;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9ad75d0abe7b644ae68c8c885c85eb2980580ce185af3222e4e2ca42dbb0f2bfd7d70317efba79cdeb1c77a17061fc4aa5787f46bdd2ccf3f1e602406355a0f1c94b58bb230e14b508f7607c28a8e6e50fafadac2b6650e17105c6a8280901c3d7304afd1154d3647a7c5e6c368a981383cb5f65ab553dfdb28483ad4d6a23d8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h661791d0d58b24dc37bc678e8dab3f5d3019e6a0e94912c6f2b54db29b4e1c64d5e23683d9c06741f57828ee1cf994787e050d99d77b94069597547d5613ba0d9f58d86186f594d36fa4ecc228ef6e63e3cc969179a7ebfb7c6da97f222cc397be847185d7a92db5ca3b3e0dba09f56c662c7c0f43b8d02d2a78cf00a8799f97;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h22677dedc13d2e409010ffb277f68eb08470734430cf7ef2364692ea1e32b4b50ecd12cdd612b53be30c60e83cc6df48d5e47894ee1a4af55df358168d71f802162cd99180f08c2580c70e47eeb716255a7e2e0c36e4410141d0dcbc874d98920ea1c196a3b470281e2fb8f180d8c17ed14c58dfb9983ae94b8c9927442388e3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hddf261bbb94cfbd5f6b6ad65f80eeb651d2c7473d09596edae483fc3285c9275c53fce51bc7da35b3a22fee55dcbe0e0cb02eb7e42ae4aeace78e82163aab70770ad126db49cdb434fa1b3d5d6b0fdd777b8bc9577c0758862a2ecf9841fb0a5b8c89a1ff202dd11c06a7eb54d74c8e03fdb2a1f2d3fc18ec2595f3b42015619;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h731e327e6526e6abb3f0a039cdec0cf5b7b40a77a366cb31d674d07f3119d40bb58bedfd104ed14010d1b7f70f94fe1d432a466c9a4f4722870edf13b92aaeeedc6bc35d552abf3467e16e1e2e8715206c8ff65b77d2cda6b2245c9b0f38efc36538a4cab50cf07b4761d022304c6fdee821a74be3738617e8abcf63aaecc0d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h229b4f2e47d13b741fc7844f147d47644f6e52df21b1d05e1f04e87d40c861cd51b33f2b1e2e91e597262f504b21cb8808ad38fd0f9e32853c9636400b825ced792fb5d3ecd8851d22421aece91cc0dbe7ad9b2b8d329f0796a3dd10b6a4a9d9aa4ad4d1ece833cea30451783835712118b29d5613a046ce607e957ed4aa7299;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he39909180e25af76b36feb6c3998882d35326d8bedc7683c2ef8569e1bcced8ae1b942091f6dd86e9716f9fbba2eb07c4c74d6322f29b95f2cb0bd40759070a7277579abc162988884a4d7a2ebdbfc31019377bd66543a7c37e0b34152d007d2970b38d2c3962e263f1aa75bae783b199b1b836d047410bdcd5f4e257529faf3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb68ffd9b9fc294c17423e717ef991226fb64119dd80beebb89cc9cf9b7110d3c6a805cc3e2becaace019244bfefdc2601870e1ed0b3f5ed238ccee6d080e120fc21cc867fa69d61a24d70cc27e2aaee834cf79b8d00b3d64660347ac749e93586173ab89aabf1671a9738de7f7dfddb93c9dac628c179e8e15e7a7b89e097375;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h645b0982574081e0f53697e009164c37e3216a85a42c24a4df925f90edebf14551310afa102138ffd17e543bcbbb1fd1152f7aeef918fba0d2ccc49f6d192b758b7b6a256c3782c78294963cd6fc5fca26d1c2c80ec8be8083821438cb426050d1936e4842f300909d33c90de7fb17df193de32a752bdd5a73e5344802d4b54f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8629712671b0711a098304bfcd0adc0a5caefd10f239c4a677cfa569a0aefb42a9dcda0551bc0a0c3c7e6ca46399784ea8c2365b66cb840b5b7b1eba7aed983d2c71c215bde0fc27178ed91991280e83931bdf929e29cb1bb3e6ec2e7f190972fce6ac3f7213d813ab9d5fd71d4b4f0371d8cd98394ba2908a03eb9eb5805fc7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha512f35c89a52ff9294d8408eb9e17d5f1ab05de1dfa2a013647aab960af0874cda9f882d50be7984f2c8720ea4a9141b9bc8309b411c7f1712489b98cc5945cfaa052520de85470d700591d19933b81354bd7158c92fb54d717828665edf416e06fad26f0192126e17ca354a42bf1bc8abdbdda876c798b47ade2555061db35;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5722be9e5f1176ca30446027912744ef1d610c7b41f7ca17cf66ac2b0006bb2177bbb44d7c5c837e74492b3e7e6769dae5dfe3bdadb30eb814c68b92cc178891518c7fd4e2f64179b3f302c56f03af1f3e5200fcccbd1b9c4a7ee5267a27fbf540084d83ba3e02d95ec8c4e1d7a96cfc7320915e619bc57da6ac0885e96c27cb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41b4a86a27f1a3dedf36a37b338e5bfc041b2121c7cf8761d78a28e1e07e3a92b82f0af48cdbd722e6de77493a32add4809bc5b47b3c3054d75383e33a26c2b6374f1067d7908cb3a53e2f04258fcc7d7203495459be381da124acded6b2362031e39e10822e08f1e90c4412a127a6df71edfc7605313a4ab1a662225c16f1d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h57b1f595aef2fd9b60e00ace9cba3522efb90260f5847cd1a90a62c741d536c08bd5436eae0980bf9d7703687d1e17d287ddd7dcf6a8e38a5b17636b261e147bef0cc0f6c246952f4f5597416bdb7c826b4e17776d11a0a18c67fc9d4c570102f27e6b35ea36d9dbc9fe49b00a431fe388a691e5dd84b3a538d9329acdc56f21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb5e59f6d22daa9caeb34d59cf4f658acd88f0e084b106fe4180d6b0c2fa08027da82d05e3ea6ad197ec7fefe05e7fd06550fd53db825a7db8463ddd5922d1523a7a5368bcec5b468c75064e7f83353523310cbf745981a2f3309c5f166eaa12306861468af6a6e458e1a3c3c0e4ef260b302fc711f1343a5964c98aaaeff0c60;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6958fa6b77dbac4ff3055b53f757dd3503685eacf28937f5e7666041844eaf0312110b0c98f075a09b5b95f33de69ceaca1ce8292f9a4bab1f3c27def6bf92b6fc8c188d50272be1be521b04b676c1a92bfa106d875c2e8c81556863c911beff13c75e091606597f6db82b619e20bb893f276acdd2259bbd614999e4417c6b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b441b6373b78e22bfd39956cafc905699f23a0ca744435f04121559750d775e20d982018be47a35f558b5de9bcfef091a85456676eb899decd539a5c7003ac68610f4fec2e53b9acf0ac38acef9f882c89173d9c8b799e00aedf8cb8672988683a19212a430d4e07e36c17853aa0bbec5b186e1ca592fec152a2801741a9abd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcfde053a5816b652b872a4a77c147a5d09f98fa9f5cca23389318768712d601541c51de7505c6e71d8a524171992cc5a9241d7b27d73d9f7f8b9dbece6fab28ee143d2f7ecb7715899e862b09d80486bb2be784b6cb78bef74fa221acd7ae7fedf73778db61a894f7625d7abcdb22fa65cfea0118906afc86f7b0637aa87a49e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha57693bdd549a9542f5d9f01d21a05837c625fe613853d8492eb7c6fcab581f8e3e8664add26d5bf7963dc575fea579e2ea490116c153f66122f7fdc876c50b0184341ef9df47073f12c3b0e38cbcd091a455559e9772912cc59264b4e3f25b81b977a41d461a0c302793fa85313eedb91f0bda31c7ff74c98be99c2fc2d82a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78c2436bdf75ef8096a6c28a4020adc8b8e3c75f6abfacc2c9516a7f1425af3058ddbefa47455c487d1be4e322fe2f25b9a5607ccc86aa484966833ba5d8b64be25711144dde34ca914771bc7e1b788eece3908ce1b44fecfa2426e3a8264fb5860568f26f93dfec3302836302cd910071c0c6873df74784dfe14124c3204621;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h739dbfff87d20ea3dddf08fc2a7fd736aebf5044b08f3534ea43ccaa124c42e6f9424e4aab2eda2cb5bdc71da6aad65bf8b4085ab18a3f881b60be7b1ea475b324d605d514f38e3aacaa1f29aca22132480fdb7babfbf8a82c79c97daf04c9af71744c767fa7683b44abd3a026a9e6777b273e3b500eeb49ba98196d9c978f2c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdd1d237750332ea2674b0dcbefd069a402726fa1826afb2aacb15c651c6133ddfff9d032c23677d477d7e53ee5a8ff1daf37788ff3aa40e9c9385842fd5168492f64213b7dc9234d374a41c14902e738d0bafed9da07452903022def1f898691fad06364dd8ae97daadcc78437b913b01a323c663b0c6d92410ba71c1f81e46f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd13362347076c1ef52d913338415169d0fa1aacf1d99faa060460de84135c60cdb4ba4f37fc82305f0dc89dec6bb5112eef6f93fcf4d897bdc118ac196fb77b5117b6ed321f0bca0ea3409e7c7eb66f9b5b83fdfb4bb9ac37c58e9d4089a03a8830c826c94569473edf38841ee08162e1d7f7ebd7dd9a4f6ab0a41c50a6c9121;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8f94595705abf21d9e44a0f4d537d5ea5158a90c6d1ef619158847bddc60e7233c5b148f2f49c497b4ab64c1dedff7de6e1464ce015622dea4547c48b5db6f0632250a5bee4b983adda563fa9d428e057e242ddd00a5c535593f56bf52c8503f1ced520906b66aec2767e4b7dc9858e90401be1168fb453137557cc5773c8f3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c66f87cfc09263500e70ecef76addb3f700fda1bd16e5c8c7c1071ec875cfe16cf6d065bd162a511ad83d5d8ccc12a360a0774d65d47de445dbc4dd06f6c8e091662eb4fc1c538d5ba249676cfcc0b9039a7fd3676026efdceb7347dbeb805dc496ae107d85bc556e17b86137775125e869af04f5e9f275df70b3c3e1ef0b4d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5492394cc98462aad684c548b2738d4df63daee8891e2272207ca014b80929958f143b2460497389af6498a8dd6cedc0d23c7fea99a05318c0982c66b295fe491a94329e43c9fa6ef5d15949e7f47333e731f6aa4a6bfdfef8b7a7e688939c6b1c3bb824580e5b1ec13e4c7913f59c86ac95c0f0a94d56c28482b5e5634e8ead;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7943e7edbd0dc3cb1b0a91a44a7c98b264b84586a36be86fde548364303fb665356a54a1bb8e40773ccbb4c8452cb172df134d0c692a18d7aaff92ff5821f4e2a19d283495fc6b30b464c60d2d383ef3f14e1ca1456826023196c4e6a45eb14832d9ebe55dceab8b4a34284ab373575f44f4d6b8e7dd0f6172393e75df4a5f7a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h877f6edf73013d1cac6ba4a46d7df0ce5487c80f6ea599c56e98fcd0f9456ea41d0024167d1358a1905647874f8359a75432158338a911d0cca28144ab99b5a2afcef8dc0c4f59f1eb0dc616efe94ebd1528d34a755ae0312fcf97e3d0403e940217eedb96c8885e0ec9eeb31a3257bb6794069e7ce1898de60fbf601641cf0d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h92b9632f88af7d697793fb87b3b422123dc1811a5d981b1c767a6894e6273a4df4c78fd7bf48ac1d7c4016f847fe46ccf563329d0030836deb61d616aa8e8c79a56619b105df4f1405817e3c18e3ba6e9cb81efe87173cc9d438aba31a95ab91ea3de73e51b24e4efce96db470043eecd2b465a0db35d01700b1d17aa61d10d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1566bcb6e67d3d717a806584e4db3d8ec937823649eba36232b79adcf7b3051e4d9336ac5cfabbd22bd0e78d084494cf3c09d15bf37b65ed0feb9dd3c02fd4c2059221ccc9d4b09eb551aaefb70adca00de3a917ad22754f029011607a02ed45f5617ba4664c127cf5815a859269c5457d650afa9103a0b4f521288f5e2c5e53;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcac38d24c03868d4ab612f294f3db4b76bd18b8c6a9e92cb01bd0357a99a17cae14ab90d7d40deeb557757711f88903bf69818d5840782b5694d182f15d292dbf60f86c5b424bbaab1ce957b0ac9411466e81bbc2a7ed81bc7e43de0e2b7dafd6e4c294be52487c239ff768cb3448a93342082962a15406e0a2dd9ceab383d56;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h494ab6aa8b9b337c2c880e47645806d56947da75af03063be24f7935fe77faecd18ab176a7dc9ca4f4ed8bd1be698633f265dae9698fbf0a3bdf0cbeb20811881eef857eb35807d8ab665dcd37dd6524f2473b3e3e92de91a188f2486b7c9c1cf0518787aeb8ad49210855ae9261a48bb95b187130b143c41e1d30de40871046;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2358b2380ebd4f17c1c3390c690b61b1fa52f5d9c27617eceb60482d85359db2b130ebf9056f53b333ff83f7a1c8664b1766a8d8f0974a5afb129db96434cc3dca47aa5bcae2e5fc581ee6704772fed4de57fcab80c339428bba147c06fd265179efd7825069ad0e88b256e6df06c2c20eaa007f7bffae26371ba0ac7d03397;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb33d002e1059cdfbfb3bfc09f14b592a2209b0ef806c4e6e6d6b1dafb1178fa7fc2b280a74c0b23a7fb412cde449c1896e6dcf78030e7a1bb1f103171df34ec5c8a620d797273efae4a40003ae9ccfa3a8a300cde91a9d5494f9839a4990b0a767b7b25f65441fb85fbc2984658fb4a339dd99c94aa6aeb5b337834aecf2cb3d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6b1294aa6d87920b7222cfd1ec39195123f0e5a1e0233565c4cdd01e87d02acf47af0303cb5d60c526405425fd1985a7588cea9b2d56488077ba8830c423d5ad1efac22f5c8ba092e296e14ce089c13944d6371d16edbaa9ddfccf1948756fda1ae419cfe4bcefb90cb6c035392356920d2240215924601adecdbb43c6fd1e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hae84bb893e96a68d3149b026dbc81aadf48b1462fcf25e94e74834e02d225cdf2e7c42c695516e8bcc5e36ba6a177ea2223a49f03f29a694d673a4c148785d1b136494273070a7fb8e3e396fabc44fe10010ce7b69ade263b8f47bdb87273923d5a09583b6c885e8684d3b4c5fb0dcadb2ada96d113d30641a1b286117eabb3c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda93a2ff14db36819b66384f0b76de36b50bb03dc1dd2fded85fe6e33fd1d393d27f8aa6f9db6850fbdaab72947d96011e6060a521a8b52a3b9877f276744c13074658566236665bf02cdf40cc3466086ba369b62c05d39c50a11d88c12583d313f002e086351c7ab67f3af3bad720d01eb72b76b0aa9df6d252d31503c45030;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h53dc24b91bf4fd896edb8c7c6070dbe8b9d5d11324ca73cca49436a820e151eb92bdf1cf001ffb25703e79519c483a0a8fc80e2ff6c721fef8e9865cdde2ff8fe2923dcd6662bd1c581fadf4374e813d43eca8d64572dc9fe66963e3539670dfe92f14c10ff1f6c25b5f6e0e8b751fd24a390ca8b9df2fc67fdedf01fdb916d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h302af6518061d3be66efc9dc4e55617c76d55f9d70d0d2c53ac6ca1f2fa68b31fc2df79bc00f341901d0cd6d90a16c88101f58af47e4e5176eb485cbda808ad53bd6110f349797db10f93741da13050cc29e051239dea637ee6cda388a0b7e5450c3233514a254e1f36ef3eebd2c8e10feb19cc2a8b4496e1ba4a2498161770e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1279637c2df8bec59d720167c6c03c3cc514d5fdb105a4193b5dda02cc0687528da33b09424ea7db990ead16d7ac83ce4ee04c4bded1f7a4e1624a25ad3d4fb0816a4c1876d0364f6eab7eb7260158c634a7bbf9a98a0845f28e0aacb3ec92152244f5510290f7ab8c5800a482ff83bf7544e236379f90f8ade165c71bc0ab5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b1fc7b4a6b1ab16b91e14ac638ca09e4b8f4791917a1d0be86bf2cd6da056ccdf9b0f9afe1e98eb0b02733e76b98b3cfbd9448b9dead3dea2849315090113031a9d9b1182c81556eb777bf478783fa9fe504b3cdbaa9b2dd3b53c733f88504c5524715e7b6cef7beefe596ea1d95ff051443451e209e938cbebce183071045e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73ecb02a7f8bdd4e553c10a6d3fe93154793e164c814bfec532bd64b0ab673113811e2cf5264a630e6cc3f125f92c05fa1b885bc10b47cf8ef05cbf59266ddfc63052cea1ff3c3c4c30f595b8d58885bf363cd518149f34da8c8c6ad646fc860a8af59beb0275c9e5d6c38e978b935e0f98b122cbd1cf0ce3fb171d462db0685;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda5880b06d9abc7ec4c882da82925cd7635eba8a31bfc698709e512329ab51735b34e4876ce4699256d28a21f2aa59ee3cc68b4dcf79b23fd52300dcf91f390ffee00b063cbdae159abed4d9da1d920655affda6fc3fa17add29b3a2769ea09f44129cb2aa8194489067323d29e410e61c30bf5ca3373ab3d8065ec7d4f24940;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbaee94c5ccf5cf680c907beddbd46a3d0c2a8ca01defa52c61abdb8faca96be37fc6fddc982a5b75c5627f6714341ddd19b9a7abdd109b0fbc928b807477c4b18e48c2df493392de57423cf5e8915e358b525f1e999ae93f572b27fd891150ac79a94b183f16dc834691fe5d014b1f21aafe428fc96207fb4a4a5d63908e4349;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb24491d855ac7ac554652c6889f4fa92854d0e6c3eb04e8f55cc2180dd4cc43ad2e21c67f9f888e1ecef1e89e5e1727967ab538d973b248c87908517eeac418eca00e8a999f7092ca9d0cff97472e4495079cd764e1c482d42fcdc8344eee28455ed0af412c152c67c0f6bf47369b1b7f95ba4eddcad79b284c3cfcea8ef3ac8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41c7c0fef3fa8233d0ebb0c851b6948a7d4a92df4d2b1959be7e2e9679aa4041bf0b365eb34f7e6988ac277961363e9a8ce37e886bd2aeda72a0c6b660dc113470802c74d75115344069ad0b7cb86e30d98bbd722becb09a93ae52f3474d3277329a94a4bb44528ea10d7c088e7f4ef24f1b2b7d2fb3a90d5079b858867388a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4fb209356cc2e45031a1d0f4a50f9822b4aae2578d5cd0db394669e971021bd6767259bbb609dcc234a01a9821b4d6797733a4418c25127097880d822b0b3972d931ef588602e0da7764f7ed3fbab6052c27930cacecc7d882e4816dee215c7fd43790677a0ab63b62c2e06de0a73cb6135c758c225499c708671f1cd5283784;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74aebf6782e524b895791abc207bc169039f0a7c8dedbce4ab76447346be31f6ba7ff01dc7da53f306bfb4abeb9b937dc2e8a3d9cace45f40068ac3075a6d98d26dfc33fd23822bfdf5d93957ae344fa3cbfc74046acdac413d16d7e774320165091649e9d7d156fb913be4a7249ef4e5f7b2886428d1b7c34bb9ab71be4c47;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf67a2213cc63ce5eed9dbf35b366424f5e90636560f3984d75a3c650d44b86ff56dfc0b143c350ec1b5a48d51ac0069bf8cf7414109896aa9dbf064a32eef013ce21d172dafe22b44cdf1089d4f73c76a54d7f35ba7fe7dbcb16bfc1e6ae1c301f7e32e390b6a0e50a8f13240f4d754c799c13fbe29be711391acf2b017d337d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2eb85382af28e1d99857f9bac2f6ae6fb32d01fb693f4d752197e1e8f90587d05956cf53fb05c341382ecb5388b79e96c33f4c67a65695bcb41c988336767c1ce4d72665434f42c3acc5bf187eeb48b7331975b43eaa4309bee302e158b4672a7671d6a0ae95a2657c5972e5f9418bb8deadeaa6d07f72b9e45bbd805bec61d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb0f472c9f3c529a684db211d6b8b05e6383f9ca8b7298e18425dced198998db4aa9caa232cbccac1d57bd55768c3c48cddce1d03eceaeddd0475da16ed233a826969658319284e075e17388137dbd44eb7c57a39e783225508406fcd3eb89f3f213dee92cc2505279f952272dd9680bc497876d6eaaafb7e9b5adc8d0058891c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h932b112a1e892d85cdb4f973a2b2f7400e046091b878b220cc249a8a6a6b605ce4318a7e07aba6dda976edef3fb5b8c6c692daaee2ff3d4a7a67dbd80c94558f02e4dd051375ac41e80a8ddb2aba20a131eac9f857a6677912f73894ecba052eefcae044db73fa7c5e271bf518c03e245a6a182a3d0555821d8cd1cefbe9e9a5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h182e8d001c335a33cbd97f69da7b11d9fa52ac129eba33d8987a89a0640f974d0fd0a59bf7d8c562b46a9841cb62b0e1c3dd21e54fb1164c8580227c352ccf0b1e23730f30826203fcfca37fdf73bdc70411481e44c0d69ee20a5c252ea453a65e9340d41731420957b0379279277ce276c07548a6cd6163eeb24d4be647f11e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h92f15bdcbbdbd176b2a8f337284fab3dfba8a6bdd70adf08e8e19f9e25e16517bb8a3e4dcc649e9a01e86989321876a7ad3597eed75e911751b450e4150466c8c096f07565b3c619f10437e760e937363a24dbacaec4a3a7d47d521aa2f1f3f7769e7bae08d7390b860583b88ad0c0facca82d4d91ec47c769aa5cb69ed059a4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h540bda8a30290155ded0940e90f3f2a468ec8a2e653737405e344146338b1a0f893f76228d0cd5be52ee484ed35dfcf88b727b475057ba3107ab1f274cc867e23c9fc7e7b967b1d0122582b1d37696c365ff81e8763c9a7bbafe4fd81981d06e17221cbbf85daa6bd406c23b1a7edd76fbec9ba8cf3349f43f9ffd15b70e0ba2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb0e0eb9212e58dad4fbe33a418aacec8d4befe9b80f96322313cb8bd1224e8e38c9d9ef481b0d0f1c0362701396b3030fa92c09d0f02b82be88350ed9d469d0039009ef0a54b4a17bbc783f6800bb2dd7e266ae8785841b59259104d8ba8ebf049cdc04534a3d96affdd3ac2919328569e1386cdb34b5334ee716717fac37a2b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0bd9ea312fd85c09f8135e6f11ebc95ed428bf5124f9e4a4b2837671526a424a4f483996900fc722194d3811afa2dd9227a02eeafa8836b36f6cbbed31a7436b3e9a2e70441340a8df2e784d46db5fb839e93e23008e8f214bf33788e2e84bdb6779980e0ede23f1d5623428da9f4c86915e96e44fbb828331623e6b269a636;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b6150ed71136793e80ee901e41fb454e34c3b13caddae695cabd31126ac67d94aab910fe18d3e8393db663a535395662a1dcc348d9d02e8e34bb333590cddeeda3f3784bc1df036d23c1a18c36e8450ff5604949485748a48a5343c121feac443b96ac91510a6475e2fa1e1619b30b90e149fdb4e1968950af6f499d6ecb528;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb7096f92f3f924a5695b202cdefc1727a904a1f1a057eab84da5256d08514b92493ab10cb789c45c5148204085d36c47205dc497080cd04d56e46e9d9b40b4902ca0fb8847c3c75171dd83b5d4dcb9a3333df0955dca3dae62e92b85045b38a8c58d10a09fbf0a1d8f71166e60f803c988543a903d2a6ba6d60efaf2350b88e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h147ce6cd40407a996adb96c793ec2ba9817d3a8dcc9bd838c84da8174651f6cd5c51ec74b9c0e6e46ae018d510c365b05f2212ec268568b1649b2cff7b5f3168d040834a8d284169fc2e50021131aa7c8ffbf792dd621c814aa9a3f3b00e67186ad9361b00e43efc97430f245a9db0e575c52237f21267ef6f0d558d6f564783;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4de236434588605360b5e4d99d127c9d6f65410ad40ff5b52679bd8fe62417fb6045a7655204694588e7675bef3dd763eaacbd0c7e8867504537fc05bbf0024fcc4faf37dfae3c77af7e03570906ef78f9046bf498e56b624fa035448a996880d5d3b30114381a2647c71003a7aa02d6ed7027df4bbd7c0b9404eb2f14117052;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62237b1b3cafcbf7b908b76be35977179ef2845d93aecba209c56f9147802e831182875d93fae5783d54d0922e4f4247df461c0b70c99b0f60530d325387684caed1dbed9714aa61373d6a19a0987180a0f768a3935613ad7b1be44238538900591900d8b6da4f60a68e2e2a28b014275d5b709cb9c484c9bb99b1e4f22910bf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7c52fbb5cad7bd6c9ae8bba0095757ef2bb4947b5ee89f322618724a72e1fa51112fa7cec04ba33a962dd14561005a85d4e3128203e8aa3343f364448e63916c1711c90a841f2adc67fd85ba7fd6d2324422f27bbf1dc5a36549dfb4f52ab875d00e95b852ac3970c975307851bd2b1bd30db9ddf1b012d53726f19f19f3e9a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1464bf3fd23148ed49b266dc22b825e4914fe026df16b5a4ce8de196f5615bd599d5d6b2fe605c4aea3d773e4f4d460d37e2edfba24c81f6304ea40d2719a50348dbd277316ceee11824e189c5e95641875ef25ce5b6ad73ffab15efaf53c41e736f42441de10f73ba6abd00ecb0c0f3861ef511b0781600184fc816fe9d155e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c23a75a3d1ae5ea0ba21c8b5dc99a4911ffcd5f753e30645298b08a07131ef1711b0c33c6585e649a32d30afeee6e5dd6606ce94b05954c5cf7d420cfe48daf72442b9ec5760f2fa93b5fb4b384c1e004756896b41a9077dd774ab6e2214f7a41a79fa45142c6d72aec599c45192af021784fc49e058089d6ce9dd2534a5179;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h379cd2ba9c9cafe9bcfc432cc43796478b4abb5c2cee94a94b9a966a1d60bd4f15f81ddd0eee1175470ba5dba14a8c0a3193b463ee9fdcab9ca2e35e804228a26c09557492b6781395d65551fcae1a6c51b4ecc1d37863e7cf411508ee34fe97547afaa28565384c8aeafba710e356ec3d4f81315bb6f6471c606027b7b6ebae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37bd74743a7ef310827eea5ebdb32867db69ed2d7f97ad8bfd20eb37143db316c60558eacc5b39c9b653bbcf7cce1e2de592c30f175aef43fb436abc7aa06b8a5f34a03f20d1013d4a906ce3c0450492d516dd6a78d59f632177e225b31329a0f5b3f62d40f3a92788d1018d0ff285bededbb2aa8b46d4bd50a88a3153762b3a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h64f7fd2609b171c03e7d4921296ac23d9875fe71df9fb8ea4a35242df24a0d7cc08bf203f8ee998608003a7c3d4af76ea0f04a53f997c3c7bf9bc37afc7f23bcf9cd7147f87e262ba5e38adecdf5c7e858f783b1656a6e96c45f1f614a28b13b1cd45c585b9bafb17396151b9efc8709d9a400bfffd8223ce7bac40ecb84034;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9b985e21579ce28bd29138de8cb4eb527f15e2bcbf46c8c855bf2a34a9765b2d007d7c5ffe34e22c25444a1be1ce143d13a6d9e3415df2f92d8b78dc71ef92608d0d6089cef428eb1748d5eb9d019b13cc9e2321df69f7e37f2406c7913c1b4025fa1c43774eab50796046c27ed3f78aad68af2aa5771e8f83fddeb76a39524;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ebb73b0b74608146d2bcb863714c963ad37f101810e2b49a725df4d9e2f137ab9d54e5f447909c4a7ef43fa58248b16f623e60f0bc6491bec9eae3adc682d140e400b6de7b74cabb9481204818610b5af3b7214f6319315e7af8766094e2a41c65e59e03b11012611f036c464e71e30b1706ff870aa86c06b75d2511c2ec2b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f833d6c9a588605233f823da7b0d6091da28c204cd61e283951feeb1c0058260ae9b7c5a784d2f5a8fc4aecd9bec6001feb724fc0bad716047924bad6cbae925ccd9d3130c8d136458ea5f03528b6df19d82ee9c21ee3d6be3a2a965bf034e6c711ed5313ee35729c4b11b704b9dcd630a31e184a318df2f6de1aac2bedc335;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9e807d3c14d67966a27a3d20a06955dd09c2d44e9b22266c9a9eb2c7689d64001a20f2ed8df7d3a4a225e3b4438fc8870c269d5115fa25bb705202d82fb71249020f07949eecc9322711a4fd121ef9ed0b52c07bb494fba7b9477e82756b7c1da58c77fe6af3c8a8c4d498f3578b2e692e61f6bae674cae7355c02c5a755f2e0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf6d1bfd11f6edc5c4ad98b785955411637ff98763db4e22e1b3a4246d2da3d11816fecc48b71da31c1315b58bb0ae55a03a275a7f360a664773c83a2507933c4cdea7f47438c9038f272c593e4344a6b7153e1e8d59272e20a046beaa0f59d47c9d44c1ac5c89b78c29b37a4310a3a6d3efe2cfd94ca82b699d947050eead3f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c367e7b010ece6b8a4a5fd729a43866d463f0785e448e51d6b8c21f94d0969480dd8b618d642112104e56bec1057975ba2a2ce706173549296fee6659682fc0bea141c8d2f1f3076bb1270175ce8990e2f6b282dd0dde96dd1b03f30fd67a8e94f0a1d9c1027b7fb34355af548b294de966f603e19903de51365179c268bc7f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4a9ee1be9ba69c37503702b4e78c04f2de04051251dbca1e2982d8167233bac2b90de36c63fcb5f9ecc8c9b38f684807a172bdf3a0a6862d8d92831699b3de10af5b083a56aacc127afa4b19ef8e265d354328dc6a7ddc3b0419220fba052f71dddf21a90fd3f2bcd811321d4a637b697b19f940a23bc7f2a57027f99e86f15;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h996e87649af05a0841332a4808d29cb54c62f173af905349a7e64fc5141ff769f8c2c7feee318f08a1d50bd47562449d73cc821d2c16368256656b4444914d9b5daa08708b1267534a33533113590f8a81a0c597bbc2f6e9da2a20ccb297e724a343dda8a454d87902bc16c3429994f23ec5a6350b43be05d508880246a5b852;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7a95432025d672ea470803d9ff530d274c183786af986c03538d9ac34c5bfcf2f76f35c3fce14079a818f823790f3fc95adefd133793eb969a561bab53359627fec7621e93ba6695cad212cee8f754931abd4f97927a763539adb506edf65e295e1e3b4944a3e340b092f0ea46a7d1fd59cf0d57a11d684551dc0bc9d2005458;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc6ef0a9c6eb41255c64aa0220cebf57302adb86458135ae33bf51a9c6e0738801ca92742e45e1ec6ccd98819372ae490d1d4a952fe65dc1e8e7984368819b39e19ae199f233392d4e05a729003ef00ff0bc8dde3395974d7d83233dfbc6bab389e55d4b026d0f038d661970a2498472443ee7cab4ca1d935ff8b9aa3888e9282;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1756bfeb35835144c37b6a91a202eaf2490f8cde530400e91ee0fca849e3c5d91bae8de5809b1ccec98d70d4797a17f71b0d8007f7d4c338cd64f28d1dd58047fc657ee694ccaf8a761011a5ea1e1abb0ca7d403ea32527d34fa54597a437ad73df2c761a5c196b8845ad3e574ba66d0a38355717e84eb083f57043454230360;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha24f3123aae152b3da0b23b738faf46e00140d7ce50fc4370e7ac063048e6c59108e26a580f3ee169e8c6149d1db754208cb5c837f5346935e48c5d3b1c3e10bba1b92bb37ff0fe438608b171856df3a65a6c3f2b64d4786373012f8485dd488412be43a5bf6064564b349e6fab435e8bf0be4783f9473447ca74e1eecc32d98;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b1c12e27c5b00607a72b2951c4688b91433f5b79cb3814555affe58af39c595f588d315a383021c772ee8f136e07797788a467d620822401a706f8b2d7a06e56fce07e9bc42b9b66f0e919dbf36a2893ec3eb6c0387930c63420cc1d48799913d546ad6f3cebb4c20227a139fe6c4b475d19c84f4bc0ea5d068f0d0bcf2ab64;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c3f228c3266520a6543fa23a7f0286cd06c90bdb365c24fc5c2c3f8d98b24718c807187ef3b1f0a3855676614c641c31dc3c74d926c5519ae74f6f09dce3141eb8e2bf9b75760204a4fde9d41b7be6296ed2441a2b30504d346015e7580b394d25cd43bfde126fe9389e010296659c404a94ed36b8a34b02a29507bed8f25bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9a70e0f715f7c2e55fbe59664cb281b75daac4e9dd911a333e3d344749593633098a8015e4002425d15e3ab9069bc757992ddec4fbbc623351d7833f021edbb3b23eb50a21ff5731d66cba6da54295a7d3a9da1e4afcba37d7d95e803f2f7c65d29e1155c6a8b77a0910bcea7ee205bf131edb90e4207139e24f55a343b9b35d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h138ae060b7970fccfbcf9cdbb320fedc720f5ecf8ae7529e34db3f5725e810690ce7c269f9bc2c262a42268d856dbbe9cec65b309530fc92e8955d5100710879d38a2c0872ec57617dc1a8d2d495557ae688a64a6d4ec5475b55d2fa69555a5a701e8dba9a85d95a86b234be62c22f83a6cc32109947cc1c47d720071d719b3c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h573c69072741c827f9e89c5f154ebc3a9e4f1d1637c4e7b3714ea63ab5fb83aa8c884819415645d3cb6fa16306f9bfd32078abd58bc156a84a9d8e8de53d76f064d6fca6622d294c5999f2df64b449e516c00fe320f56ff238e7d45ac923d454f584d925cd98c6152b20993b7ac6914890043b10c422f01b00f7cd99ca91794a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbb6a0b860102f4627773236be349c33156f0506dbd195f160cbe70512d85bce5b1ab1bfe17239bf98843b3834d431a03f84db6336abca10cc31134219093d5cfc3005ce285decf9b890903f9c97f90cd5c77996f65344485af52ccca6b1439c79b604fc8e1dbca15b77a441fe9b154c7d83ed3406d9bd205c1f019caaf0f473c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7c30850ca6f01d6f3afaa0a4af3aa00b8c04dfc31ba5c76c6d1ef7177a5312d2ebbeb5959baedbed484533550141f726a7ce4e7e152a894f9a5e0274ab9a2b587d19f25ac97ed6162a31292efe04af49f8f89933e14a58afb8acaf526998c0f6ff314b2dca6508f33d533e404823fedf3ec91241fbb7768acd0aec4f8071a38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6096e73184d3c2d1203585171b59475c26d86ea4610a264769083744c047d9605a012abb2c2d93a7e8407e826c9381056b93c3e38eaace06ce11476309320ea0c0043e11f55692ee69d4bc9213eac0cb0e0e134f3ab1901d06e19ad2c9087f291bd4c56ae88d2c775448f385921f99bcbe934cfe4390c1e80fceb22811d05366;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h800c2a3a31c61a3ce6122f1ebfabccfa38142fea344ed6da6576b8a0027665c18a598a43c339c7e0d5bd9db00e4cdbe79e824de08e485a21f580aaab1aaa6549e03e3d32ceac9b9d5bf0f2fd8e09f38864a960548119e60e6461837abdc260439fe2465609088434086c44c2e14d1ac26b68b6dbeea66be93dd43ac5c481543e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2fd7c77405416f239b7916bb1130e4d7657658ca0f8904066865f17712a5f2c07b9e6d9792a02eb594bf7411ad0565223cb5bc3856c86e3f0e329ced47fbd2316c521b619dbed97db4981b223b9d378e925a5f410159569a9d3d2e6851179423734d39bfc72dcb011d33c78c4e6d854efd0ea8f2851c20cba47fa8da93af7c38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4b6464d55581ffc730e4f80c763d49fc4d775538de7eeb6b863cf99426d628d8bd054fc175a073511a5315bcc679aaada91aa4baca12843f9eeda05e835d5be8b4ade0d66cd12365c870a7558c42358c1199742a12cf9daa67c4e0246bdb8922e0d5c9fa255414fcc45853285101ad166531756938243a7e2ad731a10b7298c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hefc48b398f3ad19763c86cdbb568c49b6044e4807f01ec5e137176eea147b9453ff839b01a2d2009b5cd8877c8d5044387a09b6e2f667230d0af721a90e1f3bee677afdc2ab11f0eb7ac3ba67b6607d36adb17b20fef15f29afa82d88ba4a89cda42e96182bdd525a73403c751a4385d111b4e103afff02325301a98da7d2a09;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b3bc18555d10c20aff585393bab94eda0d9d12624ec2ec42c7e09e98ef3aa0f8c62187377266cde6e5a190f99ab6f7792bfb255d42bd0822d0694c35dea61ca696e0a56383d7da8ad3eed4ecd6bbfa13de0fc53929d7f789dd13237a8cac345dbc0f1e3e8ef29f49f35b9399bfb955e036cc38fec62e58e5e159ae91b24e4fe;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h746b356603857744c9ca610239d3fc0cbd2b4778d2baec3f2c12fb4a10451bcb0112b0bf3a91fd566c5a63ce059fb09ca67b156dd2249e1496ce269c25cb615fb81bab064cdf3dbd2506693dd86e93b52f6bfd88fc3d56591c709faed563c2dacdf553175866573e4341590570604f7d3748fd8647e8a376ff0741662e4230e3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2c44ac600d003300a49b783ae41e27c057a6ae6906ffd86fb585d43104a48c200123870a4663e584ee1010f2f1c1d5e4fdc929afc19e60ce733ea4fbdb5a1e5988ec55e39b3007649421a186315d0901b174f6110daded739178d594964eca5ecbd1c38de404d1dc232f22e3a073c813ef65bd7ee5a1f4e81a2b27308b35b73e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h557f68893c31bd121f372cb99eab16c47292e44906b8ea0924bb3f457049ca416afd2b040d94abbf1a3a59537d9bc7cca6e5fb297bc443c1d9f8b1755e78e0eb5ab556a0025772ca1a904fc2cacf39739b71f275a48a228fe877b0b512508eb1dd62310917c47efdb3491f59c8e0126163f6d33cfe558abbf1ace882c0ee53c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6151383bb83e45f423973261be62f63dfad44e874f07f08790204d14912bcdaf81cfe9f3e4a8470983db26b0c4eec56c3e3290969c9895324feacdcbb17225e82bba9fa7f27e5f4a2a43f86934340a99b560dc47409dff4378e166953caffb4aa0c9793a92f9f1ebf4b418da285230ab727bdeabbaeaca4338199b69f43e75a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc7c25ddc7dddb9683dd10cbca81956d91a274e3bc7677c62ad782d065edac93496093c42bfe1c86a10d57f2f7ebecf1766752c02c36e219108542faa06320d487feb8464aa4065efd04f2f94457806a7d47f9486c85d08a25d1d0c33be0c648dd0550276b964d6106e6a7f654a80a3180ef103839b475026abc9a318408a4270;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3d757c8e15e6acc77c585c662c92f7bb150aa192bb3b64755f629a0095a498ba2287e54d5bd35fb2ad9ed41e200eef07cb47647ae32521c01a8c15c08e631990726f6dcd69ec3993362c7ef9893e580146f1c65e229f7c3ae0976d76d602055b554ddfa1942061f3ec3e26eaca6ad1db10cceac63a8734a14a327cd4d04e95c9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h63b163f06714244b55e741851d1a82db5c9a4cf92c7f98789d4791fdf932648aadf135b4f0276868ca1e3e5245d7915231a82ba7197ab485204dd84c4e137fca71ae818f1f0799e94f7f771893a9430e78c8e0d4e33b9f991618f99ce8465f71fbcd5d6e3717ce29297dd13534c6408e41d2aff2ca22f2f90be6d4df296abd26;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h46c735115970a06474375245a46795108fb9b58cabd5f28f9ea6659bf112ac12be2ee9651f180355c4ce97fc66e297c782bf9f327fe77c96c3c25e230482bcc79c57dd78c1f2c47fed64c2c42041c7c2d3dc0200403c9b527039cfc3ece0239f4cd4c03a4afd284245a4c692c40f7db7bd2017c9353119fd2372f264a3e5d576;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc0d6bc8b488637288740aa4cb33f3cb880606c2e7ad9a899ad437dc069811ac0836fe7ced0b98d047bd31ba3202424a549948e371f9985b025060abbe6322465693ec45511fb68504470cc696cb62b2cd84721fb6993057d7cf1e36b3286c2cf34fbc2e9218356e3aeae683455e2e1cf55f24050acfa02c350216a61d6f5e7c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h55cd3fd487db9ef9263d0ef50c38cb48dbbe4ab399fba2054e429123efec0d7b0c8c5c9415aeb8c60197496779d2f22f9db6628e32bbd17435835dbd3df47811768f23c6e622d6e7fb94125779617486bc0e97c2bab9c0949b8ab9ea1c5743fb07c77f923f974fc3553147a3d2ccafa3d8038dcf5d9bfb86578428b61e65242c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf774a8758f666fb3b604210012448609b21d6a338979024d5765f26f2110cff608d08371ca13211aa10a4b9f3f80d9e27ec95a5a67d993081efc73d9682d7d8b68c42d362cb5dabb5016deb6b9cfbb78af23fcdc7459acf049845dfb57816f2846f942a845cec614a8590bad6645928543383fa517cde9df8b21d8898be6f7b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h998c6bfb635913720834176b08fa585a1e69dc4de557a64802ab101d735e34c0ec2cb88acbbd66ea60c87891f42cd06068ce4d710d0f01d12bf9cc209336034af39f636e6ce3b880015b60f44130edd22a5c836b9e68ebd7c0a116ab96c30f251221f0cc21ccc1f770a4d6c929f77683fd27d66984441524979204baf49fe2b3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb0bc08758075c342817dc4291bc2ad7fc55a991ddca27896e5aa35024332b18f842080a1cbe945de2bbadbc32ab5141dbd58e5419c6160c03bb54e0f8141bb66fbbf329df1dd8f4c6e96d58ed6819c247bc918a066348ec9826b73b8f4ec0892a2a2ce6d11ef014f6694510919d71511edebfb0a436b6400e94f11d28b79042;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf458ebcdfa6fb042d8c9348945272f77f01cecbe6d8591c3166c6026f0ae14cdebe121fb65e4c779bd1ae9349980131748229f3c076a6c76a4e4b7870b466e24ded3e08fe94a75a3c8574d1534a84aa8e43da6b6919b78920ef52405178bc661e4e170627d5eb6cd759c9984201a1e22b9fac1be9d65a62974d5f84f6bf48d9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha6202a0a7099571a1505167b18bc0aac44d2bcc5025e9c0a24f144866feaa73a0fbb886f59eab742a100107eed8228fffdc9147fe66eb3d0c479cf009da5c0efde43bde3fd3d24154cdd5afc8ec2fe90f05419c4d79c127b4a79de6650d4329d1a15454ef459080d0c66c2c96528a314cf220f45dfcda7713b6b3f084de321dc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd12ec5233ff194258be255924b32e6d27138abafdd0efc01d6900498904b3e51eddc7eca0f2ded8c5c793d1ed06aa8298f528113e7012461fe80ff2e5002cee3667ea295c092902607141d324f2490b67e9346ba10a6f3d55aae0719141f6ccdec441614fbe34d4320ae8573916a9e89217588e3248c189bf1a6362aab76a72b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd042cbaacfa6386f7d5dd84d3c20179618492d099797a2ea7308cf83d847b4964f7762d28098ebd031f3828b59de38628de5424fc290d8009f555110436e7fdd13b751a2fe7f2bc5bef8162ce8234326ef22233d5ff757234a19592e740202193703fed41be0591301a9f8572a782244d66bb811a3d725e57e50787672577ec3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd99850659ad086af0f4bd79b446aa357713b928aa252ff8d01435c00cca9c91e9fa42b720a3991656048b6e22bcab6530d690de76f28c17cd8a9bd588caba57fc58b32ef1e06e3956eba9be3f030e4f2d8502878b47cf033f484f428f524c4baa48be01689ebe32de065679250961562f59212dd2399a84de003464d5d80df08;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h466d21ab29179c9b47e7f1bbe5b2c9600b1c7000a9da26746b8935ff2b59c9151dc94cd5ba847e9cd4d136f50ecb458ee52df369a1bd08819369294537a6aa9b04065296647fd71e182abd5647b1830226b0155776628a23c10fe6cf4064281a3e29950589be4cb84aa5074686e750faef7835fa20c1f1824549225f1afe5bd8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb8699383a142437d4b6af666cb79fe58f2f10e0a347adc0ef92e9344c050ee211eaa85dabbffa9f0faeeff30ff17cc1d7453e2c07cfbd40690bf07789554e1840238d3fb779c23e4a657fe7cc0eb87e94a3e08d7782814abb04dc526610022c5cf981383087c4a8db278e8d9623e714f2efc5c2577c85a289a5c8b93ec29344f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5694cb1e67452ae96b5b031b14076b08d5aeb91d2d75d6c6db6f5e438c4f0247b21e100ac6bdf35a74bec13bfe87103b562b0b5dede7d3c3c35cf5bba1070911112d58a08c28475412d9f4dcae403ff4a13b2072c5bdb2ee28b25f49b5b5da292902072b2a764c2d49549be4fa5b30c4740b3ee3ee7a1db0bd5a134887866198;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ccc20364cbf0f4265458eb66a4c9f83fe736e33f1559abc9c07bed31e8bbee6866f2a3396d6601943bc2d61fbc73eba5ca4d219b75087f779ae417dae5768b4cf86f2e6b6a289d000834010d0a64ea70464424b24e02a98f58db0c0dae33ef8d6f6f4d02feaf481460fcbfca5730886b2fdd8f5446f0364f9c3e9f3ac20d792;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3c57d1ca071929ef9e7d4e5dc4ad7e062ab21ca0027706e4d682a97c7c8733a9b82a1521b2c6b35ca4f3cd839e7e41947be5887bc1c6db9f7304ae4e8c6e408651b7df5bb8848c2fd81fba07b3ae1d94e0e36e02a2dc7a2231928c4c8408f5d9e3b294c1d6680b0907c3308b57ba040ad6fee3ba48610ba0e6c57baec8d929d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb619de91d2dfad79fd5a26dfd0c1e4fdd93be8578c14fc7d46f995da71bb5d466fe5adb2a655a966d1bf80737d585c4652def92c7c15b0be45744cca40181cf42f6a0778a83c5edd5a9d321f95aa4c39abc500e529fab7e4cb7e4566a4c17324062cddf86ccb5217371092c6a273e8fedf8c9ee9d412e6a033d06eed0914bd7a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39d984bbf49d771d2eaefc157e8797432d70bed81e9f9ae4ed55d222a03050b1f175a566931c3753b418d964107fd65658b32300e33fa9250a5098cbebd4c0cc9118a0907d99d0c3e887342e4bc9645a9c92586490259e454b3d86fd7ee67e638f4a757c7f47b801a9e4bd625e0cfb9c25dcfd4258b5ad377fd0bc85c4600b36;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9c8a84c849c2f0122fd3195c2c7d5ac24f6b796917890b0d0395dc3530a4b1e8d641b35e6bd58c60c7ee4677c4b7ab5038d66271ef7b30fe54e60dfbb9a34dfd2c4334483fbd47f9ef1704263c03695a9d6d5700636f70e14bcd16bc489b20d2c0a2abf5ecd11b32ed1f611717efc9ebcc78cf50af0e933eb4e3b061b03fbfbb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha21658c54726992346a94226537aa66affaccd37799d915e7503ae5065769f285a7500bcb222b882636b05fa82e559aa38424f64f2e54e94adc92db5d4cbfd6fa67116741450d110aa56fb0ce377679a46cf4504d7f7b732e5c473bd5b8285feb3bf6eb9f6c511737a56014eed6723c3d462d4432989d26aef8c87844fafd7c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h86b786fb9abf842f056de436cf55413aaf77ec9630c7594a018409468ec2ea502d4612df39a8b9249a547b7219a2eb5d7745b6f8abb7b55db2e14d709ed8f1dacc88067afe2a2b8b01155d47220fffdb340402565fd44239c775d2dc2a1900bbbd8cd49f5c26c79ea0d304e1a817d861ce701d4b451330c3c39607ce0d2cb3a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2eae6cf2cc1cf5ba3b3ab65cd5906fb76d9398f4221cb75f2dab992a56cd801061ede9a84fc499fc32cc970057dcca3b92c4a16a25e3deccd5e74704ef8cbc1f78b0254d31f8cfeacb2fd63548e486c134379d511fd3c904fb4351670744b3f7f170f6686706caae28998820878d472baa00294718b96352d0f9e788cc0b5b0d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h64c91435912178d069f5cbc6aa7b81bc1f15697faa18303c464ba1e5b649d3a823e9c418f660b41e3039ef1ad44a80564bf690653ccfbf9077e16b6855f8a9787de4634d3da840b2129c89fc896788cc200fcdb63f1211975b7f8f12f3a56f37744f48310899bcaada550880d8a181764c64b97716b7d0ac659943b251eabb8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcac81fa609858a34db6580b1d232e324b158020db63f831ce535cd5b987650a117a04d3465b7404068698621db804bd7006f1a2d2b358930d4b67190f3fb53f3067db64918309fecc72a28bc50f6a9385068d4e3181d1e3306ca8e59b3fff86e7fd21fa2df67162d9cd7ea57d4332f20aa08b24fce7ff86baaec72f522db4386;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf1f0aa1601fa7fbec0ebf4bd72252b1d94ab61dc8a9d5fbac79aafeb0b365c8efd50627d1d1c048de836ed387fdc7043376dc4010f4292cb2f77cf5d2ddb5146a1678be6e214b2b3a0be92e0810c0f966d98de07329ac78094b9433cf25ae56b054c77e1565f351d5145375462a501f96308f34788be1a2f492346e4bfeb6740;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b0276e30cb4e61b4b8a8550834385128bb17437941988c428dd02a0bda29cdae0e150714a732539e4a0a7de6679e618172c9ef3de05423c36801152a286a05ba764b5d6a55601bf2a57e4ac5ef76feb0b4e8a8aef920590402a6ce1a39ee367cfeef3142c6d8969c591da6671eeeec7aaa066534c17be636e95bdd3771a485d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb9e2cc8036ea8846757c0892317fe86eaba90f5bfcb2e9ad9e883740dfeb65e7ac074deb9e44ef397dc567d85a76b8742630b62b790c10ad670ba506bcef921aad5ff6ea59ece6a06997331a411d05ed9d9949e58ad7743be7207d7e52d648751e6490845f1b77c1ca96437232e240568b5a39377e3c0d26ebc5b1f4b54e21b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfef4910f6664185cc066293d3d28a43a591dc31bed3b1940ff547fbb05efa048c8bc28a8e7cf56715d64b6cd2a419283e20ac93b7947063c6f8d4c4d468f933b59958277e4676c0979bf90392c08efb6ab1d8689dcd85ef5a10ce58f6d17845c1a5e31b5d2e06abaa6baafe65ba7407bc40f99252ddc831d3dceaa576b4e3731;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h647e7320c30892b354bc316e2426591b98499ec2a03cc1db58690c4b36de15527fb75d77ce20881864477c7ae31119f218b90b58d0101d87ef9f15ab3a7a9d8d16ea0adc81fcf7d77cc565cd9e725b2df0211103698282f6b5a3c76b0e4fe1a1db9434936a03671cbb79029de46c7ae6cf18b2a38d177758c0f563bb71ea7c0b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5c5ad4a6de74d57ec5bcdf794d75bb3ec4800a5eb2d47d7d6356fb29cc4c207b602d01af4dd8d5e47124c8e10dea5d08f842a98b51cc922fcaf44d7e5570cb562694a850eb26e4ca780cece347f9fa3b8ed14d793d921037500d54e724659e04f0f72416b18eef6ece2f1ed15bb72a264ebf541d964a0c4ab63e6680336d4bb2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h54b73828c47988b0b33efe34b2c1debe37b66260c50e821d91e9d88e1a9e1766883f460d5441cca2db593711f5a5723badbb516160e052bd49ea56e5cf58999a29ca9f8f54e1bf2363a6f2e01c4b529a833f073c1e6fd04239e13ae2333c7fa50bcf30de8bb004c43dc1ff97abc9db993044382480773b8e41dca1c9ab3aa6fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd424c42110a6bf0b649634c08b746e89385775fdf39772c9ea0151a23a2a714148ecc4394218814c3d894f8f6a7d0bbc0f0df040e4d86809324c59d8b90da68046fc3720df6cbe7b9e784a751a6216bc6dd9f1fa57654a6f7b148ca20684a75418dfb0ee0a5576531bef7da74712f23d031a37330f206cf9405f58da261af61;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1c6357ec471e090858109d8591c6b1549d43e5d513731636de4d8865e9484ab35ae7b07bd5f2238f84af07450bfe5ddb21a65a74b707e1306ccf07dde153085085ad1a1080be5824504c4544aec57a54b9e3b0c7256a605196423df4d023e67ee6d039c38c80d67a020ecaa672a9b1c689e779184e5fc83770275b2b331d2ff1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda45f17918b3404577866e362b0ac48bf0f7b4658238412e20f7adc713ee92232cf349e1698d0462f457f6254b16c8ddd06736dd2306feeca0772bbbce216ae1db5c417a7a6483de188f64587cccb77182733cb8d095b2b2878b92eb920ca03793c2e2018839e2472b1fa318c7c608356023819ec20866965a041658c94493b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha3007f5864ec4da3ffc6abf6c061bf74816c2cf53c62095c10c645f0911d0c5f258bb13cf238e2e686a95f75195b3a28e8f0b8f8e239e7263eed57df3ad6e0d87e284a716e93fb517c42af52974b4697595ad4ebd88a0b4a5bafd882eca9a97d31c7d774efe5230753ac8b70d17692a22708dc6f659a30ae08bbba30af4a6ed5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1dd67afe4d7cae1d10c7f4a3c5e08cfc3646258d7c15fb055b4eb875a2eaaa087c52667842ddbaf1e97ed2b609957f12d73c93c44227798721f59aad1978cbf6291ea74c9dced3503794e7f3ae790290044168814d39726deb0db50d6e0d21132b1775a35cfab1f2d295a28288cfb3955434c4e210887d571f7e5b3c9b2ca834;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b0cd9c51ed42abe7ea205a0cca994d63c0f56dbb285e54859a956336feea083d59300203b925d1574832c29cc6c989649139af83297379834225f836e4a904c7aee78807f93618040b4c2f55e5745e79c85065faaa3d2f576976d9bacb3f3ee281357054988265d917da197177a6b8421557b7b5284ec94897f4a3d82fc4297;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haad839c19128463c27186d1e0f2e1c6eaa437ee508ee8ecff05050f14240591e6eb8764ac4bfb7afc72eb790c9046bdae723045d956f518afb76c91bf2f20c07de104b83da17e633317fcb70a03dcf683be13ec4eb09cb7dcf192a3a6dfce4fe9ce4ddf17a8c12cb81423cd82501e888d928f214a53fe5325be1b14dee7ebef3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha49a1edafb4918da7a1912de83b1407029e8514445d4020aca5f6cece98938829dcbe45fc14ee12ee324fb46ef3a01b6a2fdf5ba1a55f5707fa12e902c3a7c250a757fd0863ac96357cbede753f2859721e805a92ac0c5c67645815c8bf031040ba5e054508c227abc25f8e547f17cc6f1ccb6285bcefd32aabda4688f22eeef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h78bb58f72aa300ba86ea6c8c7f9079f18e8ee75d72c20d5b29f4be3356b9eb6247c81bd030987ef83f7a154e5b417faa7982bf575bbc2ea4f0d803091b63b155ac56dbf710db811e68706c95f9ddc67e045b790fffd784cff4d6a37d008c4f6ab09985007911e8350006e940bd2c2aa11d35ac060eba2478a280326d5c88a4d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1fe09dc32a31cb422cbb650e0938c472348861609173310e43ed8c2118fea7f61c879bc0d393c25ddb77f25a709b6f025cc1a9bfdca29854110dc105335e44ee48a4be93dcf017a0fad1c09842d5e67851c4706d44c6f72fde88692c5987f8a1063f4946ddc7b745654dd59a70b9b54dac0a5fc101862399c141fff75875bd73;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2b7d477e1bf407935d9ec31e240f1b5e046cd0aeac4638073d227942f57a4942c8a99e0ce27cdb310f1a1c3fedc99a7b78018cab2d14f88130000654fb4e416c3901610924d87e90d3ffc063438b134f307d6ebfb4a870392183aa7cd6d87b1eec768fe0bc9a6a21a5af905646e5793b5f79814ef2138006704f4efa953f6f85;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9b44fe53efa42a35c53ff41f77b71043010f6aa420554715cb7cacda24e6de7d922e7b9df13feeb8f4a18963134a38d4037ac1fc909015f7fa53c1461789ac0e18d6594c293ae5f7a19183c43ce608b9d3b9ffcad83e2805ca5ebbc05d71cb072912ccd62c51284327b933e1276b80ba748086d670fc90d92c8fb723be251307;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5f35c77a3ecb1efa9a27f13c0749198f06022826cdd9f84d6a893a4798247b77a6b24f1f7646cc2309b63113b34e23f929c6c5782d7d40766f5c8a4565661093baa8d1ba439944eb8296af5aba176f00736863f5d09efcfcb8ef71a384befb1b1c46d54bb4dface17850d943fdec2906eb908b05e5f2817da68ed4964f665cb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5412f8ebb4dab5f105da88db6fcd57b62861d28be529e26b921cf634f4890fc2d28803ea61ffb75bdfbcd2c4798faebe9923def23ec70308c3c68439e64364d768492f2552b93c539fb22500ac2e03734b4ca1442bbd2bf13a7616ef5cc87efdab966379100ea3d3a66285aa130bc9836c4601b9182bfd6034004cc3e6c01643;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c300c31927f2298aa3753e64d8ba2c8a5c42e6ced0aa3f3a3753171c3de73c470aaafa21c881bc4066f76902d4a25c5d7f53e3e32986a8f1e9442d8430f2421ea19bcc639933da7385cba478e77a4ea27413b9736d083f18780d7e491f2ca1b10eb6882bbecd7cb5e7504846a0e165b2419f53081cc0c6fb24b92f7dea271b8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h36334435db6b4a0c1ac45652dd402d7981af8813de0a8285aaa8025586ddd983ddd9950c3786c8abf607355e5d3a961525fc4dbaa0fad7f1d6d51e82bad3a223f379eaa7fa54ea705dcbabae2dd2b3de352838dbc2709a05641f024cc9c8fa69e3312fdadf86aff2b0e954a54f31740746d34d6b004ee106885949f146b9e1dc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5097ee7ca95f3444e1e351589ed8c874a7f6aadc488896d075afaa0530418b86ec7712d22de61c4f4666676d8e349cb5ce09bb99db254b3ccfbcc528050481fb239dfb9acc8534c6f819512eaed2a3dc8244f190607bfbdaf4f14225c0f233a4bb430cb60d468ac7601b50b984037289d732821db58fee70d373f30bdb76d44;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he134b02ddd882d9060950e2aa0834474b4236c05b4d6f4b022c8b64be573f3d1460fe8a54fd3d4380e1ca9ec2b09126fe6a93cf70ded8edc1e595ed02cfbfb8a07fdde11e851d139b6ed7eb6557bbb8869c4eabb62056b64f2eb488a571672ab7f2016d4a4616c2f6a5541b16977bf8a351ce08c4646c6a6439d5f30a7e3653c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'haa65b099faae21edde84b3f5108f24463bc5a4efefa42dc398655500df4168b06c72adf8cbd97e86413a40fe6bdee8d2445978a8d8c7002dac9afee577a4b1f0838d56fb08883af75fbfd889c0020f65d997d3a5c392245e55d99f421209a375abdbbcb1bd815b9439672362095cb960ee95c5accf8baaa6a4e4c12e663f076;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2387159aa42ff7470e58a535b89e6f545122e9651dad3f93ef94015fcae1468ff626661950e0aa5f7a9719fed2b519743587ac6291d3162270f222295fe6663045df8b35909b041ea12ab05e5a6d47194a75be395f11f66fe89070ee243e8ecaad48fc84d4793c41cf302640a581261b1103723b5e5f97d71d5589ee161fce3d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h74868a5051b4bed3772e94dbe5a085e3285e44dc68a19db05e344c6438fa54dfa6e431d3ae46f81b23509d519bc8cca23e8c4e5fb3f19ec6c45fbe25838bf88b8eeb93bd8aa11f8a5adc60d712957077b156f3b662b8e13f39cebe28df45d45630b65bebb1e9c93e4287c4f5a10581d44c7d47e0e9cd71745af5bdfcdb9a7005;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha68bb0248c7d68cd7e8ce25dfd06fcbc280add6486dc24f5e3d008839edbbe02c331edda770b5820fab161505017479b2b3b33f653d6a4833ee526110363235b553aa9b111503030305c6292a9e664ded4a54b2fd89a8613162208d68bf69e9040ee0332e7a3d93d3af48fb7814e73726a22a4b6a197d7bbf74f119d2f52110c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h15ea67f1e9450d657dd6e29ba5c7531ecd5884fd29827dc908c84520d5b704f4b634d65f54f38545f8084f8b97900cc8a075cfa2999fadb51ba0760b75bb7c3b44498fea98a5013c94a75dd0355daa437bb7be5d6f9c7ca6933dd991b1d6e7d79237c90ddac35426e85e3bc7d8bbc5a2a08aff3ae173cd8db7e373938775ebc6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h229b983a73b92039a07d62698d8ccdf7e076ee303fed66bd1535957781cd61d8f49c3cef34b052e30848426f1059e784ab90ff3a5794882db7d14937cc855351c3324115a19e1791ba838fecfb87fb1c2b4b7f506c548dbe005333369126570f2a5c0e5c954d41a3c808e9d1004e3b8ee36e887d80a9b4d8698e0e2ff25fb11f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6355b21c8b37955f08141f0d9b787e3b9e57559de891f02986740a0a50fbcade5854fad39e501810144085520a7436b38a230ed6bec750364722edd0d17b2bb11bce220af9448da181e003560deb6cd020684291b0854cea821a2436bfe012d7784322e3ebf76a7688ec8f682d321d8628a94320766b5e3f305a835b8474c91b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9bd01146885c141899c2fbd9da8cf4cd32b2abdc7fee639dfd21263cf3ab67653fb1757521037ac0fa96bd76140c005675632f9cb16c0efd91deb478b6145f8f2ef85c00f74e752a7a49b302868649d62869f5bd9324d9db24b0b39a13c06884aad543f0719c82267cb6d847e5cf50a16a39bac4ff2d5edc8e59ecf281acf47;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb89ac8f947ea7caa3eb8e2bd79a95eb3a18ea9eb55f3bca03cc6d75f87703a52ddea69f55b555d77b98e8ba90de03fbde706e4c31fa962b62f95d0eba5b7a58b18f6a59541093c401cda4b194e234cdd0e565e3948769f45698ba6d0e2706ecb30e77bca3c5fff2da9e3b6d6d0c64b32ed286d7f8fbc0be68720fcf039186cc8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e854d5986fb5fabe4a7190cb7f75543ec8857c02c092caa682bfc12d49da692a67b84dbd172be28f483a3000f9b1fa906f895c5850a1179e4e64e12a36a0f898bfa03c06e4d0a83161cf86a827546ba11cef54826cac9fa9f8eab2789abbc84fe1cef8ee47f174f562d7e9de86b98b42b20715d4d0d5d9158ed7d04c8da7621;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6bc54ea4005ecb69c0cfb3f8e47b674605b2dc688db0f68c3ad40126c0df4fd9c86f030af7ccf9c8de9ccff2a7ec08098bb93966966bf30850e930ce566fca670c7c981d708d1550af53566c574a58b88310c27e973a2873364cba457a24e81f68c5e85cbe45a59e9e8a58a83a743bdf1e7c68ffae9632daf43ea06d117dea89;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h835f3436b6f799577655bc9606af9aff29da0f952688d5d0f84fdd470d6dd6026f77de4e9b539ea14c6569bea067d36ccacc838c6e766b8340a20a502eac2734e9b00f946379304735885a8d4622ff7525cf78d307d80da6290738d368a63b6659c7134c62bf1629ae4cab5a56c966ea9d46bbc5252502781bfd6531a9b22816;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9755d9872220663edba0d710507ba03f4237caf26cad9fe72776f21bcd830b629f95de641c513e70d95f07859635a03bfbd520549b4770fd29f7fd68c7cf2bf0effee6d45aa3458e0d93dd1cad87762d960df91e008c8cf8151136647a1a1da67f99f4a46891e174b2aa31a34b0de9eb74d69a5f1c8e728c95469f2fc3b810c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7efd20c0fa535f69be472ceaa70fbac9959a2a58fc3eb1fd22939309d48309bcd30e2b721d57bb86fa6b91f363c0e75ec433904cd020fba470ea3c2aedf5b70f0af4eb7ce43649cd3a85b2ded58ac1f4ac205ab168e32e34966514e8af8da33e004dbe8a66fcf65b587680a55cab261eee481cbc468dd18d4bbf0bfdb305a8d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6dde5649e6a1d283c2cfaec93747b18333bd8270d5d9ffd4f98468e60926cfb8426dfcb329a0ea82c1c9125aa36527ce7f2f5a22698a4217c435afde832909c112ea6caa07d7890e55d05cfc3ccf661cd62278f45d1a6822640e8a6061127ddd19ead3e19558c2406cc892eb888ec3235f278dd827143151297c9a5503d01b2a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h744a6f469d65cb0189ba60bcefd8cc46769267d746eaf17fee7a4ab41be015c5d0da2a48edfe7466aac7060ec4753b068a784577f5e9e33add4c79c838b0866135e6b5622b9d42bcffa0f8253e472ae2b94aaa1542cddfa43849db164ff9bfc346ff0714de340660b5eb4288e241451c5e9c9f848c9dc6886e03f053020cfcc1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2a235126cdc6729decfbf3da51d05cb72974b929204e49fcb18105d8bdefb863b70ef5b2ac92646f6b8f82e6b9ff94642b65b0f9865289d404e233d29107029b5b738553a64bc87b9ef979a718c3520c212f75b03ce19cc4c970cb0f32900809cad99885422f59ba67f392b3a387639b6da4f33b1ffb4f6163f4384cae34bbf5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a886549a915e2c27b90756ee1d165bef68799bcb12b4014bf3e53a96869590663ffbf44dce739828d9078ec3653b118de3541ffa658e671b2c16bfad01fd8f1ef68e0a4a732558214d7b25ebd7b3af79bcd65ce01cfb73b116cb157a7a2273aa7ef6c3b568bde906314ed22739ff551766ec8b4859b41e229ccb0f879239aa2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8856dfacfbdccacfa81a014b85c71e32adab4b98ab4bab6ffec3040675183bcd0e6b218bfad0208f364ac950437da79d2a60871b91bb8773a5b175ba1d7499378a37ebe4bf876b237a90c984ea7ad3cba5d5014173e79c5aa7dfd3e04f288c1cd438cca9845679b530c92b191435c9aaae30a061ae77ef10ddd7147d34f47a6c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he6493d18e401848ad79dc229b4deafd19f6d5820fab7049ca172e8e745ad86509db288a515be21c35d77f6e04f1e5aa1cec273e92f048fd08f8ded9a9b30b5e12e5b4b313f485816fb9aa388e650b6edce73e56d7eccd75472c9b945983e043e52601e1e99fadc9718f2d3a32c68840a48705ddcb56bd2e0c0d2ff171a009e48;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h77d203669b8d4ff9125fa8eeb5c740a57cf6b482546dc9150911c6177a30220823a48ada4205d2795e76d4812b08aeb20855d8469685fb3ca9d07f0e0f8ad5291482400633b01c0943f86ce7e778113ef5262fd9fa5684316708a4f5b297f256956d2c5ff713edc5f0ed49937297eaa337527f524abb4901202d1cd05c59f124;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a16076f3945b09dc873e1bdaa20bc62d0c944a39eb0d2fbd5ff2a7062baf8a5f457ffd513e7de9155186754784312f1d7221a196b894a7a565e5583f292b4406dc41e6e22d49b6cb72f972f567f119e108974b2d3bddc64bf4fdfda3c32787d75281c0f798882600b0493e7f14a2a32cfcf1525514e8f10c9d622d0f75431c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1b6a820ed9e3700fc97c50f6d92b2ac3736f633bee9d393bd8e89d98b85cb2120089a06d895703ec127b2a90272bbba32a68bc945e41e88746e76b1730f50079d266bf89e6fac5de7970e72f7383b6c1d8ef3a1a8d9f0c4d73c8d3816cec083f619365b95099e522607ee163aff08809c77f116fb6e133462e7171086486d86e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b593e8267967d2018bfb1d28f4e751be2f77b86aafa794e21af7c3b65e96dfb00e154416163e5dff4471f7441569b867e16bcfe977c6f6b8ddcd7d41bc968b22654cffbf67cf368b56fcc27dfe0dd9bb8fccabe49f2825ab72e4c63b2dd869aa33a3603a6caee49233079c1e5a3f9864dd4d6837553f30eff519310055d5b0a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4582ed69350443cff2db8418a459124d3bd5442270279f11e24bdabd343efdb3b69f9c9ebc762b2ad4d40326402482bea7efeddb406aa7b2b660c52af61ee73a748fcb5d65fe3415122376ee246026c867001418b0fbc42ee0f678340cfc2a1e9ab3172d6af004504271955c244bd901a905c968803d4e9f9cf952a98db040d0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hea085b4975e33f5ef60f584315726fdd8052474c99117256a3347b9afd67f0f571eb25896a962a943a39b99f29716d4584f52f381a2f88adf4fceb4b437fb1b927f4fad254fbd77256dd9b21729bbb9d856775b03436f2c48fdc39f5787ccb551a9fb3cbabfcc064f594b9f8683c9581c8bfd7400d66819dc98b2bd75135237d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc37e83549dbdcf8cb5ba007860f7e3cec5107949a6ef25400d8dbe7e00bc77d4c58845625fb806d567172118fd53bfdce5740785923e2e41398b1adcf70f6287e76462fb09739d685bdef62606c0a956638cb98f747167ce80de77dc230934b4f6b1ebd9a5033cbbe5dcbccb4b428eb8b5b263b2a146bb8be42df968ac5517;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h88ede38855ebde4a521a0dfd4376f7760f348edb000bc2afedded364e436be0fd1c506132fe63aaece3d06145bd1d59d9b24d8938ada4c06bf25db4972b92db896a7b238faeeb43c0bfddb477a30678abc9e5fc779720f39cc6fc190e9f779e1105ad53a7c2998d977626c0a4d25843f6f6b1522c3c3bd48c7bad4857f8f8fdf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h61feece52e3f30cb63ecb29b2bbeb7fd16e5bddebfc32cb088f241910f3129071ac340a5c6cc26986b46a04627701f2053cb98fc9b712e3a81857e99364068ea2ce6d0c31187e038c1b606d62facafffca054038e9d196adaeaed0b1863ecdbc44861545ce8255ba05c94fd1c89d5b18caa97abf5ff8b7a8bfb389d9b95cd4ea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2488a9eecfa2ee53d97532ef30093cb5d725fd130e3e08f1fb998a17ecf403a4699aa676392501a0f9d910e50a293f0232e77d6cbace5729bfaee56abba43b316ddac7f092ded08d726759590ff4e8c966d91241ae7d2cac7419e8787368d1c24933a5c8a2411f9521ccf8152c8ec160b4579bf655a4e1039f9b2edbbdde055d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7c806ec312d803cec3e482572bd15b6cf32cea60f4fdc0949b7afe05c953e76ee1b1c205fa2cec541b45a4b96e2c589fc62fb56ecaf5b81e782eb637e05f58934ed077582a4342d019f0d936bc0e53978b93f320da94ca96cba787a532f8dfada88723f25ed0faeb38c148b7b3ee2095f30c9d3f5c161ab7eb2f55c34999d24;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he9622e2a54f0461589ead046f6a28f049f2136d0523a122de34327a1336318db50f0f112547d72ed243c39ae9b05aa684f23a5ce7cfb0ae32282b90ab9222e3aee714a60f2cdfe82960d8e549772b258f0ad43eaef94964df2fba1c0ad01bfcee00f25590b838b2f1316f0651f12fb32610b980f2e8afb8bb24d086414bf6038;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c5020087363d735d425dc70fa07cdab08ea5787b40507e760bf69343251542dbfe5249d2aa7b5ce87b916b9748004d5554e89ec0bbf709a095be30b852d50c69ea0a57a9d6c74df7c7f74001f29d2f2f67090f652f562861ec0ee98c40e622cfeaebf14800d57b6ba079980e1c38056def456d4fc591adc85c4fb9194722398;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd58739e18361ebdf44daee032e5fb49815a58be035d061490579274ea2124a216933136abe1c653e7891daaa9377e4088482e5d8d335cd55b703b40d568f09b8ecd9212019668d5916b7af29103b273360d9faa7fb1dde331f6c925610f7f6e61f1ed3decf138b62d6466caf6679caa4cd61ad8cc923ac394e9ee1813e7fe55;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3b5f8d744da0297aeefdf54ee273232795da66b46ba4a5b46e8b4c48bac4b420187bf6e23fcdf3bf48d55b937c26073108b564b996414323649471f162535efd7b9391b4aa67b52817aef9a2381172d0e1e17ac0370e1c9dbaa85f0d495c7c0e14b10b747a42b6e5cc7b5802f308ef1b883c91f7fcd38c580dcd3fb147bd957e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h476c5df09a83f9269bef27e8f22d53c1f2a300fb2ab049ffd31087848a480386443ffa315738098b5ec960c15da3e401f5637c1b3af5a20b95a237357461e3dab283916f8346b367b8737b51b4c70c51c9ef74a68f0d2af9f3393250eff90376d83e97a1be10c40827b1f3cff1ba2060f8000db2262c14845600aef41394913b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8fbeee2acfd2493f87fb1cc40ff682e33204f5d22eb0824e415a1b736fcca0ee056a5c4d100f69bf6e82bb45639a402a205b382f49775455b2b134314754f60290fa1394d062288f879deb45dd36aa32ea34674692d9e5bfc72233d4a6e62ed9f06bb41b0d48dfcdd9914fd0d665362d61c2d2b14ac27823e9561673b0cc282d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4bfc3f08753c9cd92ae93504f2e4f5e5a2d192dbe831305e7335178fa664f7be58542c35b52e306eb4777f687a07b850972f1400378ee9782d1dcc7f4d6548e0f553ab8dd7d67622d4ce0a83e97187160c043191665009044bedd60bfe24d565a6b9a81bc84f942d550c37c4e4aec707e3ceacd155c0921d511075d95d00948c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7b374581e3b9f3486f6925b86286db29a42cf34cbc02a3e4bdad513d9630484fd7ac7a3f52a28237ae094f39e97edc66ac5b3cb7683e65d6b56f6c6a92d951edf66d879fd2d2f896442353fd28c5bae4be50d23a1ea69f07d3964611bfc800b06706205ecb21c48a92bb2df9ea08f7aeda01e169a0d79555b6bb383c84f2f82c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h968242143e708f0e1f4adbe1a05b4c14170b41169114b11e84c1b2a461f9c6707003344fa4ed67a4ba1b44abc0abcd56df2fb64fd17a31f1f002a7fd85de824512448935acc4c364d973a65130c652bc2d1e97e92ff218e21541ab21db40ac865a1f9ad643af7dc9b9e7bb979ea4919b1f45a54de731293720d2c39d18ce612;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1bf6aae9295006389bfc5956483285d7a63fc218130594236c070e4b334149f72db415b5e763c97fa837234862665322a500f15b3d07ed2656d31a76be4fdeaf007d4d0dafc385899bd59284e4e0aa32806e8b643cb489119913cd074b396ed0e35771a4139c0f1a3890435dbbeef5996f1d5bb27875d9abe88fcc6ed8d3abdf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heabe0130deabb2b27153dccaffec637cd0064f8facb5084df84430636530899abff9c2ad8e876f41c49fd5d8660028d11ee0e07c11c40ea9b27d68b41b6bcf9ae3967431cbe851f49e3d4a157597abbc30d9fb7301f8e0de80dc73db78c4399a4aa3d35b2c66552df1269722bbb2d067a5f132861a769e50c8e23cfc796cc32d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha91912813c1891d00211c0d66842bc2d3e47ee7daab8b007c0eacec332482dd20ca4e9a278aac706016c1535606489bfd43c3df5c59efa3e14c783fe2826f913fa1d8b864774c184b6bdabd5386c0401b557adc314795ae7bcf130ee63fbabb3d71a94e7ea2d9fd042552158f4bc9d64515b630d0a57f24a1a0ba64ead1d7d2b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h683e504780b5c5649e841ff60ad3d1ebd6270bdeaf73c105338e5acfb7839cc97f7ff4d63e7b0c6873808bed54f9dfc301befd7a04860a7201bd03ee3ee712462df00e24218b267e00cc6110cfcbb5fd96ef020a2a3465a45e700b25196b3b40bbd052fa1a2d64614a59ab32780e8c80cf466476604351935ec8f84b9310894f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde57b27fe3375177d2a92d5b3c0b817a910bd9a5296d9c11d9df47fdeedebb9bf9ff30db789acf5367e4316085a12c4ba47776cf58c1c1bb008961f999e4e113bf831f9996ad9763e6dbfd2ecfb0f777803126b8f8b240f2fe27cd6f04787d0f840c9baecca82b4f88bf92075ce57391cbf03e271339feda51249cc63f638275;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h73e058e4b8eb70548ed59879fa9b44ebd24d482f6a8d3809842190edff75c11fc7a721ff6790fdf70981b8a081258b3bfd0b2bc5ca1f9c17b871d2d7990519a6cf754ac813f757adc6fef8c5eceb79587f1e1d37191574df5f05373d168fd05fd73dd19b8d74420b3edf0ac48475d8f23c943b69f8b3bf8cb3751a0283c299fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha6e7f9926244fddeeccedae6d9dbfaab816ecb92da979ef08cf9c35ae15fcb25ac25664b5973e3ca2fb5bd8ef6f2dfc19d92a10cf3fdcd16294b8bb4f05ca91897e0be137cf47ee87c63b8e2924612965a7d4e207a91a6457dbfafa44e15969e477bbdeb97aea36ec82039f1dead768e8cf5cd7f880fea2103d5b985acd49b5b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6e7e49134114c8c23b36aa9e8b11d6162a264c60b87620eced4817f0b089d340d05ca8bc2263f2e2aa9f8a7277592efecbf81f7f4bc61e353e75ee4457430f163f78a6c34f715802f96a514f7fa0147db9c7ccba7ca0b992d6116635d01587d5894181d31d2f21628a215fc174ac52f3f4ba277dd1888c6baa728ae1c0875913;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hec36069eda5fb71475c6d1d147b03e6f566e440a36ce85a04c71843c629c93a958433077853af1bcfb455b240f32e804664b255ab661cf7058300766e5826c96ea566020721f9ed2278ce1143994c7da5d069d04a880bc4b87cf5256f4677645714e1ab11a73573e6999d084167196a461026a31fa38210d3d7bada4f00ff026;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb23f5110324c52ff67e611bbe2a971342d204ef137d45984ab7f1a743eb70637a0cc574d94e5f96df1d31d3c9b00549f24b3af046ba2ac0442d4f796fb20d05bb12082002f46dc582fb1fed8fa3854367d87fa31556b025710b841704c9c36d6bfaaa2195b7da175c39b657a82a541de6d25b2d18cf5a50cf59eaa88661ded51;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5094460bf64e2f2ed0e74a3927ed71abae68ee4cfae0b5006d7e4e7e7e84218fa061ac6e84a10c9dbe5ced25e4d3feb3ceb456f3cff7dbeee4bb18007057b7d9de8a302443a34e4bb457178d6a063a034351b5153e3565444b3700380091a2805ebb43a200d6c784d913e9749435c46812b3f94f120b68b67e88d15d08598dac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf8abc58292dee8bee391253e706141e6da96b819bbbf6bec5a0780c79f7b9590f7b3131e27c2e4664f344cc4d0ae23ed0990c035c1664b3a4fc46d6e5ddc31ade04732bf0ba8b64acf64be0efcdb01a6b251886d77292cf10b3d1689af51d70916cbd8ea9ac9bd4b93bcea1462da4a729bbf28c8b90e2e3b9c9279618b3c1b25;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5b20ee21b5568f4d089bbeb6437698fa71e3f96b5d434b58c5551613a76db7488eab665fffbfe37ad878bdeab84d9aa57c7655e941d8e5ab4508809b15b5fbb8516f51914dc5ec056dc40338f7d9ceeb12d1119abc7d197a1d6871d9cfa26c4173df356d48a4cb2ddf425e896b0de0c8c35059422dddbdc5b9e82d46cbc0f948;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7e25a3a432a664bb9660313c36a2556aa254be2265a63485df77e8903941119b690eb3b5bdf713583778ca9e166a31fe6274f8dab10d6a200892c5976deb83a7ca6ce18da173ea6d74ea2fc2725a440ff37e5f224a28d8423cc5030c5932aa691ec409e2d60298823908f0db1f9eb70da8e4c9db765814024c95ca7594754a84;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2ab57e2d0a1595afae351cda2ec19364c93c587e4c53bfe00a55f5a7f2fb84c2b557f62a2f7658e8cd597cae8fd3af3387cd77cd0feeebf76bab0b599ccb072cf7147961366f4bba81a43f8579cbec4a718ac7d6d91460a26dc366a17f2c43d06d626f9caf9e6090285b37723f087050610385b549ddcb7512b6bec0a41888ef;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd2af3c312b5751b89a7a38c6e7e312b31b92756809ec3f0887602e10c690aa595db0e3a2771a318ddb49ac7966e3c76ceb42cb578a0a30e199c1fc2dd2a392ebe05350fbe6c77b63fd7e0c17ccc1736c61c03ca3d6516d7af0f21f98fdd2aa0581184681c1333a28c8b8589897d1575032f452b84c9356221404059869ab3fc4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc89470ad156a3c6e5409f1fa316ca83e63b0bf8ce512781f47b738b2fc1b80dc6deeaf97f077cffeb849b4671ec6b031ccda760d37b2d4bcd9a4425ad7e322174804b674901199fbf1b081a15fae506e17cbccde71735cdee313b6c1cb365ae772ae8a8cac257ef5ae040310198b78837154557c13823574e682ca2d02b13406;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1ac23bdb19bafa29235fa6952bff6b29adb75c2929fefab96b0eea1cc457dd8e0c2cb3232143aca0cc13b8cf6f19a8df029192245814da4deb7a02b7a52bea146cf764225d6e7e7073ade780dde2822d5e856557d86ce9abf1d7e351f925725c4d52329434b7271af7c7c42cef23c0a3478c89375776898c90fd73ca0a0be98c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h392a796b155b896648e140bad6aa6479ca4f01fe86d61cef44969e98968fff2904402e6694a8bd46f3f8b56ad5fbfbfbd7fe36fac9318fd94578eced35713cdc2b7491b7793d915809ca95f40f58193969f0e970af5ec8c59fe4a9f33550a99bd54e22cc2d8f67177a04376748965eae2f9b3e44ebd357a7448e324b591df678;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdfdd9da9940237ae677f26d3ae3744db99b80d83471f9dc22e12ed81b1079301b4349c31b36a2d130a61670c57822c10821877dca3e0d2252534a075002ae848112d24fbb36618a3557c99d8d22945e28a4b2899cc50363e4da5b049e20b1392feca07e3e3553670738a299af91cfdfe02c53a808469652187c83ab7ae626855;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h143d85cd60ab13e68edf52e222ff0e415ed8316abd624203f54337a9f6d0d7b0e836271d190a2d4922a042bcee35403d28899cd33157db34ecbfb469c0b1375eb2bb063d10dda16bd7c3f4fc5afa163dc67ecb1dfd638347109380f63bfb57fe6cbf99544d75a175c5f365f728b8d1e79f9c8e50c2d5898434477d2019516cc2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbf877026a906763a5a545c2b2f16757c204832f783f20d31dc0a1928801eb2c8afc26c142cdfd06c43da53e693074aa00776b809c6a98a75ef56bc88b57edb31a34242946bcd518829af825ac7542294f55cca20217944291dce60f8be2bacfbbf53743ed2cc6700dc2800a8263c1d707e0908601bc595452f34a57b01032f37;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98f075934f47aebc5673d7b51855a651748f7f3c547ffd7c36e05640e084346cccc1833b82e39d7656887e2df48d41279f2c99d57597e055742bcaa626e1c97259dd3463a430f5dc86308ca870c47a71ab2739b68aa5ed8e98baf7e689ca807fa8fcb4fa15cc359c592d0c74abf06fcd086a3f3b2345a7fc4bac4cab1e2725d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12625c9f120201a71c862099a465b4fabf9d9084bfccec796f5e987516ba6489fd961f773b7a51139a132b5c2f9324d132f8d7bc39889a18f98e20ec3b1cb3cbf9f6b68d9be68d689a98dfe140a0d5d32bad42800fdc502922edcfc8795b579d91cfba9e5d500706f8fb14ae8d011b7a52726649f603ada208cb0a017c3bba24;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8278bf028c4f8ad9701cd1f82f1e99d10d023ccaa450a8b72ac9cfd316f76cdda16469ea57978ee848f02e9ad5cc97dd1a131c4161dbdfbd1ef92dee38b398f66263cfe39d064da49fa1b45feab0f503d86a6f34163d96ecdc81a88c596d093228f81b40a0070c3f857219df25bcc9515b11943942378f94cb95a96954d8ceed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2cbbeba1e5ce4dcd0bbc8aefce93dcbcbe5d02b31d7315d4da82b0b118a1cbc6692edf2784c58749f9c6b75b174eb99e12977fb413c93c26b349cf1e5f6b2a2472f62e6dcf930e969a3d168d6bbca070f82f391a0e556531557415c240df38da9992f47c3825db5f0e10338b0363cdd467aaa5f3d3ac76aea95b53f071c9933;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h24937a0510ed08044b8099d4148e140003abb4f64d465a5095134a0c70998983448dd3afcd2579bdf1b85448b9420972abbe568cf13b7f3987bf3497945a857447c9be4c50d2c0544f1fd94f7f0353215852b9d570f2731f025776616fee6b71ffab74fa02a63631d8a362672c16d592128668c470065971daf71e91ba3d1214;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdc31fe4b507d641f48421d65767fe4992ac3f27a54bd11b7cb3d0e5b1dd1aabba3621a34b1f358c6fa4b1f9df16a988a2e90b518822d59a371f5d430bbf20eea071f368f8cca53f0c7d6225d2c2280ac9f24028ef36102a0ae304e261342a14c27b69266820833e27025a3a87d0e6070933a988088d57b1c13c836b9dec89fda;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4f3eb3a9d3f93e073c2184378f609b9272358a9e9bc5e8b65341e9a7ec6f99dcc23e65830b7fec919abab389acf2d5cd3dac5543b8d14f228771b500f3e9d7276d2c58d208022fce1833610228047f20926f6a7f7b1300e70c990f9f473da19fbc42136f11992b4786e8d314e75e103a843f46738b0246958c20c4e475fb4dfd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc3ec49faff52d479008d3e0ded598fd8fbd3d53cc3fcb88bf21305ea9670d60d97d9eeca52c72f52d6dd12a2b6371b71ed99e5d4e7e5e969c6e3ad3c708dc2c8eaed7fa45348fc191f6ce3deac7533f389011d0c974229576183b666461607a4cc2d681a4fbaa2822855998aebc457f5da15cc49ed085e7f3f0ded472cb36494;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3416f80bdeed215afd1495635c7b56e4319c769a6180c92130cedafbec7a5c927f0f977e708093090e7bf22bc0048f989a7e03b031ecd707a235fc0d3b831e94992d5cf2d4cf54776a1bcb355451bd30c4c7b2bcee3a2570b0faed804dfb121e12b946ef41efaaf0ac783f04bab3371c953e55bb71148fb927c00c9c97bb622;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb576e6f01e978622ae22b2fc9133b8152c70d6769bd2b440e2505ef210b3f348ed43d02f4dc7173be98d5a72886ed116fc1620e403238ae39e9187ab37a2c6829c226a7a8ece4adbfb330c5af70daca0978e1098ae27feb2baf44d7e63ba77be8a8139cb5701d009f944372f1300debb63cc699c6848b54dba061f12b86e5044;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha91616fdc667978af798d00c3a3ec0755e1aa408b582d4c141b445df8bd504b445cb3c916872b45f2424e14af02ff347b4b2fa3e05afce720ea5bc45a53d6e9591e62737b4dc066e069cd90afd2a2ec0aafcec1025320ed867e294f3a10f8416b53af2035f0de7bc4fa5fc8dc9f2463769cfac42f12784c300e212cb3284ffaa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha5fde9f047e58cced0a58ed1213e347977e0f1171a9b8240aca0e9b729f54d84c09aee82d655a6297d3abae62b8ad32f0d60ae7513a405164293c4e82c567e1de6d05030b32ec61313de8fd073e6e3d6b93b5dc64e1631a0b3114ba3bd2871261a46ab5eefb02b12463257862f2d42d7618aab5d020517bcbbb3ee81ffd7a82b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe37084783c58dcf1245b9656faa02dd8091ab28dcb42f29bef37915edca656de53aab6ffe9fb6468b11156fb0a9d64aab7e25214861b07225542cb333fb7d7f6417bf8e535528a5ca6f90a9d138686dbd1648fe6c353af78a52adc2b4b621ecc9a47af69a7f760ec2199a738c03fbe125963526731c83b6ac1b7fb06c2d2559;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbfc9cf4a938c29b241786c295ed48c52ebf28de8921ff606ad7320176316d042071c0bd33ccb1cbd41b4fe88b7af5de24ab2aa41ecfcf371491bf38d38bd52035c73bbd5d45b2b4956710c7f41288f97ff5e90c7adf532c9ab065552ef60212fdd9f8be0c56db1bcfe1c9cded1764a75cf1d34f559b3f9941894e4f7a2e9a989;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdaea54fc851aaffddfbda4da377b175ad4d92798f325cb7799662674796d9381df2b3f060fd68499f867b56f604576afacb7f2b426e029ca3d5a97b9d1f6296d802e072f329030d01b6af81b6b02050ffc9b844a83baa80d478ed4aca02453a28bb9948402aade09f4a41f9470b5672c98fc17be37c5f848c83f7c564edcf177;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h13a16b26972269cbeb9bdeacaeb949fa42d2b267c558797b567f10c16a33ca99321843c38d672deefef74e6a8fb2df9a394ac27af5a3c70c600e0af7399fd77799e3121e2cb0cfa8130193c918f92cea52419f567f062f2c2cb2aab6ac2018253dc57765ab1911fce6b2d304d6d72e475b323de2dd439ebd92b3e2ebfb24d83b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h718a0f24163bbbbb26b6c38b78dde4b2c1132363cfd00c69624a2b736f4311b811cc7e6876748e6cf427723e1db87c105c4ce8e52cc171dc5e328571b2382559041833e6d283e836c92a498b39980fc3d6d0d5f7a9b3528cc7140e307a09b1dc1b12af4a97a4acbd80eedc81a1edb30e09edcf269b722af5b61840f9e559a6f9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcc48b91d07edb020a0d1143265b4f318b4aaee159d0df07c1a5e050bea5cb8e62261c4533f7d2b263cf8c07ce634f37cda92a217e00a3a87f7b837375690a23f9c8fb95ab005857494df1bf35e277af70f3397ff0273d2be3f095374d0b6def9a4128abc3fcb6c5e79b935b3cc3cbde7e69c669cc7cb5e12c2fec35a4d590a82;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e8647ecc22fa1d250435ae355972b87c640fb10101ca8eff6d1c6be040e5b3209f87a14f91b72027bb8a14d205294a1e6277b512857b79b67192d40abd375451e4c7b396e1ee026c5f9bf17e5d1418c2cdb11f30402f739ec3c1bac197c234fb676d09f8c200d0e015b84d68a10c233d96e2fc7169e8aa87ac99c337d867b6d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdcdce0626043434143c3b9c619e76ecf3f611ca74ec6cd15eece9695374523b36c89cc0819cc3a77c545ca56223dff78c1f3e6dd4cbc0469d03c343f56253583ba345885c6749fb374c8d11380dd147fb1dbdfbc54f49bb83fb360a40e4bf86ed0f55d037ee390962916f4b7e9ac62ca9d1b4c78f954416028266b8d0253799c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a58a7555d703b0619c3626c1cf43a62e6f1bf99c98ae11e019765f0af116c423c270582cf257f51d9e3bed341e09d3781cc7a1e3161097476d3a3c421991570d51bb8ee685241255574878fcb9bfbf3e71fc083440ec5748a79388b581a3b71828476c88205db5d41f3a09518359e9dc19441a738a0d6ccfe6981f9a7ace1c7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98853a443bdc0f5450d15854bc05c0f96a36d931a43f01e85ebe83f6f06e9acb765be429e61bed136a064f2f21359fd673efbbb63939cc10a9c31328e3db913f69c97e9ceca019ef791debf01b7311e98a2dd97e04ffcf2d611fd4844db2f98ba038f706be205a7b15fc069c740c3bff927b71909a1dbafb618c63691e30c4d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b79ebc51b82a8dbebc1a78ef0c6ea56df69e9f09bb25be508e2b1af94ac4599958416355d3f1009ba60edb59cd4f13ef3693f4eae4a9aeeb9a507d7f5ba4e3ed2b48b86b92499dd89bdf9bbd792afcf5a947256179cda324e3af6ffdf3a35982bd2bf35790b23bcbc9767a461fffe60acbddd849afae84c2c22f3976b9c8703;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6120f33bc68e83ffb49a5b650a03683d0bb02d04926397cb4599cc88fc93cdba2fbc8db67b50cd9828caa0bbe94b4e7e4bada10722b263a0908357721d453739426d65d810ab112b57ae2a10572165c274fa5289dc8370d3359f7970683fe3eb9577c1f3ac4dfb6d0a98a3e7826d825cbddcbdf71756af961142584be40e180e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc2f69c0d0861967e915302c682fa2cae89f10835c751ab6805733b8f2a0f842074ca8f41f6f1cd102ee8e9bebed356e278e9539c5f498abe56ee9300d0cc93d1b33824b5b4f6f39fd818642d3c098b020702b6ab9304843efd51c233a4ad38cffc52bbfcbc06d8275fd1c91cf5d414fbb90a058c1a340a3fd96028c8450016c5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h193ad4315b36e9f9ffafb7ad3d6fc923a001fa9353b3d4d086bb3b35e0ddbc6cfa0588abc990ae025a32378f69ae4f895b8fbe42018117be5afd832927869d50cf0c33d964908080701bf44126e48826f50ba263909012d3361d651c6d61f3696ba0965c6982a7af96e14d6c00b8b8e28e118af32e40969d1063b74c91cebbd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd4e7d81376d9572bee5db31a81e64ebeda420a61b5561dba1fbdeb02d0579b79767c6362b6f213a312c09e71fbd3396264aa9f18deeaff03bab475bb4f0e8a5efe3b41df93e94c76e9cb467be9cf03ab3b22eb7199f4479a119ab092626f09debce51a35b5147b68ad83083f1cc5a53b69666c2d45139e621ee0532767a72236;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h7c83220df2c9bb97627187cd92cbd1962fe851079dabcc52bfb9c62ea8fe08f89c9fd1d95617f5c0ec0b822212818b4662d66849985dae2e99ccbbdba8d0f269f020c97d441e7a098dee944c0b492db74594975aac9697de23ed4c2bb37a62a20b007ee727dd7adceb74cd1106e3b83684752d264a091a2a38fcba993961d3eb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h27275e0a5cb5d24d30b7440b3c70d60f26f87015b8c76e0c65203f4fa04f9a8c5cdd0e33ef7e0fe3f3950480a8b2d0f94df4de5a3b00916d2893c9662aee24d258c11accc37db297351b04fae07ebe27a90b592ca7dc913d087a6d7579ecf9957e018e81d779ad967d896c3b2a3183465974dd95e3c7c257d912d12baf5f9844;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9afafef6429805963209836807a36eab91acd7ab55e1534432531d022f6d298efeaff7253821adfc5431e6f299b706b0b748f03ae6171898649ecaec4f90b249ea5c8afc95fdb7e5d5ae6265a85c230fbd316a192bb03cf7a81acd1683364678d60f595fb38d0b06004e860a2b5a4e247dc8d361b88ef619bbce4e55d0b6677e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h70bf12f0cff72f170d0ceadf4f5edb886be8a42185c58a3caee94453ff01fbe59e6db8108065820b33682ab6ae407dfe7a5d808231b20efc02c33519d6ffd87f4d6e3baa7e357b5d81337bf302ad274f7ab1ed56c89c8c618162b3894425fb90eec5e33b6624aa63fb9edfb3eeaed1343bb9514a11ffca7b5fef30d6d144da0f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h639220e4ad9fffebbcb0491ad96168b47cd2956bf4d02749c50b102329c774a944e9925061c0abb2a4c56bd4d15571fa5f655038278f06ac47763ee3b25f2c7c2d90d97e5db46bfb7da34a6cbfbf7316d1ad4ae9a22743249c3d2723746dd4a49e02d44cae1f74f5a32f4ff36cefecbd11b182861ab913bc327d772bd44f77aa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he18a71d239bc21b41a5b5eaaaa999976d0a1e191f305908a10449405cbb3e87bfcd07c7f50f92ee5ae0b10cab578ae65ea5c9bf78e76498f40b472717d7ba3fd46f83eed8829d1db01505e4239d70a348bc6a25a38cc3ab3c19e1315b2bc81fbed760e04a232271478bbae8500b8ddd4ef425a8ac5e1da0ba6cf7d0c81ca9e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h47dd2e3c216c8deec2e63082a5c07f32cf768bc0bd2716265c338886e037762c2b7044889466b370500ee15ad41098ee5c9d4dac706e316abae54cd8af31e2926f9f37de1dd3b50ee23526760754e38ca8da663e620ba1d25bfbba6aa533c305e41bf1e410b1d74d032883b675f9d2225c8b650c173da6da2c4bd45895867db3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd7a358059afe0532f0bfbaa843b8e5d3927301b246468e2ae3ad502f927dad110d602fb51d7dc34b0e490c6de32b924962c7d43bfca91ede6fc0f1a8a77073a6e521ef649ba718bbd6d3f9e52ac262ea302b34d26afb7600100c3e1337c62f775d25f1a7e2bfb1fdf69a724206b46cefe324772a948a5628be2d07c039f8b844;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h84d75aae371c05b845d11f6fd777bf690b91186a08c068c375887de73ea99a34c7853682bbeda4c1d5566e2b873386d311cc0e794c365326dc8acdb6f44b7b6a6a148b0a050c13fe6791de8379487d5f38fc33a275caf64032ed6e570a534775bcb969b8a6987e941ede5bb3d38d13d420334996ba3fc969cc00a92cf896a336;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbc7fa7029edf522d011aefe4fd0d0c8a3573cda81f3b6a5e0b34b7550aa7afc19f8e20ece6d7afc87017234c2dd740063920ecd68b5eb21c0808453cdb391e7232c429fefbbd447b2e8bc26133c9ab05e3abc5bcee1ddd76e6caa1efe2f9aff4edbdd84e77c1e3bffa3a1ec70fa03547362faec8bc3d4ea322f3505909eedfac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hde0663f12d62220842503a7a0ef211abff9f187c2c4fe90b9f069af90f2ec4af86bafd3714397d9358403197bbefbf398c98dba23b7e116d1f52407e46c4653762b71761e769661662a26ff2dcd410d33e50202c78347a4f2c89ff76e3151690fa3a8df0b2f35e4a84e7e74a12df18af268574c4e53204264343e0f9e706f80e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf3e11ff6521e97448c172e1a6dc02beafbb6fa07b006130476f1655d640992406270d494a1c99c43d86d4e1b404257f7f51dbe9141c3444e2ddf5b5c3f411f59e69bb937677ae7705254c7d5d14b0731f15f7e5918dab021ca07c5a4db504ed8cb869ede0e280376c19306cced8cdb5d87bc9484a32f278ef077a7c49cbb5c17;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd196174080681fed79e20d4fbd9cbc8e8830b9ecdb228a2f2467832f501e3ea785751282070ef6cbcb5a6c28671d76c654f5985d718dd570387ba8a49fb839e2028accaecda6fcdb8af88dc5f2049c70f68407c64d40d228a95dfbef8318ce0da392c99d326c3ec60b13a0609a5a4ca519963ed7defa39c7dafa96c998063e3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94bbf8f7ca27e21f6d9df7af2b5568f1c12923dc39fc4493a9d111545a2580388c2d4f3d61018bf7f8406c9c5c10ce7ba8ce79aff1f044216a6ae2629f0951fedd16f0c24b8cfd504904523665ae3e4486a6265d61c0149dbe536d98d2242cd45edb683aa68ed60b7a2b223f748e1733a48583d3cf26b5030895e1fc52c0ad6e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha786b6672cc2e0e1900411e6508f426fc0565bd36165062215772b54cd262518266a95927e6a67e4d8b568809bb2dea0aa1b13bde1775fcba5b38eae8abf19b9c65c4661cff143ef54b5bbdaa36cc4a5b28bbd229bc5ca864696c0393380f96cbb948e06fd9a4c764fe957eaf893f206b2a3761cd966e61ece38d62bed577a2b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hba5fa7b9513156c3820395842452dddf7188ea64edbaee4a0312101adff70e2544258d947816967eddf5af6ac9b9c5c75d08e146f08d1cb36eaa0eeccbd4644dd1928a84c7e1800fa5226d980a7d3e442b9f32c93e66d0d3d4b28012030228af07d197fbc482226dfc4bd825a55cbd7817f67a4ae8c7ee4c188f44b81f41930;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8ae972f87b5c23fc35108299bd13c64e0ea00f99f517a77141425e17a90c03e96c1a5f08b2271300eac374cf624019b3855489ad7dd8283dc21adf06cdec79375fe8840112192213106aecc62a42138d69549f9ed660c0fe3b448253ac3de3755e71eaafa96065e15fb2e2bc4454e2ec6575852800b9b1fe0b933f36cbfd9c16;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94aebb2e6f56ffc3d5795632a666f8e96bc90a60f49fa21a1bdb53d6ac4b5cb7218e0004635f4c6552862132d6d9edf1c07c6b7b2056b49dd1d93b39c7e7098a0ec7dacc6554bef1a18d4203713061510476212080b864261a0be2721e0f4ad5d53850b6e80ac367b578c4f60366ec311328b9f138cdaf9608fa17d0f8bc8da3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he22c61534d42624b7fd41d933f76b046eb07934332d2093fd14b87ad8c6ecabc7f668e7afd1f2075feb1709693a37b7c69057d4e976153e96c794d77a5e6628b3ea17effdf8073211357ec085f68a183cb729a357c1475a073194adf361598a8a636933cb174826bcdf1d5cb2e70837c94d190ee89553dfd580bad567445fa33;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h136d4928812f99ec909e4d4515834684289ebde9bd996ea0ffa0b216595857b374dac835ca4e0ccc6032d1355828c610b49396a609e5e2cf213849a421b4ff22a9426d19703001520e7d1741b8008323d73515d6ac2551d45cc60e3cb9f8b6de1427c7991518a80d6b60e431dcc542e40e775cefdad8903405763ff80d6aac38;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h865e295888c756c551dd10fa712c07dd5d2bd9fa875f8691dd575ea00bf608029bb3bbacf59349e3f67859bbee8bf706b0b0f5b9ca646b5ad1361c2858f3a0a76bc625cf6a29889f885b2beaa25582d21aace9f3d62771fb8895bf44920cd7a8e1ae307efe86be2d3bda4feec7936ea1fc6d65346b4aa3e9a3482ac0fca49f8f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb06f483aea2f4c7b65cf467f00755a26a27e13031790fdcda1fdf8038860913e9aea163eecbdd8754b9fb81f5289a4d242bd075f69ccb4300d087eaf87e53ec6ab3ee4407c5306ddd1e8dec009828ae3725c72c3f45279442a17ae5e8ce350e277a37586a78f4220662f673609997a0fff7bf2ed06af3f558e6053a598fc1146;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he15b61713a046378f0e503e7f2a336cb0ae633484d0fd00cc0d20e572c74291dcb0a03b4a35417372a690e9f2c6c1b0ab12a98f450632b2a9285bfd977995b22e3beae5ed51c1ef5ba902824de4a440cabecde904a2b15f4d164113daa90de111925f05509ae5fe6de5226ddf6670d7caa7d4d76b836ab96e918b7c08602c037;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h121384233f7bcba818214a42ed8428b129532eed8845b25576244f5c3b56835adac3575cd373f18dd3fd4c7b2e51e50f288ffc8393fc07ddb6817f3d6069916ac5da11dbc04243988398dc25a4a944a83ccdf9d80b0aa5a3e6794083f8682b2956e6792bf964fd1230558e89e3475866f08eb17d5b75a13af950ca8b5f2424b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h563fa55b811bcf66d182bbb61e4f8c73cb497d43cd525f43965dea675d53d6308c638c15e77e3ac623f23b28b9066709db71f7360213d84858ccdaf011137c407a80d2a33c8215cfd79c053c73f9f7f1927fe306690766cbbf359ee4c5b79a7ec0b183e7ab06f0f27904f3688fbaeb4fc81232297553dc4da72b5ce5262d2e80;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5d9ebe05462076492d158a7cc4d25a61a5434e4e7e55ad18071c6f0e0efa97abfcfe6c612f57e422ff5adac5a5111171ddf325330b320a8b2429c7c52c17a6cca4fe7e5fcdc374e1f18f043d54ffc3a15f14834aca94119564518b1659fbf508729fed955cf5ca30fb56d02e758c5a77e58547fd46ae1e78c103ba81d4c5f792;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a5ce91316162d490de04a2b14d2444ddcffd9dabdba49da2d1b7af32f94f9c49acbaec217bd377523ce6dff6d5db10386d77daa77385e4603522659f2c9da83e6a2bbba36da85991ea1761bafdbd736938940f8d9f97f2439d38acea43e1f436663d22d9c4ea276976f47f775272e1861c9ef55fec2f909e874711ccfe1c872;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h9f035f0470f688daed61b1ff9803d45dda65af12cdd39177e7177e75914527ac5f8a231a8411530d82e41227f7631a6aa6d3a550a28bfdfbc916201a524cbaf3edec274d3e92337fdcf9c39a3c4a716fd81a135779383fa604efa98c7cfcf870fe26076ef7a5be4b55ef5da9251b7615eed4e4babcbbeba93b0bf4925c643e82;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha86a4e5ce049664d338b90946a7b8b02a433b1f203fa0364cbefc58c7d6382d47bee96d48766d4fe2974bbbc1841f1e1fbf5ea442633f8f06c829aa6980396a8a1387b75b58fbeb1f4cdea97be2ddb1b8160473080cdc819c5383f1dfac8e3f2c134dce5416d959e44b4ed68ace5eb45e9f3f50699f78950d16b37116f4572f0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h18aa5e745510b7d05cbfc2501c7d3ae13beb672e5c326df1da9c9172ad393ea3dce0745a2e5039744b4f4311295a3d2d5f07a6f3559782d215978915843d4f63242a77a42f33faec9972b22eb8fbff190a713340a6597d1dd284c986c44f5c1b2ab84c9e17d3afcffe147d9253a3efc931f6bf3617ecb0f6175000af27e1bedd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha4c7a5960922e47100e8ef1302df388c2099dad54186c481125bee5293e5eedf74710e77b995d62da46cc32dc900d04d7ee25028e50223ee324cde7c86835a015d52692ae2691f874b06e783d49eb1949c18ca9d90c00dc536bfdfac5d09242c27577d93086098dbc55c95c71b1d3284055a2ced863e5e2c3349f6386f5d635f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bd4680daadacf6e2011d5cd077119f7a8e4a036dca68fd27b11cb4cfecfda36dcfbcc1e3e24a010e06b8d23b94bab417eb9c578110d31d7b1276bc33f2ea058bf5027e9cfb8f46a58c9e36e220ccb434825c18ca2fd15b73727d323c49d728f59d96356f60fab8a1de1f9e507bbe6a9ec8059fb84e53f93f1a2b72ac1bf3c5c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfa2bdf47a814bfe89c750a86f13012328b303e2174ae4491f8ca295cb2cf1836c8fa22f47ad1ce8f62c884725b188f1698601677916eebd642fae88f985cc145420ffe9546fd7d561247cb9ccd48ec4bf8302d0ffb2e5cb020745d4a0363cc987b159d5fd797de822638e7675198b9d2e191526c8997ce1616c53942cb5f0a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hefcda81a7a003147819ef8df0a11d635f57481ff114c817a51332db6f3e113bbbb17742c55b7f0abb6c82b35f881f10a198a5116714d97b3094425ce59e864d545b4de06dfc5018ee199ca870b27d30a1ef370d6dc7a073477c752292680290f6f385f27651bdf23cb549eb1a9fe7e2598d8e0283dd68cb66bc715bf58f87f9a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfebea4ce1b2475508b0ca849ed4c5054b13ccfe8c8c2b7bb0eafd259cde69b9068762364011f2b8076edb4c2f38d7db1f7f387f3ff643826665540c9902633031f604e47f36b70a1689d85ddfb337fa9082a2de58d7f95ddc2e1eb293c165036c8cb853aaf2758d5c9b46395581269450bd5e7f31d4f435c8cef22695df99527;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc1c397fc3c43322358a5c47d054b8efe4afe2d2b4199ef6b273e430617cc6a206aa3968e8895a03ffc7bfe6aaab687cc4eb39199f659fcd28dd2012cd069088461c299709437d5eff1605b95861e56e4b45337fea66fcbfba4ee1c163e5ad4cc72642923ee94c1b88b3e9dab0fa076ab6e442eab9d578fcf775a247cfb3c602c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8b8692500f18d9cc289b3bd45d84af06369c1ba41401f0633aff48a64a7f60bf3b44617376d369fe6617d2e6d3fe95e16890d068e6885e683fe29a4e20c8b63911969451ab12669ef49c8ddded2a63707dd15570c25ba30958e85a929b06b093be24b3c73a4c05ac8a51209e6409445699ac4199d93a394ac13a24167d59ab7e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8e25294b422b399ceb2f2d25bba4bf80582c378ebbf0c2d38adbe41608961151ac3c87de8a673c85e305552b594b58f5dfc11e6fc7f21a6f1e45ad3c14d59773a9552449f2d13bcfbc999b52808ef95a5c729d29c8911c4c067a2099aa4ec766e1c6b2dcf3d34fb5d899e480bd9d5e67acc08674ec5a3d44bae2b189b2b57adc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb6500a2c4350ea409808e893b9359518840d7537d277cdf84db50d29b26220f50b5c48af70d075f4a7922a0559f6b8f833718b4e6a060e7f82b9d002bd05a6e6286140070605126fcea584550a54902b3dcd5e9536acd474d42ba0806b81f64e2eab7c90c6dbd34489b8697763f3b1adfe07f4154930a8194e31709cc69a28b5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d54175103e14dc7f90507fcd2e760b3ad4c1c0020a6b168301a5331cab4a07a0d3ffbcb6bd7250bf2f3fb507e89517c1a3a7f6205e5d20f28d8b82ecb58b934a9cd549dd52ed2ceeb9ef1efa0d8a208fc56e2b047e42082d4c1c2350af44a0bd598f11e17e69d30684bca1662d826f6352560891b9ccc676b6644404162b7cb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h665eb272f21fa12fdd77034fa13a20119bf7ba8d4107267a32621f94470f1cdbcc061ae693923e22aa960491126c95de1f6b657bf4d5425bd4d0cbf26ab111f3835fe39a689d09ea5c7a6e2f9eaca52ca61a4515ef1a2101b3ec37e22266c52b4e3beed076195b75c09d201c567a208f81243bd122966a49fd0b30a1880c929b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h549a7d3cb457e95eee71085988c68b0d5350460f4ddb95889c7100570cb9b0ec77a96e3f29a4f472bc0a6c1152347f463f786e452ae6845dbd923df993142ef2b58a4baef0741a59969147c2c540624c1105ddf5d5e364f49dc91360ca89077f20c9c988e9620135cfe71b0a804488da4a14c1aa802c99af4e879e37f088f694;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc5c19520fd52c5a27624472630ecca465a9db8869b59e898f9859749a80a812a56d4f4577a1d5e65c1e6c71737a26b73bd8c975973f0072a029e252c06b17b2d262ffd3b330c97212cd833f09ee26a595d31b122e86dee2d8d5d0cb404c52eff499e03b334e7e09ba0bdbb60cb044a6b4792b4c3ee0279549b8dd09a75de7ad7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb08503a01eff3699987e26e6a860b0e10db43bf49be6b89c71eb40aa3e56d0dadd76d75d1a3ec242bca9a66d58006992f94912825bc6881b8b156b2dbea0eea7d7efca124d06b34b8bcad35d8b960ffc564e97721cdf177dd6a8965259d149d1608db3b4dd5998839ed40dacc5a311c5e54c66dc860755f6782de2b622fddb51;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfbdfaea4704bc956c65d21e8b42a1fb8711b94bce6293de3d18aa4fdb5fadcb69770e22f81706b82c6aa237d9ca8db73d3b586b71d074af60c0433d346a3cd1a473e5a85994b653290c531583836330e51ad46df9202e0f58106a60312efd6f9caf37b47b23159e46e6125f364ed64a44390b306c3ece6032fb19e8429d6d9e1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2da95c38cb842ea8df6cf2cac5df45bad80b0477cdc350edd41281720a623c0b6f92b044e1e0487a7b2ae50d54ffe9661164dcc16d4ff9c6e5a4a0c0a384fd19c43d6a045104c87fb5ebbd696c085e31a3e75c31e8878b2fd884314e8b56ac8f2bdd344335aa2053191de3081be698032ffd75aadee87f80db84075db5d6a6ba;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h20b0b4bcca158e487797a2827b6ba6c8b78104e8d5999df844ee5116f7bdeca9997e99d07fb08e8d6fa7f95fd7149a7bc1d1abefe0ca266e3668370af1fba9772add27d1783bd8dd89131872b46eea2e9e9e1bbac7bd03ac4f276b75a4d2ae407089f65d95ecf6d0cf2196317724710594142d44af555b7ada2f10a759bdf653;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26d9cdde412ab743dd16ce42f59c45265d8a98d872395bd6bd95a32d78b6aa52ba677a67d906872a74ed214f916b173f51ed4ece1f95aea287314f1e6cf8567681788f987e5f49f0e5b290980304d6d259a14a79e490e8ade42c0c9a87f51196b4d71b8d78a7e4d470ee4b82c7adf1123bba58b29f7d2f81e5b63cee569a6b90;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f8f097f12e4c9a3480a4f90440370ed5e2d32673926539e10dadd459f1e5d7af5dbf888a2af0377cddb2b3d48f5042eae344636e8eed09de96c9928c58b517d508b3292c548b8d716d784bce94bf7f4ef9a6dd237e0b90c347c9e0cd95524bbfd06ebcb6561d3c8ad3e861b9955ce861fff715e2e0d09d0a61e130da0a3bcea;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e73be729f236e1d445e866f77c0764ac4383a1fdfb2497750fba59abf4586cfdcd1bfee7d17732946f8857b2ec664b072cfcf0b8ec03d738a29c45e8ce710cabe9b2c1403fe6aed7d576cb487ec9a163ed64b60a73efdb144d083aa337e6bfb09cc668a7ace6dbe28c3488edb0e278a94ff1682b88c6fd682bea47992e5e7dc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda180a578d43a63fb31fd851d0c97c8116538a1c03123fed77ba432273212287c7aa5638726bf9ccca507df390d2d7f22ff3c24e1a308c264503147c17c9693a9427160d59b067f058d0393388c66f5387470a5029efde6b8b8e80043b4999ed25524f38fae08a483560ec4ff920bd825dcadecb35318ac204c68fb54eddcaf4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc09aff022f9edfb8bf08526201fd9c5848c42080f4fadd892657fbcb44602f1d79486e1f7e8b5b5b4ff066ff70bca3112c25d5516322307b5540d0d42e4265e6aaad8ed47e899f1a9528023f86c32d07343efd6875cc60a42bda1baf80232925f1e0c0a3be8246e89ac5cf23ae08cff99e546b8321085b7ab775500b91cbfef2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h91a3d0aecb7a210a2c3679a5cab1bc03c1d40988c11d68ef88fc8e7352502b077b51c468bef984cefda5afc7dd2e852b2df1c6f3ec565d71f746d2e4dcd016aa0703e9af46f6563956c3e4c6f37e3489708739802694b5517b5f67745988a574c263ac1bbc3ca92992b0788e04db20f618e37a11ff4fbe5bab86ea9b75b5e16b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he03e6d68a1878eac75630cd1f9583d185b61d346bbb0c35e976f387a680ef8b690dd6c8a358815034990ad0e0baf43f53e6bce1148eada33dbc11295921e2aa6c675bb793cb2d1f40766e867d8517e029009b73569709d15b40f342c2d3718d66500692f319dbc700a81859d63a591f92d65abda2e0612cfe4610521912fcae;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43f0119f6054f821a020b146e5a83790ea0a64141f41bcd44b9bf4a58b17b63114cd31f302117173193f6db300458546e1ef5505d9f445df7540a15929bab5687c64714f16d4e60fa90c10df5a5bec69440c42976cd46de8cbc5c98782861fa6720ce583b46269d1ba536ce63ac35ad1c0d9325d148804bb6510d5f4da9b270;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdbc72513d6b37a5edf95fbbf92016300c75411b26550961f608f6509b34a3c54007b6644f520edda5652347e0b8f3b7f21b56c7e2dc5efeb418a6f732a1c4b8fa96be8ea52e65890fbb6356a2ada597f4609fcbdeacd88d164862fafc2095b28a19f01f1480c7c6c0417de98668f7cfa3d6dadc1cd5e586dbfe75c1324a4bed9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd129bf3b581a59777414396fc0393e3a889a35c66c0cb8f4b4403dd84ba922a3a19506fcbf07756c5563f665dd703109feb32a9981cb6462c89b7907d44f788040499ca8aeef18f63aece46e76863ed0ad5268d4c7e0d76bbbcc0be482c3b46475d0bf667a548381afa7b88195a31ccc64f090bd4b261cee786394578b46ff27;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6c3861da2635e89c44f27a2343a51919ec423e3ed58b51886fbe74adcbc9f4bafb38b9f30d91888bccafa8ead80118c72dc0e93219cc4aff0c2e80d032359a62ba28cf07de8bb0af1961afa581d0a9b20c5d7cab6ce7e03160a6b02b43d31569e5c9adfe0bf8a75cad9c21a6f165d824915b15cd733e485c47567fac03b8eb2c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1e53a9c6e1d1044f6deac98c41804efb848afe554f55daa1b2df2ba1554025265b8cc187e8ef465f77c7adf3a37aeb7628ea4f56d77e5ca2416761dc4eac4f9db2b69f6ac2dd0e583050f44a71cac0afe25486f28a0fd83f113458ee9b1cdb59bf491b6b9f1947ea18ba312a90f9fd91408728ce04224f3cef701eb09cf3ee56;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h62f9373cd1d9ee8ed03ad4847a00b1b7fe484f38afafee3c00b27296282336a61d43d0e1b23327a999010f6e8c15f8471c3820f10bfee66e5cdbae4a36d6ccb6cf00089053239d0896326d6f86b146842df5bd71bc202550e8f26b5a3000a4ea5e33c0b6cf79be6695b57c96e4414012dd7effe0ab18063fe214eeed6f54b9c5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha65abdb9e25d8a71b21224eb56630f6de11b7f2a0e677b173572454a65aeddb969512da6787c8e95ad8dd5472dfb42fa5261fc08dcd94e7db7bbd9f02be5801d3d30cb1b2d9faf75cf4ae363e86c846e0f5dd1e1a1b487f8100888db8af0ee2e7038f1833b7e9e1d841276a99867f11adf57cb1441217c4ee9ab8054617912c5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a1747ca45b86dcdd53cd1edddee445271f2cdf1fd4d899779b4db67362ec027d54b94698648ed53437f083dc017d1afc2334e7e40acbbaddf016483065c6bab1f643cff3f42d645b5655d97d11070f8b3ff827e7ddf1ee0c1e37d44c78fae862d48f526eed04e1297d2bcc07c8a9fc5c92ed9042ea84828b2b83826d2fea24f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8be9e79af81ab29d2b749e83e08409cc4888c7714b33112686c541f7592d2e696aabfe651631033d64ad0abd414e79bcff5350647b22cdad5066728c2dfc35626b86cbe9df5440e8f82348ce565daf11b7f213988839e76e4c45cbb4d72848d9550ccdbe63d8bbc991636316776ccca86adc71a2425449618988a21f27de210f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3165b09a37ec55b0d8cc6ef1d2d1aa5878246f8b9bf3e095c7244081a829caa1904c4d2f2614c194cd22948d3179feac26bd2cacbb658f72c394dc2a5209773484d96a666e615f583b81baaf5e0747c59661b5e93cfeaa445de33efae380a2dc9e827378d5fd1b4cc13fdb6c1e209f27525935f2cba1a6a8c366a431b905c214;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9e9ceff3662f087ed327422fab19d2fe79fa9332330e67762ee05e376ee05b2776a851892b5d53c579f02489ec7795136795022d7c4901df04fcdba93af16d7faa5a2cdaefac4a2846283c9d39fa840ceaeafe060a5df3152210c68a86269d90004b0a2ea1f9f733aaca1de2a5d3c5d070c15759d2f8206bbfe02114683dded;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f2d0322a29369ac3c07d548c17dc35239cdc2b75f6d27f0eb8abd8a64003f9e41aacb53431e1a92e45ce7662e3501464b4b5c063e0f2b0dabfe17cb7f8734680f7ccacfdebf7934c39b0845b48ffce7f1a1f8354bb85ea61ea895b95d83dbcbd4f38761972d25e35555ff3b5abdca32844305e522f8783e2dc6f6df118016ed;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he786a14cd047ff6e0f6d689425d7ac06cff207ed7aad4949e15f8bed37332aa87873e2bc3f7eee1937cf4ee9847130fdd1d5a25e967abaaf6c7460febf36bfecca521ea4f38439494f252e94ceea6d23e9b7263dcf329fec8f84c46d8417376e2e91ae9fd4a0e4b05a6821b15a46b6d7393427fb5295b96d8c681b930e38c158;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h35c2b7b99fdc6d2a5f9bfed2142b298be928d92de5246f1d5be1671c99b4cf8df601242fce7b0131f65ec3e5e8c5fb259bc451219d791a4fddbd95e06a4d5820f3eda5237f72a92ea7c8833ce714540fefb1fcee1d6b71ae3ab7ac32e171f938e1beccd79b7a2b7a7cdd92f7c6d61ab676feb315c162a3c7fd38c6d41ec0e7b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c6afdabd83a9c44efb8efb1891aed95c05e84be614d01992ae5d77d4b3d74db035bef0a4e418a45b8beed0f386ac8dcf472afb72008896ded60d474b2858db9ceb2a2475a376529394ff7b1935a95d7f6dc47619c02144f933e193e492ba22453f7831ba13730b21fc5afbb5f5b9f2da97f95c1bc593b74374c269962bf4f7e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h239e8016458b8344f24a908e6147d677b251f131ceeecd064f8d7a85e04fdf047bad73ee95b91dab006b7d1d0771741ef035205e02f274148c4dd97bf7099b36d35d16646054e62bbce7555f4871744f4e4fa5a9a275ea0f1d0b235c073ba231edcfda394d1943207b5832740e9da5411ed3b7cccceece460c221d4bbc78d6cf;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbe98d2913e067a9f50393f835378205124de85f1673a851c43a9e23a8c491755486e3c742485112a4fe309f66dc3276bb1a77262b1090c79fc1d1c10e2afbffe75ba9028484ac802a02e765b35a3dcae36e7fdf0630fd91e8d147bbfa1163d5a6e0411a342ede090c657286159cbb545bbfb219cce245ad125d3528b0b430ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3c5743ffd002beae4cd17377f43ded0147bc25163575e01d91eb700ad06d13a7e64753445bec1bf8c10d953fa4753321c9f436202144e93559bbcf4ddd07622596ae918e9ae09f46f855308d6e0e2455f2ec613ee21be7833f86f65038171ab44a20ead2cd2ab0f3f2e6b7e29284f87ee200f0dc380ec92490ab6842e182f8ab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3f0d796bf5e913e6166dd3c7610e6a6d9153bc9515a14b8002d96c0ec05c26cd0964f1eb9f2ec6b46ecbaac255564b6234ab665434f9d343ae0addae6e22b2f4a2b51142bb85b0b1c77f12ee10c646c3cbf437c42b7908cc19bc45599f5cb1895df5df30b3e29e69d88030c5ab23875979534df164476b20e3ee904f9facf0e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc74d58a6bad9cff81c9b898f0fec30cb7d29d9ac2badaa2a9ab7ef2f0061b4a1b05473457380e70a7392c18d630cc32fb018718d99c79fe0508636236fd49b718538038eb8912220bf77d2f45dc8a50ad54e0fe5e73c1f5e5fcf901a1dfb2b6c4fc3b4afd97fc8a2cd3735251ad40f4e604e9859d8c4c95d1aa7c001cb64dfdd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h17fe18f83980307caf2f286a5a9da83e90d029aa61a3a81fc29846af61b8c8b4353c7404681906d0defe0acf2bad757e2c910811a7c097c631fd333da2a925a35cf4dbd370649f671f12227298a0b216b14a40fbcb17943c7c8eb78f6b2dfb73009d47a845b957f0ec211781725b31414b5fea856d2fbb5ec329ec964bb06ea9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h72f6182341754257a44e2977aa8953c0a2a7aae2fc217c0a824a8979efd1c8c5ea598367f3240afd00613ccc8921fd61417e03149ec86af91715a21ba885f5e40f65208c6c29b73247bd7a2224f95548bdd46af8b5f006e2987b16289e94a15163e0b1058a98d3de0212d83df167bdbf32523feb8315cdec6e930dae734850d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h26e740005d8c5d967688364abfc075e9fec645a343ea69f6dfd30b25721ca9873b2c5176e35cf9fc336e34eb36d271c097d50543584932a787b0ecbeaa3c82a228699c6172ee34d0f8c17115cfdb0be5b542927288c1141f27aabe723261ded979ce6af44b33261503834be10dcf84eba2f6a5e98c7e79db30b42f1a1e992cec;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h96c45ce2d7fbf1ef323fd502f7e9eeb2d7768f4a92d26d0f78005d5a54b63e3a23dfd6952915f8e81a38978dc844365da9d60e805efb972cf93ad5cde008c7679e90d13059602e51990a63d1d334c7223b2543a0a5d2c9511455fb89489f2e5926eafe8b138754c73b317b0c9afc78952db7214f4bdf8ddf0c84e8e9a896b9d7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbdee85aa827773b2e9a389c1d060a9e68b9d72c42f5905e481ca4f00f5b5c0bdeebaeb0a0e2c8dd69f4990290f60dff2c4c858273e5a569e212f5682426d1fcd505f58caecf5aa8ac162df9dfa644b403083ad6bcd09d7c5f03aa8168a40f0cbb2eae312150725c2bb1852e50f3b8e8dc651f50ed728c9cf86ca6e929375a902;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41ea494e42838853605b1327ba7e14b24ac0b67f5115d6a3f268b65879458153729719b35b627cf693acc7ab575a50ed61e4f62ff90b91dce98e2f274fd59e3f40109793d922973d0f9e9aaf5beb5db315fc361f1604ac2213473e2455ec71cd6e4a83bd22b79e1ddfd59032b9e0693b67ca027c3f7bba5098923a3894047c5a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2247a88e9130330a1ebb69ba1383935c44b6a70ca386199be9a7a9a019a22e2a86bfd6240179836af49f5920b90a37135223d1c1cbf25281d91bdaa4f403e31fd12b6a9532280c5e32cb8746f2a11826329b30d20f83d159c3db282e8cd1f0f1f131bba4fe5fd009b6a06ae3ff50018596c666fd1c47e8b44b9f2e88fcd2a1f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd43ef816b74309cb8ff8cddd43c56570f8946bc2c695b4e18341762ba0732bf5f29161cd19126e9b6db592a647ace2c31d31196aa26c028cd70cf2341c4ba1ad22b78adbe61861c7092ec46070f7ab541c1248ee80c36eb63f1ce404bfec0ab93682e190b59716aab6e3486e8942e8ab9b9cd34b981d320204cfcfcf396d5804;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd856a88703fa17f6c2324783adb1e8aa63fe90a33d5da599d1e73876ba8dac769f1433f8895a68452eac72a39ad18eb45325155ac4f2097bba1910a8facf3ea2453fe087c567a50567055ccabeb20b07dde7af97e44ab74567b2e9f67565905eb8ed5c823fd516ab4b53ce5a47b91e41069929996b27f5ec9835a29a4e25d2cd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2e8f62fe833dc3fca9db8ca8ab9ca3ba299a3889ad21838e141f5c6b5d862daee48c85886852f50fc2f6109656b5c06482435ed8cc2e72ae5c9309994971960e9331375753ff689662057753731a101160e148b7c8d0fe0bd88105b6d2c4ad35f6681f71e17456badb9f2daa0330baaa6d135191c69e6c1dc32ba12ee47ec9d3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h989d4a6b31fdf1a4064c3ffdf8534fbd32d86afc3e3d18942b0ed22f7af190ad3f76ba21f10157ba8a4861cd1e263a766c6ac98ae47a2a929e8e0b042098078ee71b8fcb9ba435ff6a8c431adb36b4281ba92228b8087396a7c56561b9775c8c128c4e27e4207e345e4585fd18d9b850c08e19c71996cb93de936829c447c96c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h43db7d3d3b44bd7e186482f884f58cbed26c5c58f040b4cfe0cb3ec20d7b91bc354fc6b696b630dfd6e246c809b532fdd58e203fd24016a972e048027b5b09de78e4e9fab68f6ccf132c95ea52aa1bfa379b7d8ccc0806bfce139e8f7735dd517fff960cd57b7d024c1ec14483e2ca9883cfb0de0e63653fd2cc03ecf8f81f03;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd367d7bd704d90dd37131eddfd4b4d3fa64fa8af572b474ac504eba73dfe63d7abeb3e2a87a4944581aa1bfc4a4772e6e2320137077538cc4a0e2cee4bb427b21c473e28eb061f911aa020d1dd4fe625fb675947c5c7554b180a3f6569be8fff4f7462fd1ce1ae486e505168dbc62b8c1d7dd56fe4a7ef68a88ff80331cf941c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h52afa0772564993d2ccff669a9361f5661169d1225225794d71adcd3a58458e7a5d1783e7d26ea100e8c8f7b59559e37777161ee03781df9d3db579e154316fa93198c414ede7bddb4d99eec637e7281f5ac3d5560bda0ffb6d8a70cd00e56d310d0634fd139b3249cc560bfe02d21f764767e242546cf213c5d1894a19965ca;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h312d8eff0290272e9ce59dc0d91105f7c15d276ff5eaab38d82fd4ccb24cb797cccc504e3b80f2f3a25dcbc67b84365b6b4a1daaca0517532e63a879c54ffa5fe8099eba64bd2b4def774bf7e83a4cb229f92f474be855b5f33d5c399836cd992275a510b0d622e70108c93e98d4d618ef9329b3242ab6b1c3da37a2136a9783;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6fb401189205a38ba58d99b37aee02a3be8e0a6a5a5d13f07a37a3edb31054880fbfdb93461c83c2541bdf0b39d539519420f440000b75528f16573c4c23f242022b5e321a974debe0283da0522025b94861133ee52c03718b2986bc7057f30160f77bb55e8dadc71773dbdb5da2b7dfafec7d25fe98648e42da34980abc6379;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd9b435c772eac2691992dc7d53331f048f9d7f083b4d7571a9c77a897295257c445f92ea20bb917c075857bff8253c29828a24e8b28fd27e63da15ee6fe4ee0d21d426e87160b61e57b2d336d77b801873428b74ec8061cfe5352a7045c56f804b88e1ce02e07a68599011445c975b3db43a3da6dd348d34fbb3ad322db3c72b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he68bc444a2494b7d71dcc648cb0893daef24a38ca99422528d7e8f272765cfcccdf36e0c8f55d2fbfc001439b0333536518acbdc839e387b3e37a8d1c68f745aeaf3509f30bd39194e6084e290dc679122c366ae2a650c74a79d453e5346cf93521d95c3babc97a40f55da06a23b86e12388cae40ade0bac25e8ebd641d761b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3e63da3b6480e491aed29a2d6746db0d0183b54767da07cb5b55b8f4f01dcd6bc48d059785d58e0c01bbfe5028ee79377e0720a9af67c400a367d516b72560c29cdf6633d96329476fae960700ef02feb56198458ac622adaa6bdc77a88a2a156861243c32ac301e7e565d62c25114988ac4d3663712227a3ec90ceb31a750fd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h40d80a56b4096f234bac0242cdc8a85fd05797ed3c94365565368bd0a825be363ea57edef054f712308f64421274c0937cc57b57e1daed000808412d5eff2c55259bb5ef91d8f5e35cac69cd28474984d22c1c930353916b1869d554d713f3d43001261dce2246e78d418bb5792ec5f112e9ea90a0a2f95649841ce41f8628ce;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha463a8a87c44fb59012a977aa16af2034fe13333d5f0d62216c1014385a606517a0fde10c3124d61381f6e03f259cb999665dcbe7ae6983be2d8a46236baa8468fdef99fa6035a1ea6d3dd3427dbc2ef9b693119c0f89d7abf0d297876debb8e0c0db807cff8f376af38cf9ade6fd43abf0595168489756edfeec3e46bb71d69;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc9edda30fb8e305f049e71e7d48c1d674750c3ea229608fd9c964e36fbb30d6b528135dd7b60dfce39c027191f4d79714a84855b11f2c78b054e527fc27404e02992ba85331a011c84d05b66bd0500529cb32e2a52312b9d25cd39c01a7187c0bb1c685517b8c2869a81e83241489da0edf14e4eaf2c3b3938d85a5b9f7d96d7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h814a41dd1931938c2e33e57243a8611759d32058cb82647e097e5f2e49e457cf71c4040462657a14633baa010f8879bb66d424154f8eafda17a39c9b0acf622603cd5ff98398602c99442fad643c96a9d392688fe98d40b5a1391f05e82f81eb070d2c33276e8e8e3d7d10e0aeaf007d0d0e5b3d1a24d5b6cc7f8bdf065a6a51;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h34e61a13ee7bb6f8298f18a0aed4cd38341e44e568d13ca75348a7837d1e67592b420d7d23a80909b21d682dfa372f4eb3fe79dd7982efc8c946afbd8c38379752859977cc5c4e6646c0cbd5b405a775ea90618a6406f63530f6aa95ed3ef0d9a8f2f756b4f696a5242e86dcfa0bdd8492735cf0765d8bd350cd730c4be48df1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d1aaf04590105f2c3b07df3df3c52a635c42e0232aee88606d8d0239f2c69fffa6a8fb7a41e9e9f4af86080c120a8f5fece023ab4fabcf0808dcdaaf2c8c0610c7bed8d0d3be518832e3f1d1feb989630149b99e4ce6917d9582d6c6f609b5a7dc4c9b589eee1a3980dadfff187eabb8c389e9526209a47cd65774bf96db4b7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf340d84159d52cb4f113abe2448a281d05c5d83aab8c14d3c88293c8abeadcb9d234f4b6b8511810f3694b2f659e13adc093b3e4296303e3c06945be1f8269c83daebcd6991477dc6131520611f4fe0432af44dd92e6ab679f698cf08f57a7f9195e7c6399352fd2c09249c660880a7f1bc51b799bc44c5496c53a270c5bafe2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2458c889414f7fc2574c2979a92972c03309480155267204fe6791880b93d2b1e20e5aec058f194e75ef4a7174aac27d5ef0f35817bad56040b1b46e2925fa9da34de9504c777b3767e7a311a55b2c9b4e654aade80468f1d9287dd65e407d18f387377805bf68ff7cf4d63de0422ca384de4bf71802d7f359f5e9a3e87b8424;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3295b547054c3a2a861d88ed0211ad3529d85e211d25725c9cf91eb285a7fcc93572bd9c3bc50eb112d9f9d9c9481c30e0bc50a57e4c93e5716426446057efa78409a45db1b5d0fd842530a9068332277257be7adac17fc99a5ade60f269b8eac58b1ab65695cb4a4fd512d1aead09cfe1e14e7c7d79041710498110c202ca37;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h902ccafd23bf32b08a48cd559deed6696068884330b9bc366e999cf36674eb9c49bf26efb84c215b4651e8f9ad899536622ded9eb6ec4806e40b0474fe773b0a3ffc5882ebfae218f0f8277c45c3fb55d6a1f0e6fd47953be00320110d02c167f526d4e80182a02bdc91e6e9ea67cc2eaed5677d04da86eb9fda1008efed360a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8f561fb56298d19cd3c9f708b5ca4b2a47e2f362cd1bc97304bfe59c4c7b18d60af101abf225dea046696b8434c97768c4a09f4b71325a44f75a22f4063d00c7506e04cb3ad272f820623c1ac3d955e3ee2014358eeba685a171b518b662ef82a05d4611ba20bbc3bd36485f1a7d9efb1f0c203cff48c4a69861741e363ab71b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4cabffed0b48fa46b8d75f41ae92669e458de3cbed3767c2276446ebffdbb756b547ac1647af89f5d6e2f95aec44a6e606aa365ea819555ae09a4bee71de800f2cf270991c51b6062762fa2b7716e93882b8fa6415478630388b431b2eb139e7615c3478a582dc3b2ab6a4ce919b1aaf1ec316eed3874cc02224c5f2fe109dcd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2490875620a747c0c2fea2130d3f9cd9e216bc8c4bb6c0e0cb764a09a59d7c922550ee04cad6de6fd372ffe03d379900a94d373431c33876d5d0dfdb740a5f747fc14c54a730bacfba6296801d60787300d104d0d674688dcc6976185d19e8543ced8da724a5c0e105d0c5aa57bcb48567b0cdf062533c833485d7f0c33b4d18;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he3faa16f7149c25ff319d3421b8c0c0c86f3bb3f2bcfc05ab4f94a5c6a74bba7b0e7ffdc10dd062110625bf5b3714858feaf8a02b7d71d813b09ccda4d333088cdb234635a3d834dde364c9d3e231f7f7c915e0788cb284012667f8691f6cb8f269aed91cc2c3c8f09644d00b0d1afbd5de905eb3f95c0d16942ff03eba78345;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4e0d864da853da6442e6d17fb113800595a0d8036138ca84c1af9c36bc40b241dfc7748ff2f0741f93e13b8338eb5e99078db813e2f550e1428f65fc031fdfa8e723ec0862a28e863a3bc899c6f98ab8acb310b9bd2aec352454d34f83ca274613b5ce6d55416df999962a8ce2334a208729df65d766fb3624b06486a0fef9c6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h4c6733610f4f69757b9e829d8072d377407154d08128a17b9eecdda8ac3ac3622e0f299a0290e95ce8ead859f2b5def304b46be5bb5580d0599c8768a39666da8f538f387003c07ca5c720cccb8ccadd410f8b72247090403b488fee51f4ec675d1e9339bb189bbd2530a7c04798e07b8191157473c54ea4f6db0befdbe3586e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2f5fed95246b33f8f0b74806c668ea433744184e382deb2a775d8cafa45a9db6de15a559df3d97d328b8b9d5c23f0ec285e37bc04a61556bc177a028b79c2038408ae672c502aff5fe5bb542ef44d89c1e4b6a7401139548e51f6d20c87ae448cbaf779675d57e6cb0f4b97d83025529576d0b8c61e1d67962184f4adec57824;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hffa861e6b2d32d4e47cb2b7bae95b9e19e334082b548a96c6f1f4a00ab6fc2419bbc42ad790912942a3f6221c4c950abd70b82b3ec01fc69e97a3fddd52693199963145438b610111dde85a5fd8d23cd5a0eea420ab4738ca3497de336e748d87afd4d5776c6d4b69f29b6a1db25d90bd1cb681199f121131bdb8106df38eb45;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfff41b221bdcbf29d42e264668ffe1b131104ac5569703d7df969074a9ddbf488d7964e5a4a09f5d2230622b65b513aa9b8e99a1896fc3298d9434545f3b5d2cb18e2704b8ee72319104911e20795483a795249105fa65a224761ef6e39e9b83e18a3bbf3ff9cb1237d5968d6c41cbee23daf389eed33d391ac54dcec31478b0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h183f5e62ce9921cf15d841511558a63f5376064fef73dd79feff933699726a639228645b8edfd848a908bb486cdaca434955812f1c37f233a2ce4168aed8dad3c9c3eb0b67d9881432e6011bc2d72cb6e491e15ab8d0bb083e3df642f292a3a4c811f4d0d16314f4518b5f827b639a6eca745c7d62aa76f5f299fddba16883aa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5a732762f0b2d8ce9bd86dd2419b2179c44d6a12a132cb5094352c6d41017bf60e67bb341a61885aa1068a5017f341509f4ffe1cfbdd672046665ec241dccc52370548d15635e9dddad7c412cff29622107f4ef429d691fe5f4a4ed0e9df294ef84a958d0cc0ea202ad30592155b6a5eb9f6186e282a18eb10e0318603efb0e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6dd016be0706c6a2dcb05d0e217c492cb4f6c798e6c8eeecd6478c17a6174dbf981cd3d83129fa05bfe7009e2f6e0c6b1cdef6a923e0cea503c5b5a4ff3518e1cdf29ce4d5a7307748af4097fcd2de26e21835fcba3d5b1a07ff28d9f21bc852689814e5249c2a0aee0e26bb43da2f7c5e37a8258289c93a832bc1c7d71012ee;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h985ee5937e4705bb7e38f57d2f749a0853781f8d1c740bdf1b090dc17632095f8a798043b3deb06e52811cc97c4a171aed7d2f9630f64b21ded87a708db2168171cd60371fd02f36e8d08d8b6fcbd11726049cd32f0e956d79fc46a91bddb850f3b62f220bf68c04ffde1af4c73fbb2a470102fea122a8aa9e3021d818618c8c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd55cb56dd57767b23bdc958072f8995c1a3e4100ae99fa6bbb34b61bb04130b51ec0c991aa821df6f544d2680bd11fd94afe6431530a142e43e7e6b7f431cc36ca169f63ece0e329e437a2582451038c849205967168e357157bb4843f09839f2bd0d3fd0a6fb6e401abb46f557327134f6ea912152e3f4d7964057daf29782a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h142d02e67be3c4a269ba3db6b64bad778f5bbe30a44324a8cef05cee3052da26fb31a43f6ba5366b8005eefe75022e0aaebc5ec62a7c5e63863dec88df85266344eb0a775cf9b0eed3b14659ee4ed8a3598f0efd95538079a5bd9f19a0281e03a017f122b1144ed7199d6988b50682e50b3e72ae0b53021d8c4afac65020c463;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd22cefac254cbbe6d4f7b04b9c87711fd07eaeee5f944455748e70248eadb30b2a6192adc443c443248e8ea0ca039e2c2f7dc907529080c1e614781d5365f87eae0d3a2e0ff867e9e8f88bf6c9be0d5d8e6865e147f11f49df9449c4aded4548a63d1d058119a746e9e2ba797a59d8bc57d4598589995fabf1556f108be69592;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h83e4c2c324a26e0f3b8d46c97cc7c63786355def71c67cdd1dc35d1c552c8bc21010e7587783d8931732b05585bda4e7b8db3ed866022fed7ef0a6b2e04e834473bd2547bde50e721299b133728b864fefeeb3a31ee9139992b05a3415974bec1676313c008dece5ca18e1a8ab697a1835cbf33a220b56240a571d8116cf634b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc30c674552f8c05c69a5d3789d574ed0c0044b74a5e287ea509312576a9b47662cfebeb759c75d6a654a78a702af198a444efd938f71a76129b87880ea16066d3b500aeb24bd477eaf254acfdd0e815127b1e945c9ab3d2c6704f77d09ecaf34d390ab3f73a5667d64d36e36cbfa6453e88e32de2b706ea91bd0d7cd18abb304;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h98b986f76f598e85eeda57a3daa217ec5325c1c2abc50c8d95abaf1d0568c8b153ebaa1c44c48b305ab76e7750c9655fb0668cbe8557bee460f13f19612c6aebfd06904073a83166dd7c48c9f9f2b20f74f77a030554880001d188e7ac45632f1cdd115a020ba2c121f93874744e23a8e977b7d433e9b51ef959c0055c636d43;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h8632d5355f7b82685c6bf921725efaf9ac430e1e5a1b2de2568f911ddec01545c8c91def6a72eca3cf01aadc0b28d8ee8c3c08b1ae23aec0dc40321ede5c61cb9066c1e5691aa1968b7efce47c19c9d2766a09213503fba57d8d749cc55fde967d25cc8c2c0ac792642b5543c0e87a2bded21993226a3ddd7141ecc7e62d4479;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h251206bf7d525b0bee431809ce712e7342f746684444d70e75ebabb15d0f0428ede33e74b79f732458595e4937689b2ccea311e0dd81d1d408b5ed5c16b1a0ca41a1c0a8c5821fdcc5b67a4b997c8769354f8065393c06dbd4f0b6e679ac17c2c56b925e32c2d1f2f1789d9ade7def4637b82ceba5cc0283a97c3b83357af361;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd0f44417b67c11ab69c2e23ed9cf7fb0a9ae2a435d241c66abd83472e02bbe2b82cf8bd42863642bb7362d5738b1c11576ace96f9ce530a3da83e0822dee58e43159cf5d0722b4e1e0d4944ecb3e54869d85fdc5afe22b6b7a43d852d2731d5066c15353db60bddc846d548a53795180687024fa9199698dd4e31081e950e4e6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he1f26d2a6e87778547a4b3af462d5484efda6077f9fd7e9adb45e93827cb907c43aee1c833c18ca72c8b8c84345bd1a8c5c07448d1d77fc81afa6a899d0f0f5722ff725285435766d25c61bc0b87881b95400b0c0e9f381a1b058b2a60d2af72cd8b2cbce17a6e604f06b85131a332b9fb602843a3a444ebf9961a14e92b9a3b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfe1b1efbfca5fe14ab7f1d34b5e34402b31309ca22439cc07480c6dbf6055af8985f7a41e12b37e4136fdc8682620e8a66face9e7cf3ca9abdaf7e5a72eaec94419efbe2a99f5a36f053764b969cb677e378431401f0dcb911afde7123302e6dcd887617be9ff3e95680e799ac29c6d82849b6195317c717803135d4a94f432c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h41036cebf25c5500309024436c699226ae84c48181404e956b3e6249efdf87b63bab4e38fe94920a35da794278cc46f2b820bfab5dd96d4149b1aa051b7c2d36b49e5aeae4c734fcb3a92f768d5f56bcb9a4c2bdcd7a151f8e1f7effee550255414532e1da6b3563c0c6acad5f61cc3a8dd0a7f3ee9528eb624b434bdfa285e9;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'heb78093efb7d3d5fe00c85830a8e8db5a352c91ccb4e590323d618644a188ca947372ed4a1bc84b2c403de9f9b3a8b87151716650a9a204cba553361b6325e11bfe4aecc738fa4d53527adc589eb3356c6a340deccff0c5f90ee7d488f03157c8cc035948c6aaf586947781cfe968c2497f3edd7bb759cec8ecba53328cb39f1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1974ea4e5ca84f95f7acb19913df622be62249f7ae886761af776fb8f320c680500c5ceadc2d69e3b7e3bc03b4ac7bc0d09e529889b1d1c76fd7f45b2822fc2d90c0470f5da47a2b4f0b8cffe681989fabe3ed0a1e27e9cbce37bb3c8db0aa7cda3ab6de745f80501ddb6ebc59697a88e441c381cd024686e2ef74857ca4124c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf7dbbc6af60c5401df37926fe17d6eadcbe0f4abba6d058579aed965d71acdaf2f16df2e0bc689e8201a6d412414af030a28f46854607f7271c417ef9fe3fe231a2c72bf7b8f432be5ed354aa95a502c6f1c3e1b286c4a4874847ee1454323494f8b91a27d23b5dce1d991fa4cfe01d5ad961510dd09e98f97dd8d5988ee64d5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hf488507cda80f561b2835d0f0f1db10b72681c4092f2d5abc96ac8af2a0bc54bb7c1ca8c5fe1715537427c04179c7dacdc6ba0e4f25fc1faa118cf5d0b4123670fe34f57bcec2738da091b5a44ef1dfbcd193bb24b4e8138014dd8e6f67c8852ca944ca0677bfcc784c7c8ba7e7156cc72127ddf5d19245f6346a4fdec48ad53;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h94355bee3c1fc6158d931296fd84e522cb0bde75790a6d1836b36dc0a33f6adb9fcac35f3ac7d510005c8ff9327114aabd144ead962cfe3dd4ce5412181e15e90c8577cad3c1e21e6286141b1859b6ed5dd34f8172ca6c79812ee7d5f0071b7b3943e5ee718493b5075f9672e7d7d7636ff58c8b3062fd483648a305af77953;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbab2911dbad0d0eaab0d400bf1b595b163f69a7a66afed68219b7015ef0460fd42b7b3de83bbcae73abe0e9657dafe67c429efa8602166ae8cf35cb83978d0eb59ef8cf8d7c328a1ad7bbbb2b122050ad67772a5cfd7f0d05dc9f18ad545df8bd028c3ff7f4b079144b0a52fa7a729d92fdbd28ba65a0deb580c91adb0506bb8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hb2aa0c1542c599f1f135edbf0d85c44cc7cb0c99f5957b7d0e21e9eee77df7d711e709002ada044d280e4f9fd0e164a52069bd99266a1c722a38cc399f1a21e80974242a8ff9c1c719d639c8b022552ca81149808bc4924cca81324d7cf75f0902bb2cfb00cbf15bae66cea83370509c274dba7e21bda305b107f856f7cabc84;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h93c8dfea3d79a0bae5f23eb3b1b005cb626c16199fd9953c2998563acf0e0891a587c362c761e6ed7016fb3377c1e910186fa0c7657fb5ac5bad856c77c0599bf033abe3ef6b8325c1fa3311a3d544f6b5150b4c2324d76c48770e428e271835d7cc7e6d3b63be53014bff1299f3aa18a302eb9d9f75ca319ba4716512140ded;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hdca58d7e6aa43698e011005ad65787116e21766ad91808475e35c1f00ce6ca65300f71cb1498a5febf52dd776f5553d074b993c613b94719011f6b6a1ba04977f5d57dd14c2d7f5b83f0b0a521174a1424dbf4533176e857153b1fcb0cad17497c5ca4bf32127d32d10bdd00540b6dc4df2f644478e98b7e786554a6af83ae21;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h10a3ee0ba3410b3b7fc73d5028614d7582f1188dea6c30132422ec30e8f7158f79bd4c5ec40e262839a1ed69be31ccdddd1c7d49668764dcb01c6d4ac3fce8db629bf89b4da9dcd97a442a0b0f575a7bbcc2e9ecf7dc93ceae4919a0518855367f42c791aea9da67d4cbce9b0e2c3c90b1998fbb030072a94228b5a5e0e26fa8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1a3c510838326a4cedbc5149e2990c9163d8ca448a776b098503080919bf2ec2a98415f386c86f5dceb1610d981107c0a709a87fbf05d0e240536fd1aa8a17fb78f6020134426defa962a5f5e9ef65590840a85485b27e1d454d9523a256fd3d9b8428aa4ab0a390b91b4c3de8c72d1a52b22d9add100a8e9947d3e36cd247b4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hbed75030819f09accb17b1fb4f0bf8c7fd9e5497add842a7e9d6b94897e7e4ffec3df91551af6297d116aff8047616f0467bd6977d4ff2b3d456170a2fd2ca316c0784219cb98f052f08cfb8098602323e0e9f14215a0b637c55a865c8e49234337b8acf26003a5eec7fcbb78a97c10ba45e3df9e249b673190a2ea67195298f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha2d5769840173ca96917a38491638f7abebae33897f2f87ba24919df7b960e9738a5a070dfd3ac11412a0cfcbe676de906aab81aa04c40ac694b7bb209af982dd0d9da531ccbef70bc9a98a2e5d46fd2ec1dc65867b2c02fbc6dc020cba9b68847a348ae9d66a7115b779fa07242623919aff8935a834a8999a287a9850433a0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd991ba2d1bf7be7bc8d5758bbc627d33dbfa9b28d96b7c4494940c98ccc2a127876653c1801d644a395075fca534e979bd67933808a112922df829140afef7fbf62b15a7b6dff54d2ff757a357d2a0ce4ee014a720c61b3f38f47d020aa05cec4baf057e6f3fcf780b8c8f845b58f8ed5d9a57024e1a6e923efa6baa3f1cde64;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'ha22838d6e9e549660204010f791549b8a37cad2fe5516e55bc85b348275c7e32a6c8b0a5751db5402ae07c3b7a9131105585ae1fe7edee0003f48ba32e62f05d38be3d1d6d6ad464d316f3c0f8a26f276f5cba85449532edac934d6561cb285e7a50a09ea00567f691eaf876a70c27d9542a1edc3c019b027057d453135e6581;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h1af8dbff20cf043b161a043412e376b8a29791f1188045441dbb013484ce6bd8b333d2f61b5f85a728dd09f32ded7faa160dbfa94ad8b10e744a7fba560533e4e32d381340346b3e97130c502271ab43803272adf451ba9e362438854a4283ab0f36a98fa518a2a181b558610b97b64c7f72bf77bae874ccbac87192dcc05886;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h194c32c0e61b0e4137f79026fd310916a99efaf1e3e15a14c0a72d1902c929518fdadd7381a325d2036ffbf216eb6e60b06c49ba8d0760b0df480e953b9692eabd3947930edb34cc43ce4d83b8117acc08133689240aaad5944ed7ff50e7690080fb15f6ea56c75cb1a97760ba6f90da4b542aa6975136cf915311b330e88499;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h483c35a46f9ee07c678341be9fadf3e746887a15645f2e0f81d779a29bbfd69c125a4541759c8a4f48eb151cfd9cc7c366d727ebbe18e08ce00fa547a0a598591ed96b50f457ec5f8bf2faec8d086e30637e5a7da9b0d67b95ef29c3c9c004ab4247bb17bc738f830c85a01928070789ee6c212868cb2a13105ef37be6db5684;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h547a992453f1886450b7b0a9ea884ff97e43aa55dacff58eed5afb86a546f32012215bd617dfa60c64d8deec731412b20d4fa48a0588c3f5b8ae6b98cadc30f335c5577e78d8c4353567a7307e5ef02673f3a6e605a5182c72db389ff4edcb8926ed68a92bd0ea217b8f037af604931bebb1b87fc3d9e98d2e9b2961c8020309;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5bcecb74c2a373826f3e015048f4924df4f43bc9b8a316941012f029149437de8fa2e74018073b4f4f2676b443bd1dd6e972f0289ea477e4b8f3af57781ea7706e6ded20fdf328017f482be77a8a5fa7d846e4221a4f4f6a7d9ba299bddd8bd749a5aa255dc548fa9f7677d36be85cb3e7932439f1484d16d065fdb70ed06725;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcd6e9d2fcd53d78878fd4d921f348d25afce924e8d8db5503b85c030a371b27c3c11a6abedfe6466adb1909e2d632b4ce9bfba3198ea910c467b8ff1ab8a9a40a4902dbe3caecae516b06ae87500bcc9953a4d43e5e5cd9207acdc68042378839cf2e3824a9fbc36acb5f8edb73f964d3af2718fb70ced79d40aa1972d6d2483;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hab91a71274bf621c2a4c72aafdfac64bfa09e3d637820388a08b51b5a5bb495c164e0f2cbaa4ec087071d620283d3aefe778481ec9584d1bfb92377487b53558ff3052e8face3e67d9df80796b9575a6fcac16f6863fd7c6a99013fc0a34a6479b0d1a39656d17cc062476ea2e84c0cc7107658a75724e4159547aab58a57d2e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc259665c07f8fdbfb81451bcdadd3ec7d0e602f93b520c5b8df6366596fd37afed45341cd5e45d82f2e63df483714f00ae35c888bb7c144075c0a62ce2f4682cec75d0150775ae4f4676f28d93d6558c68d07fa005e5147b0452895aa71b114a987f67ce56463fe271ad1effe35c97bca66ddeb9a4bfd31a87d26491c1777d2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hda68e6eb920f1e4d1299c007ed18a20c87bd3d285c177dd11536e19927e1af91b7293a3e23a1254f0f8bedb538cbfa9d926087ba10bcaf0490fedc85c1cba6abc451aec281c88b838239cd7bd33123deef15b93850950c4e432c328fedba5237fef0886ce2750cdc5ce044c9671a45d9adc04f6ebd884bc89a2bc33b72c53b67;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a6665190d830d4f3a595029f24ae41514cbad121e8e4e1c2d88710683d584e88b8cb540d8ee67c3468dc6f60f5a2f5019abec6fe9f56da7669f2241d174f7b9907ccfd0bcdba96bf4dd09d458f48f47a3a094c9cf2bede969714be4f0f6e6241ad314094ce7ca6afc389e52d4e56bb4e46b806e0024070ecdf9136a3aa0c7f2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd10ce25549bff5a5d76db19e68937d2b6dc4f5436f76e87c5037e077161ac5a3204e8a801c8ef68fe92ebd24ae074f146a056beb1fb90540b54b277a2588cfeecae8b0add52bb49c2cbb01635efbc0b73537523d9bcc8ef2f67841de0161d46f92005cc9ad4e5f2f6845ab93bf7d1985700d26d494d5cb15ae49190ad59d1de5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hcb868cb14f8b6966019b27f0a8cc1c903065711593c1490d8827214b110bb70c356572bf7d4035a4e9493b7f4f473ad6516d7d8313ed141eab1b02d77b5c2307d73b1437c49262810d38aab0013cf5b23eda2723704246bd7c3b5b60a51325be02fa85cc60a550c482ab31a459df928fa96a250a6d2ff7122b548d94dcdd30c5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h12e5d05ce12ef6fbe6d71f7d4947461592cc6285775ba8c6dc79d50a022e7613579c5031115b824858c9787401b5ac6e0c3077b13116f5f0a4f3a39ded311f88fce1e121626f9a6e5bfaa7449d855c139b0c3f80f2f02e1c54aed19d062221e6630caa18a0ffda5db53e54a1f7569e8afec0e9aee3dc18c490356b225996e721;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h137dd025ce2221c6ae76f752124eecabe3cc0317395f3c4e684f9b83c5c0fd16e8cf12abc5ecec4c84e4131508d89337f59a69683ccdd8889455ddca0aa998deae3cad5057e6b3472041f8557861a249a99173eb86e345e7836cd41b1f07233a5c56d74c06435a780911e88c8c0ea4d962e55273fde84ff28c12b546b5c3c311;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h37314fff085da2a04bae763c5b9e04da021e8be37481cbaa0718a98132ff7ef33119bdd3aa234a99692207b781459788f866898fbf4f01e065a0e8658c0682fcf0c415bcc35569b2b6cd9fe296b5774ca4c9ec5eef84fd7c827ea562d07c8c7d8b4aa9fe592a55eab4f2706db2a99f17c99fe4bd491626c2368ec3ce02abba71;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3027307f7f5a2f0723ff09758a79c9b152b521b0def20696750c65f74ad55116f7f4cb36954ce03287a90fe6a54f097f805498d00f520a588da5e351be8f39dec51f89a76f6c288a193453b2158403eef3428e917b4a0007c7433d0ed94594b386bf440323e22b39c98cd98f57cc18331a663564f18d5553c8c68ca8f4b9106e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h255bfc443c276cd2e0eae302f35f4741093fb2b2be34fe2bad1e03c7dd3b42786178ecf5da6f81a08d04e8446f2eb38a037c440e6e031ad0960df1fc4ebda8344aabb7c726d06ec35d2e6faacdb48bb58215b349eda1aa332a78dea6ecb6f941c0aa4027b2b9432e5bdcb74358fb1a1901682f23469ff0eb26b50fb742ae052;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc32706d1c5b1ca2879602e618dce484d75beed558d2b5c4b3ae543d81f44135dff9061af9910ee48d90b0e320f354150cc9131f0a28f9cf382685471e55f79ee9f3391dd73b7f545b72ce59b84aeb563e968a63321b1563ba748ccc2d517187d04ad3260bf000b0f99a68ec63f138479a350ba9e10e0cf0e779db8d1f06f0e8e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd6d0c5103046fd82f9ae258eaaa3fffa96faa402acd987798a8a242c5c48c02cd806a6f89e4b844cfa5afa5a1dac5ea17855747e0c7ae34bda2dcc64204ceadcb07d760fac5241611c8c28b5a17cce65d27734f01b7c921c36fdaad4f01af3e05b75184d3639b2cda8d7e50b7f9c4a74b140043cf696f032aab8f11279491628;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hd8633e1ac8704f99ad94f31f202ac07dc03f4643ca7ec520132f309e1af190e7e8dd1eb4a7df2a4dd84768c460e86b80e92084dd7ea2444ce62fb6fe53ec7494f8665373415dda894af4f13b0b05b124bebc64cb256dfc2419e8e06e1204128aa75c8ed0237721f41e58f0008b31a9625d033d3360b43dad0a41a5d53081bca1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h39d30aded4142eab2e78df6073ca59cb4d1f9e7567ae5b5aa9485ce5e73f0e23fe61dcd88a1f212d8221d8015f75c2e081a6271e0d459458aa2db3bf22189944028556744129f79707346599b3c6f18f8565ac0c90664c76a8e300de2c28f4a9c26562fe87e9fa1de8af6254fa28ef816cf8ed423dd85e70162efa5d850c37ab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h782da7a7bf9d26563a28be5383893a3122376aed5d4d40f03034d6246db7b93f5094aef5a587d60a0d64dc1b1b8cf91ba6a65451c93cf019cf21c953361669c6c156fed983a3a9edad46da2e74a157f46ed3c287145de507abb09c4f897a791fc2e770ee04a9eb88c5d7d447574c78071bc91a51992aa8e5377505835e5997e4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'he4e4e3a996593f9f443d154f3f567accc6be280d6c934839a5786a9c9f6aeb1900e950579be959aa0caee932c09b218d89f58a6577d7de9f320617b568b76f5cdeba2df3fb9e219e366fd700ca2b99f79d2ee7e656c497b8e028bd9983adbfc7671e2bcf4b30ae2d85c33824f34274ff4b40b2450b488210dad5b01c354822df;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h2d996643ae513b89924c6d57a544a750165c013564065a134592dab6209a9ddedf2b250f298a7b145517a87e8c930fb0ced07a0a133204464e585f8816a9a82ad8d6bf158f4521d324bb856f03c1eacd50f34d1fbd7499efea3aeb2a90e39cdceaa69c64f5437bcb359e3bc55ce4d0ce12799d2aa15f35a06bc957f2d1b4e725;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h5e0c5ec15ac7b2c622d80467d59a3d5a06dd4e768e8f25b0022f7cb4dbbd2b9909aa0ffad2ebfce61707adde6bf0a0b97a8e06d82a4821fcd73cb6d4f2b7d2e20058a81fb4364d3e519da07e078731f3d19f550e994eb855eac919e40f165b58930c85a4ef36c13cec4673d386f712f32c0370aed3647be7413ce870c3fc19bd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hc14e33b351c8f118f55dd2792b76fb364d6ef267ce6132fb1a0a91f0904ccfd77504b6da5ada5f9930c3b3fa0ecedc8ef2151bdf548dab497d8d465705b5a47077405e63f2da9070fc470905009069d9501f8f0d74d5940a251c1550f2cbc75eeb198d0ae582bf7e3a9d72f3f72e223b33e1403976036bbb08bf68bc771de48d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hafad6fbaa5ddca9af73f23455f83c1e06b67bee8fe3d3bd8acf63164bd4d3c9f70149be024216951128d556cacea93d95897142485dc555e277f3cd782f6b81d48457d6fa9271d20e342e9cef054f0f843979f5a646063d3aed230215d6099ea7fb6e19798a90aa02a14ea3e008ef9d5c3b3136428334f9157ee042bbd57899b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h3a6b69bfd59f52434af972bf69239e718a3061eb534a098b36932088c1ea31c5d9cfc207392c314f4e076fc71314e78b7f2630ae53a49d754f05ed81f87b687487e796a85012dea3e875d1e4bc892252c37c095d17509abff9d55d2200f44459a7f2a13701d8db0e6fcbda88f17231fbacb50ab056faacafc34cbb30bbd56a66;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'hfeec10f6fa5fa1980a96f1f78d656a70b2277e3b4ea01f8249be7cba86d36e76a186e48370e92ff7f2295c76658a01f0838bdf45f422d048566ff9372d72880477e2621e521def87e957529f3d551fa62960e0e31feb760f8e7667c264cdda1ae3bd1a938ab4247a4a1aa5e4230ded5c7e0ade4fdbec1f848b01f48bab945b1c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 1024'h6a9d5a1d6917c024d50d8221192ee89ec927fef0abdff2b214afdbc9899215f40884a0712192241e1fc62f257ae506a5bffca4581d3180c0736beff1ac0460eec67cfc9c38c1302cf73d3683873cf6a1557ea067e3d16c8d18683fa95202c340c47761c80f261c4d4cd7fe23366ca86589a044709f4204d798c7254963ea3a96;
        #1
        $finish();
    end
endmodule
