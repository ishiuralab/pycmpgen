module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [10:0] src12;
    reg [9:0] src13;
    reg [8:0] src14;
    reg [7:0] src15;
    reg [6:0] src16;
    reg [5:0] src17;
    reg [4:0] src18;
    reg [3:0] src19;
    reg [2:0] src20;
    reg [1:0] src21;
    reg [0:0] src22;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [23:0] srcsum;
    wire [23:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3])<<19) + ((src20[0] + src20[1] + src20[2])<<20) + ((src21[0] + src21[1])<<21) + ((src22[0])<<22);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hffffffffffffffffffffffffffffffffffff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f961cf432e887c73c902bf36ce496d7489b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7825ee8079d34b47e9e39560d2473a3df22;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb396a230990fdc8afea3e0f8cd2fe05e2ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf673f0788e84925ca9a83ef4ab11c7424c07;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9449e37f0d79fec31a76ddeb75bba4ee0225;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60e409c1edd773e4eb705b8a6a0216e7042e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he77d7afb7280a2adcd9250cd389170cc85a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h863dc4ab405869ff98557ac837a368d57ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81d37cb14588eb6add99743a00d6b89960e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5bd722f20d45a110d63a4789f0532e33b324;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc00e77d26808feb2153c7ac0bd2ca3ec3fcd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5a313fd1f409ae7e2aefc806ead92c0b49c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he07e39882328532f131bf24c08b6bd064768;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd45576334bdc044a9a58a0106f66d124cb80;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h145a661d56f9f1f6c50fba728923707ecc7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha23289791257dc841d01e3bb76487fed3538;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6a9d69a27565d927ef8e17c95fa15aea4a15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea4ba90763f057038e56c39c5e74a94bf294;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0b79814fc1e1b47c568959116d77c0f169c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc39b7fb17b07a366344341854c5d808e0ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab5d13defb7a26322742742ae78dc4286bbf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee1c9ffcbfdacb88575107a1b0634ef977fc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd292228e237218bb01f456138c59a550673d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1360f2242aaf73c9de8a42bd66c30dfcd562;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8bbf8c30251b0d926bb28f3e5f98591b685d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde3c3f3186c0d2e81703bdaea9cb11ad5f2c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha63189f1484c0e982815e37a631d443a3931;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h92eead07fa78e75917c101f635b64bc18396;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc916a6442bd8bd35116631a9a46664dbc331;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7ea11ad661a1aa864f940b220f2eee668645;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he129bf7e0b96cc0478c98cb200b922f479f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h433ebd5fd007aac09edfe3eb6acf22d6d5f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea1391b9f7da66c8afea64bdf415409b5d59;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb816218284cca94ce235764f3cdd77f4faf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h303a953c52842381ce721d427fb187e4c98b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a88989a1cad40e13fca22429d5ecff9168;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hccda9e39085c3dcbc2463f7ee83a9743847d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb7e7eff370bd185672b1151689462e6bbb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d493b3a72781a7d463f778042bd6e9f6b41;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1da18a9b103b5bc3720993cc79d4bddc1a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8bdf129788e92a206094f4b2a40b88a3baa6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c3f528abc13030a681ed47b67311ae96687;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb801f5662adc71ca5e2d79bd378217d9bf6b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb561040cc97abdeb6c094b3b35c01e6a3253;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4632d275e9b8accf352f9c60edc326afa2d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9cb1cfc5fa169bddb48b6b1bb5fe8d8e8c3c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f9268a913469e6b6c1fd1fe1ad3b43e88b4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7c1b0f29040aa9236b29aead6c70a9c673f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d580f026924cf2bfdd7c395deaed354a367;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hddb64248702a36d080e160df099cfe198931;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha47bf693a8f3430cc5951dae3c92e5db097c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbfaecd98adcf09af6fbcd3096a386741376;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h667f146a09c7d1e2f6672eeae02feb89ac5c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha768d43f33e3968b92e8d1c6d9019b28d301;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda32c81d30fa61ae8d7bcae80716ac78fb68;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe5ada7261b57504986a933c0ccc22c2a38f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e4edaaf4b222746427f7a01291c04c5305;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45164b72fbaabde63ac5b9d856de47251a2e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h924b2653377d8cbd2d11a91839f067e2e1b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he9fb2f46efad3ceeae30342f8c03c70df6e7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd9fe7bc9dd67e114d3f7d84b70fa61fedea;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7de969e2a2b46c5361d42a8aea1e07646ace;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he01f684da0d2d0ec07d6b9385d085b71fcb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h48078f051f6868540273497f3bb5b52119c0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc405ba88f1476f426281f47513d4808e23e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h837a50064b48fe2d60967257d8a3ee2fd9d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40138abb7c6b1fdc46024b93e8b70d78cb17;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf48a44724669a62846378f78468e05eaeaba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7dd58195cb7171248479202bc3756ac840bf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hac9e5b9fbf1c84d01f87377d9f3abae39246;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc8d3b19b106cd81e6176f54824e11516174;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc5ef8b883ecacfdb9bca9185338f415de7d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d0ca899ac345cee6b84e63ac56714462356;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbb1fbc01e9fd13afc77db34a4d17da28fc00;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbce477592430393bee7c25976ff22376d61f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58abb301071b1cce0925e7464d4ab56a2e84;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf686ebbc9a1bab28bfc8fa8ed68e3f8cbd68;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc2e7d53420bfbf640fb8e6b58a6b291d61f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfba9abd2d535bb7cff542b5bd3e5307db914;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e791463b547d71e43ee5665d4918d3ca5f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h885846029e797fa4cef813608f13daf42735;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he6fa99c5c74a20b106939a90111cbeb0531f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37da7972828d65c94450400e26bcaa4eeefb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h28a2832a9b60fdf217b748571bc3449c6689;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4728ad2eb23f15debbe436b3cee3624a45a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e8e17f0cd6d60479f98bc058005c9de3f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h38b99463f3876c570edc091567f5d8b78a7e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a2bbed8d0b8ce570b26373895e1d0dce9c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5eb70038292fe0b6567d01b89856c5f7785c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdef23dc4a0951638e9ca266bbd45f74067c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf63ccd92b45c53f7113e7e1bcb1b2ddebac9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc8e7dc02d25cd13f9b4cbcda602106db57e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd6933385499a50886511ac024e557140a284;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6fc51df70ec01c9de1afbe58cb8ffa40fd29;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40cfe8df8bbda6fdec0c51a5eeaed54aae2a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h17f31002471b50bf1756d22a6d2eab4a581d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he51f2b57b4b62fdbf6fbf86d8a2c66e61b68;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf1cc78d0dd6c065be290e13591a4e7d970a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ca0151113d1976f0ffdb54bea09a1f37d64;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55271b52af465f5c0690bbc97423805fb82;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ca2e2127f7a68d7bb358668d39ccd010edb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h821a39a01bbf350d704224555bde4710dbd4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h742564dd31954f9816dc6ec4f8c93291ece8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h52f1db8055b5744d2b831c6e461a562a588f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca89588363de44b69ef1827332d4655c1c14;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h460f569baa74665dd98fdac68440ff77ad8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd2364a80520adf104170f6f040c1f30450a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ef412b17182fb18334b4c852c4aed394d3f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ad1e1c926e6557fba30e7e2ed306655cfa8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed642b1b743a824e61c9a08a92219ddc07d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h187249f767a2521024776487cf88eec8e697;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5adc1fbc4182a7443e0e654d01e77b59567a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h290fa657e37a7d476178e03d84c664449b93;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5cd892cb2eab23fd2438bea40743ec41906;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h202d8e99120755adad3ea049cba2a67515ed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5edae91d0cee61e69c18a7a0d13c16d8f609;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b7ede568006b0d8615eefc6f6d8f86b68b2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfe3f7c115402c11805687e0d08fa90d0408b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf83a824f145fc9d13c4bd261fc79144134e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb30d03a66a330fa06e29df3d3b51ccf6d53c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'habb4fdbd2bef7a5b9756481cb93ce5f95432;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf5280eb73d5bca831e8b4d852f1bff9b194;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb567f87c01c72f501c770c05611f74f5693f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb0b6cc96b3c2e4fd5e5810eeafaeeb2e39c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7ffefa5b02dd1ef7d13de7fa1f075284364;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb50624a551e7b58cb971deeee9547ae68d40;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2fd076b8268afd4aa26b5a78578a950c19e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d749afcc4edaf3d3394a7a694cb445421ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf18b190e3d38af92d7cf561b084e546ac89b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5e07dbbdc26dc3f3ebc5ae18bc826ef559c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hccaee8876277ad82f199064e212d9db692ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf218c33af674bdc6d0b5aa68cebeaefcd81d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h78282d137495963cb32d222b6c5d72a59fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2dabd1e056f2f97e105e85012c95a02da3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7810a321a6c450eff03331aa2c590fd9a76d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h503ea48a75e177c7e47f798cbf983ea59742;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1af6029b62eb61502f47b047072ed5b3db37;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h228ff825aede20486bae1efda22c316f9080;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h207f58ab171414a385d93cc9fd754419d5ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f1511b0dc557c42691c8d239103b5fe47d9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd5a8629659d9c5380b783ec9cd449e6c203;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h78b30b191ccb3905ff50b267934f8cf2231f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54803bbbc80dad5740b7d23bacc7692dfca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcf312741639d25df28d761b2d5c0a2f2873d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h706741773aa4d0791e7311e3902ad3e556ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc4416d5dbabdf224efa83d31e4fc60f6f078;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he33f87981ff202e55676e6587ff8229cc136;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc43649c81429fc92e381dd2f92101adf27;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c3c56d2c52e2656bb6a034b2eafaf43203e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h302c6f02bdddeb8a70fbd90b847b8911bba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h66533c0606045ed92c79dc914def77ef1f44;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a6ee59dfcc0dac35d8ded01158a6cd092a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h83fb522ad543cd4891aec074689702575f62;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6158a0bfc1a48d96e641fdccf7bcbad4c73c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9afb002993fbb7940fdb2808757ce5801dfa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd097c65474b141d07bebdb7eb2d9186c6ab6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd910b92bc7140241353452b7a21d05880a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8277607f6df0f6837bb8cfb405980425b7c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he6830c6af8ea7817c82eba9605a0083959c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d35701cac217975e3f654837015c9a6fb5f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd70970be1a0179521af197d3aa731abbf12f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7be99cd869c2c96fea39de220abb7c4544d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2f4cc6ab25a6e3c03335efd5cdc7a598f47;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd681bc226e3a66189e564ab30dc0fd6c658;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h651717ec93f4835a052e94def2fd12045194;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f24fbeecd8935e35d1098432c3d92d0dd65;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h992a5fd3eb0627286ce82c39272ab9a7e9f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h86c99c66b4882d4f3f28bc43bc06aebd5656;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a4a9c240ce5a7c6410100c34f3ef9271356;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6fdd5ba724116c072fdfd05a281a41704bad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdaae584b25f4f570d0578091aae11a1721f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c021e90cbd2fba01d85120eba3384c1f509;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h972e2ed0fc392dc04340cb63d8faed1ad4d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h24d2e5d109e4272d6a04d070e93bd1a802b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14d3a0356f96c89890064427714f9438ff06;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5032165c6a8b8d55bbdb4a4fa7ce3ea1c34b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6564580efe9768d3baaf6af1887e0da8c4e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1ffc3a2503240f76a32d8733791844e9f8a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb0329bbf3b2d859e9208a3b6d8008b36bdf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8dec9dcba06a5d88ed913cb1391f95c07707;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2264b1fc664686da5423fbcf750fd99f710a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf29e3bdd738d7754c65a8512e36fd2834024;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec60d7a0e17f3d72b819830975d9ce19ed1f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6df2cebf38c5e6f02730711743edf7066f77;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcbc8a1501b79e8f089c72c7fa4c28c41e242;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb6de76ed9e839780c19396df3e8843f7baa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he77d0d19a0146f24d1bd3c6305908279b574;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha6a51420257dd11381437ca79fcbac6928d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec54c73459ecad8c5fd04dca2cca0601adf6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb138ef18d414e5e285eb09c47bd455389a3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h83112da6d91cbaac137590aad3c973b6e66d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f758085de13cf67df109010eb41364a7233;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he9b6900f91d7e98a30bc2256b8267dc2808c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1244839d993a501e45924a5c8d8421416c8a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2f86634340e3ee670fa8fe7e7bfbc76f087f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4d9bc2624cb15a20459deb786a5d48c510e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4e648f3b3d62f84a7527c43cd8815a52ad5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h64e4d5d2746d16a7a118ec32f1843e25213f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58b63206378c6a597ec64cb4cc49c3c933b2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a256063df67662a3078ac8fa22a14aae1e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63e6a8028baa3815afa546bb3824a19aaec3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9a9eceb6b5d0f716a5e842cfb47369a325;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14fae0fc384e6b23ec46199e2471c456fecc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94960ff32165e5591688b5df19a2b9150691;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42f497b66065bcab04766f769427d245f33a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f9dd42a2f3d08dcae6e4151b24c66cf270;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13817e87c2d0eb12ca49096e8e630f1658e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcccbeee1cd11db5f42d333d4283a2088d90a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d197f82836124d3836de70b2ccdbd6314da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35110a31a95ad942d29228ce43dddc8f0cfb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he928022c2d2992c38d58d9fc4ca801337603;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c0d0509f49a7c0053f62173229cd96381cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d55d48c8d7ece6159068fd4d56bb6e51c4f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3174f224a62a8468cb0780a346e8a1d6b179;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h774608426b62215a644021484aa43bb47926;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h644ba1e0d517fcf974dbe7ce022e7088b21f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ee1d8ab412b67383b27782b4447eb4dee7c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e537c9118665689d2f6c038c77f07f83912;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc585d3ddd28cf03652a5b1541d573256fd33;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9abb11883294958de29dd374697c4c9ee8f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd7e38d909b790a6f6228cdfb6a2993f1375;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7418b48bb421a1c82fbb21e539d7fdd08b2a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16840dd2b8c983bfcff69903044dc0e93860;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14aba64e04b8bc537e6919abb7c4d2696779;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1933aeecd10055d0cb0b74a39ee5393d9c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h40d74825c5ce47f163ed0f579528369ddc02;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8541483a917353913064776aba31f10a3f29;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e8c5c9ec3144317f6f7acb89049dc427623;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3d83cd1dcbdf372fa1a5319791cc61a567e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbd7570b345fcbb40e15cd50aa26f6b095a7e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7f5cc9d7a7e0353dc88e616b2f34aa66724;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7507da1ec9fe74dc6031fdd24c7aef4c3aba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcac218fab6a297b49fe184cf1c5d51d78053;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc8f5b3ec5c312fb08a097e6bf043ebc0cb3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9920aeda6b0c8dba68254d219f949f0783e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2692610b319439ae34d5a332cb078bb4be30;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69623b3ca97bab81780a4888de48ab022794;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7f0d9350adc607f02da8d81c98e51a5a61;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2c1960d2d33ebc4e828a8a225621401da79a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h458374da90a35fa2c53744d0edbac564487d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6526b85e75a0ddbee8aeaf8e5dde08d7bb28;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82144febbd4ee8e416908075219ff1e60d37;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h731499933de79321a0b605b3ad136cb4bf3a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba1d6bfe4814ee42c739d9a67156f9a15700;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he658b2c4357c0147ed22b354df1fe03dffe8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d4275e17acebd829cd9176bf4d513ac4484;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h92654fe69701842541a1d07265bd0d370efd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d673a708ad72f42d57cb2f72648b13d2808;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9921325dab7073339da37f0cc645a9e35482;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3661f8fcace996e8f9906e202fee485c25cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe2c07a8f89fc10527304af06c2d16b1c15b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70561d3ead7ac969802973959397daf69191;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34a28e830dee230a420fee05064764d260d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d2d711b5ddf5cd00a70e842bf8196ad3699;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he6a687576cfade492512f101475c6bc7c2d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73c8da8757914585e64d2e3277c16974fa99;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2b13476872314824ac3dab165164e2478d2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h93f786fbb07feba731753ad5c2c3647258c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf0ab2fe2262c9c8d072a4157c9bdc2904cae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h24a69caa2aea63abe74a6756e99cec27c6a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61396fbd979ac2e8f5cdf98b78b18437644c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb74c5ea6931f8d7729b885ac7899f44aa00;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b66fd29dd4dc89917d9010a81eb3debd38c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h841a809c96bb2ff2fce18fd068582439aa7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h75acd39737d42fb67eb25df9320f3c995b1f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h984c37be44eff63cc3afaad5c37e6f240c7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b454fc80071adff498a15f52467457e236e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5228e9a3b457777954f65f090f6c48c0ccb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6caa359a538f92fd1b580ad8a0cec2b0af65;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1feaef44cbfa0d35b251dde0a85f9bba1ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d1bda7272f8ba07f441ad6ff8c9eb2faea7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd76b55db0aa63cf745d332318ba66691b73;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h45ef052548b4d02e6bc25fafe81687a7dc6e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a1730247047e6d496448253d07ddfd4d028;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h52b990883b7a032518fc1e3c191966decbc8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10c193384e87b8a3a56df22129d31ec18c12;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee039c427e7fede767fd2faeb60dd9b76c24;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa7e4fd8a6f3b9e25808c3f8ed63e1bbbdc0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7160019965a1f10cabae868a3b973465fed1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ec2718fe8b96c0afa7dfbe2fe6e6be8e652;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ef4f9440804f1bd5a8ad5d11177a08d6dcb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he9d301cfeffbfe31eceeb672eed546b5df4e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h49ecef0080c2a79e8896710bba234f4a85da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h174080f2818f3cb3887eab0439a5a2dc00f0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe56040a6253cd0e51d1dfa73a8b06b41567;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd3e4932b846e25cb5cc6f935059c1a5d3068;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f98f981b7c6f8a097ec28c1489a40f78778;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc754604d1d4bb606f8bff2d25cc8d07c443;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef32a0d52699da28d316bffb50f3e338cd61;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc0c008f28747ff86e6156995391b8889d605;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb2b63c0fba5bd1c01bb848d5cd6d874facc9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he9af2fef0a231d0539fa90e2514ed9036b15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6d674309c5584c7a2fada4c88fb596cfcf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h751a7191abbdc8c7fe455ad6457f940a8759;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ef526d7accc7f668c890dd485c457cda005;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h841a72e11b6df47f8a7e24c58ed7c25a6566;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb3221726a9422fc264ff47269f657fa8b77;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h177fc91ee38a83ac9a0e33295000c83255c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a6c234124da472694c6d437af57729b18db;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25efa295a728a3c8391c7fdb6b9aab6904f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h49b398ec02b003629b7878ee70192a88e76c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a004197d732bc02de89937d5f4d060df4e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd8f1090f6a8fb6561cb7c8b6a64ef07d1e48;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1278eaf153563bb2cf76683bd456fc3266c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8793f17ca21f8d6c1b0a358d3805b501603d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa919e02bba35e8e91e869369a7a336fbc23;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8f874bf9852642831f2a1e36cb0d3a1646cf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h381ea4ee228322623b0e0e7dd5ae1b37f498;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7bb3c4245f8e082dac6af296025ca36fc396;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b2556ea3317c7c7f28d799ad8fc1f2518f5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1cc83c2711bd5705912831c95158faf5484e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd8a1bbce50b57defa213066f6bb133312f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha74c1f44e45c5490a75ff3aaa41b9ac4a8b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h61b4e362639680cf25fabc2b9f59752b2a34;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10248e836033858ada24f3e322c1f39ac95a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha183676bcb1483d2a40e1f7ed326292eb036;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b779ca058b4b5bb728e861fb187f266a767;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd66b758c78a305b11fb12c4d0d464b13d9a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3bea4e814ea9fd53a38a73407f9cd2189d0a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6abe84bdeed68bdbe75117c542178b179a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b79903cc96630e8cbd2570b5d4223ca47bb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h648cccba70721469f9c3a0794d7003ff2873;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h85cde5d9d7c3ab8f9718f9afbd33c7e12432;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hafbc662a7b1de9534b5a7d6bc057ae5f5063;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h277b5c72dd5b0d5c737d4e11fb220287e27b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda37aea4b95f19c66cc5baad67dfec221bf0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5ebaf29cad655497b11a0b713704625d349;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91bb00ea11e21488c37c47d7995d2c2930ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d3d282296681fbd94c326d41fea55213;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce336cb26a043c9022822d3fd6572c86944a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3d7668316cdd887f2341ef4b68dcdc90d6f6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a51bc2a98568123ef39cb7b983945c9fccf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb62f4b14d0341cb48ebac9228faa5fbe91fe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3409392ca257c8c9060510b7d8366623da1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee394cdc444b694194c016b984747faaa004;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b70a6c997cd727b1e3849101c755a5406b7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74aa22811f195737c3a4315138bf3f4af5fc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hed29286eb698b217a637f7f78cf7910b70a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56a7db8e816ba7580c3c13cc622f456b6a6c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b19bd9b12be26ab18e083bf121a29e5c1c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb3929f38ec707aa7a796eaf9e1a88047324;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbd0e137617c08c335964e9ee43e535fd8f16;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd88b787fee903467ade5c52fba3163dfbf5d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha88754c5234c46f7421eba0e89889e10135b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc59c6eb4b3c1c6f8252a87e7671ef43a751;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h16f429c2779642eda961a2a796036b234f06;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f10204716af98627b591f8de907cb721d3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf84acc72f1c67a31c67d0679a66472ce5f64;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda8419293ef4dc98b87ccec641460b59ff6f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda5bb53530581da931fbbd566a4b895618ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hea58a5caa3eb863eca5d609b4e292b351dc9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3af11ef5511d4276bd99c92dea845da1922e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4b5b3c3289dedad9a8d3c95a23bd6d7bcc6f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ebe52dd7bdd79daec8a9e62a3f6fafd6979;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13a9f3e708e9d14772a9a2330703cdfd8f45;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3828edf6e6bc434be3b5674eb3b6e6aaefa8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53ae1366a4b7548529367ab3000db638e010;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h27ea362138a3804be9cf56c2286ad8737200;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h927c7b2e94b9a6ed3933740119465ca01c7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d34a87d137a4ab3851e5db4ca3c7aaa63a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd1a5e0151f8a71d53a68a5aa862b3c765644;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c9a7c2d124dcb475d37b1277687a138674f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h96940379442c08f343bb2dc46adcb56ad7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h95d7ecc5dbeb11be5a56f799c7cdca55de16;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e6034a85a84b5d9b515f5eecdb21e1170b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d1c4249bf3750a0a74c3500435608f2f6ff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f30ab19df38d4f4640d0337484252e01aef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e14a0438d4c290c477c399e344dbf79bd6b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9353ad07f6859c452d96d8e7da0ed17a5b6d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb22418ff9bbe72406c87e7f5baa936a3419;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f2a3649c0aee210bf14605bbead913545b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb7e3c25d9ae2a3aa56cb59a159a5ad38eb3d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h49cba72ef290307be51e3bc2c2f4bd4d38d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h66fdccc0c373efdd80bb1701f457fefbd199;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h174827a5dff5b82203255d94599379ebe424;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb75d34c27f0bbbd0e02bd1b8393a0bfd7547;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2d9664bda3f23e5eb40a4015e1c6d2a2ea5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa40d471c08be6f7ca5a7762be77d1a21458;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c4f32dad39a973123f449b7b8cbc36eb8f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc818bf8d6f86a03ce6a8279f1c979d7aacc6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd7864da14a9d3f158ea976e126e5fb9a07d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h75ea82536fbe42deacf5f594a02266afd032;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h124ff170282abbd83240db519f9443a3fff7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94c9f349d9ddc31b405165f2695a35873a4c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f122d2c234addb47ef27bf6a9a4b02d873e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h519b86e43ad7c7a952512d8df864f73e1a5a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2dc1d5608c9efd746acfedf87e8e7c2d2183;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b9ce73524d61cd83bbb8204d96c69d0e3f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h38d3b482e21fcc04a8d8a1c96da5dc37c607;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44fc74cc28bca87a6eda403219684952c8e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h66612b2502d6a8e385a17cd5a521de074c15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6f45aae6f0a26bf1446924b2ea5de4c16cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c91e016b78531a10266fec71421e63ea701;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb61c73ec347b58098f717eb61c9126bd6862;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7511a4ee016546dd182e64dd526015def16;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74e8049bb7de0ab770d986d8ff5bc42019e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h36bb49223f489928fccb53cd01dcbe261dda;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he27738230e473fd951a4c666e6c7bffb94d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11704ba08643bd77def59cb78f309bf9a012;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heb6d2f11a64f8680f0fcf8fbb6fc5d9a4733;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99aef8fc7048d6d601d2d4d42ecae88b97a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84a7b31d6c63e3e090b8219f9e04f87e7b7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h669f554c046b37852d613d24465017b546fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h75555be776a6f3b3822c889a21e4bd07bb66;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd40572c64c5b021442b6b9c36a8db8510c63;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a9d24a50f08dfe2926371355e30d03a4b25;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc460788b1bce9afecbb16dcc52c138f2470a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3cc422e70ba577b88a85077c54bb60f1d9e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4cee4e4faf5a71a35d094305505ef4384c15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h19aeaa55fbd9bfacf66f45b0352b63af047a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb242c84ed7e146bf5c2352cc4c9193c8fe04;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h17d05afa668a3da00649f80f71fa6a62c269;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99235a1dc46944ba2faad2d95f078b4cc38f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha445b14b886b2d4441303eed63b54339249e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e0f88f656290399a91c94e5b19e4b3f43a3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf0c204bba370ccb2a845370bf89339320a65;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h97e23deaf2fe331ee0ffa6f3131f7b7d132e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4045a28a65cda8cb665a47f79119a873a818;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h96ed54de3300b604a6e8ad028b22ef9c907d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6ad6b54cebacd3dbf1bd5c3ba6b3d97e889;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h67e2ee24249d108ff592ddffd0a13af848ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf6cb90c97d07c175acd97e1ada54862a5273;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77366d7693a5ad73884cc02ec0794c5b86d5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37fbb20d08609fd61acae87482160d5b5f13;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h998493d8cf4da3326d4f0fe8543e3fe9576a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa939b3a4410d42a65037f62245537305616;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7989ea9696dd9304cbf961d90413ab18cf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h65336c50ac6e6b6aae40dcd5402a62e31385;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha03b87fab8aea6d42e1f11d61b877c040b09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98ff075ea85b30e02b7b2480e8502a49b0a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4a9f4c054e82ebdab25077ccc201ed5948cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcc8ed8182d8d0f80ac06618ed8d36fd1ff0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h548fcb56f69e60f167c611fabd392c002383;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9b0615edbcd94aaa9839a1978152b7552831;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he402b2970e35ad372cff9b89cb0f2a49c596;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6cd59742ae9c26f298c7c5f53d18b8ecb624;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb985045f48057304c271e523cf4e2a4a63ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb168ef20edfa84faf95f97e94f628c2b8c15;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ee38b0c24037d57e860a129ac4e060f60f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd9581dc5f87a87e1847cc517e351d442f0ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h373a49a074fbe7aae372508f6fc3632f9ad3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha367dcf1e53045c9bff21c6979f5027e2e67;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha105bb9ddc393fd3a101cc1ef0facf60b18a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c1fe3775af70df8c8d7dc49cc0bdab59eee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he4e2ec1163c32dfeb5eacce167de204ae5ee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f341c83a3c939ce5b70cefbd341a8e38cf8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba8166ef85632a697d19797b8afacf40772;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb2e31b5ca596a358bf02202bc7c7b89985d9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he857d8863c2debb619b5a65a9dcae0fcc7f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1cd70cf1cf5a6b4e664d306a39ef25be1b78;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f962f5e4fe140d9dd568dc893f5c569a31f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8223a6575c86917c0ad7547394711845b235;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hefd0e877b7ad02491f8f47a60f7c47c2e271;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he522222df6ec8075fc72501ba3250d69acc4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb04081346b02befdee791f76f7c280ad80b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d8c3d2574734745c343388b77e5c919e90b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1c3b0f66f8726a799948e512a5c2f8985c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h742a8fee098cd4bba671577c7fd042fbe990;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h78d115713b2b94dd1e300d56f5749dd78968;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5386cbfa0acfa24a4a59d9b10bc890edcd70;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf57d0489b905101cdc5053803bbeb2786aa5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf03af0d7bf75acc51a7f9a63ee7876a10778;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfd917f7a488e0b310eb86aca49fc09a360d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdb4802f841962deef7e5b315432e8e15f0ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h884ad88cb2ba48c81ceb043843c2efb07e8e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h89815696269fc873f8d0595f19693c8ea3ab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h80b44e2943f48321bd14d75a8d0c9d0a78c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2abfb9b697b5edea2032e0c414f55865e543;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b9ec44ce04784d204a13a62f15aaa530548;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he0f7da7eddce10230a1f52a13063a45723d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a84daf46e1ab6e463c305e35141dac2532c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdfc8fd7275af01541496596120e34afc44fa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb77e0c6a39c7acecf8c60b96d700385677f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h576f088256e6a765d444bc7e2b27908ce964;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc2975523c75df63070f2a05ee00a46fb9d6a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda90f02b523a6c5864645d25dac8a9d344b7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4162e72e26c55407d7d88c1934f254ebf82d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6623e5881beb8cc8a50b81e6c3d507a87d22;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5ee130f203f76709cd3bfa859083f9f2788a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7b2b79d30443d907e73733374705decccfe1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h69a48680220ecb6de8de343c678e0130fa6e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h285faffba2c81214d97b73fb5b91e1c39218;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54e427ec6785c4ab35e4fd7c9b67c7efc466;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h242cf99a25e60aaa3e3fcc54439155dc7235;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h797fb351cfbe994942768ec7e67c4b2c6d52;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he446172109218afb3e6c51ee866b498e9220;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6078f240877a8446396498793bbe3bc20b35;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7361b5648e4dec5c9cf64e89a177d200dd1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb4be092b9acc10d268e389ebaa84db770d52;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf235efd2b93f9daaf7d77b0c6eb61203fc66;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2b5f9e5c9885e8b6b1d33473be627a7c3bc9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6258dbdd2f544b72f13308276c933a7884c3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbb3f0a5d80793ea3e01abda371fa6f5bd47a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c67dd1428cd484bb3e3eb3baccd56a5369b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb0a18660d45eb860f83f6e84450c07dfc6e2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h272ebcdc7f123599a4f3a0e533b4098113e0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb5b0c6171efbc5b6743fb019c48f5e12226e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1bdbfb4ce63702f17ab546391fdcc53d245;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha5ee345dc185bb9e66bfba95e9e29fd6b258;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37a1a6305f9e22a82a0ab18c8442868ee1a5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2d347c64d3c6e8dc7a19ff78d9ec146366ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcfce476aa342cea416fdd192a09e5cc4608e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8672ac4cfbe53b71c18890d662baf9bc58c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h50726578200dc220a71d6c16f5c5b89345e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha536cceaa85963d2d079936a7c65381148f3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haddbf04ab2a34d3c2af549becab336aad334;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h68dcbcce59c2a605e403ddabecb9ed3f121f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7fe4b8ee982ce26d694b3252cbb026710dec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8bb609f8ad4abf5576749229649b4e7707ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1abd3ad4785571a4f5f4ab39e39325e58881;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99ec5a0a7c74081e941786254940e4c0e389;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf5938d2b5481cab9a0ae3ff7d8664851d577;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d320726a73900c35866d5fa2a867dba5bd2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h339644a78171fd9ceb2cf37248fb87031d9e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf990dc09d0c3b12ab231918bbe2db82e4af5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h38f28d49a02c8c74fcfc3690ee9393584532;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf9232dee8a8afafcb46b9695ddd1b95c5fa6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63c3f6a998e46637848d3a3c9eabbebe5e5e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbab0cfa2fd20f9f1a4be2d4e358316725b82;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1ef0b09675bfbd75dd5970fae1d68d700b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h11a2e4cdc101bc99af5174673f0ad15fa811;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1c05d839415499f62ef9c0016aaec7eb2142;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h65af1d00326d8b61517bc50f3ff2be754f39;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf25a47f3b3f669da46aa00522aa7b47c51;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h752d043ea3e29a3be4c3907a15defa36d04d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7adadc7e9a885868d61cd8b13a464baf0430;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h43cc18f90e5ab0128d7075e118327ee36866;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h76ed51ea507e217bc04e0c7e91e0eab50e79;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37007b14ec275a418f52573bd764081ed702;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55e1fad96fdbad8da078d5aef8e972cbc907;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h224528b8f56cd081641765a98a574ac703b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd563296bc3620ea6ac0ea4aff42a70a98e31;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1760855f42136368d953cc049c678e2f212e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee048a9047b8472544569fcccd2ae0a0054;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5f66d330eccafb0072210a3fb52f9f5f7987;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hee539fb094eb982f9a969e822f6d3146a16b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33b94f3a2d96f7f0b72034dac0ec8dd02582;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h443b55e1e9f287c3fe4c95477f5fd4e0e3aa;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb53374c5546f8bc71621da399003732faab7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce510f93506424e6307dc9d04c18da3700c8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h208e75e045d42f8da5d53b36bd3db2e8473b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hded5135aff14ef9a47e021bc528f1dcd88ba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h96d1745cd75c303d3bde91b2f05df5780fb0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf924fcb3b9feae33a3167abdd9e429892099;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1849f63fc39bbb83a5670b4525bae314bfe3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9949a4f84fdbe7cc15dc5d97d2a63b53d54d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb854b3e3b02b1b2a1a8f0db6df9786eb9039;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1b12c6b16e7c478485410b3d4afda16a6700;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf568bff1ba96cf3a042d0ae83360cfb25f05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7edfcb195dced05419ad35b5a7c0adfcd8f8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ebe61004fb524bbdf109285b6af9ae253ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b6c1ffd6f5148f1ac96f5a87c6300b04b9b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4f670fc26c99e0bce8d03788045e70a8b92;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46561e802820189c3a08c6e721eb6248aeb3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa74db9fbae1efb439a742f8d602b22adf8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb1640cf5d4f2da98b8c0aa282187f28c7482;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd9ff8500e2626d72f784483c56e63f5af59e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7e994695a15d2b59f36c90f3b5e8f20492e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb5e169bae1935e87af56a2c067da3054ea8c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf14e8003348b6bc1d9141783455e65ffb20f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc739364b357b83e9c074a329716ae386a1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7b4e7efe9629ef97ce6ec4bdc75f91cdf6d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he63f61df2847aedf10018f1b1d40b0df653c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h47348583dee8072b31e66596e8bbf208632c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h299643d279b956c7fe28c46326dec581d41c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f42b934ef9db7ec42911e7f5ce6dd2af923;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hda1713606bf48e249c96b27b7d98b43b5ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7518faee52a1dee5f3db6b08051b0cee4868;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3a13d793fbeb871f30645e3c4a91158aed5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf6776b4333fea6a984eea71d158e37df52b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82888dc382fcdab9eddc6fc7ea0f2cbee571;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h230a9c590233c36e19c455175695afce7c0c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5454b95c7ec1826a2eb6a51e87737be8f6f2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4597e49204fbd22a242dc7b10f6453ab1436;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha79a8799d86204bd28b20106e2d3619771ca;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h400125af0c474e89d5f0229b437a4371f12;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc5cdd10a72c581225d8cb080a6bf2870da55;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h38c1460a869434e01a674f524d0bdc9327f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heabf1e0abf6ef4cbb01de59364e655cd408a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h27e1c147c43df24a40f25810653da9d22bf1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8195ec0b0ae771ce86536bace2dd39e70412;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h17d39ea278e0d25a3c2e3067621110dd5de8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h39f7561d65be6cf81a1c8aff0f404ad304c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha33ff739d50c68f0dc0b9697f0e3b8abe13a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h33d06e18b1f61acc71c7628a05b087208b0f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf535ce0270bba0765d373cf3312f5798782c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc8d28f088416bb9b9b2f5b71f96cfb1c5d18;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha53b8731cdcbcd92e9601fd62d7e0bb27b8a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6476b026ffcd74e2c31ffeb746d8bc29b47f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h327ff6516844e7f11c20d65458cb540d0003;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae685742c71fbef645b6a4b0f997a284e8e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h30b0d15e9c7eb93fb54fe762604c5de0d005;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h89517c4e4c8255cb5aa090b0af49ba7ea887;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7de97bb701b735b343519ac1f06e34dc0014;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he1ed26dc15e7206308f5608a07876fd9624a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hde77ad7764d17c01fa11744f9bc6fb937a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc88efd7146b05027ba5e4dfeb108150cd581;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h363db7e50e42f2cefc0a9aed782eb1f0783d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a30fd19d8881b76a315b7606caa80f2521a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb21b16e3d4df5be4b8083a512a4e69600b9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73891d7f1b0b275a7113124dcb40cdfbf3ff;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81293bf9a44684c866bb14392faab6ec7033;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5695733cfe1cfb812d89decbc615f1609592;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1a67fbbce7270d8e86fa895727d0492be610;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h48a603d528f787dbdd0811a9278072982b71;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60611ca7df8a4c0b7920251b46b17d3ca871;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h54e7f20c2db03f4356d7af6165eafa1713d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h56758a404d02a5328d2d0e4c64d4ee7fd7a3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h55f5fc481dece489213a82321c543c8ad40d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h485bb68edfd21838164cf056835b8f06bb77;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h26e97d58fd0b75b29c51b1dc7e5b26e42bf2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc4fe8ff0b3067e8681278fe283d7954b30ec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf17c534f1f239e088ace5ace816060b82540;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e48d1845e8cd9b4bd70debcc588550b18a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb370ee79d86bd4ed9934c942f2b9535499d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e41e4b2970b23e5fc18272d6060cba4244a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he432e8246970781828d1a6fb46d8e3c9cae4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbbfc1a4d7342343d020262c941acba2e2923;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h29fe31149a68a01d789139f8546b87f88e60;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8b400f05f2caf95d802976784861a8c6eafc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf841c71f7bc0adf0eb0ffb35f309075d1363;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ee595c4344fde128b3395f1bef38703b5b5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h15db4598723afaa0601bd380f16327c60be0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd97841fecae58db0747d170cdfe7da5e73b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha23e55570eaa5bb433b62d3c8a843ac564e9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46dce4c6ccb639506a54463066b17a189ea3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfca60a3e63c2266f65b9039718e4d680b6d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h869cd3d4e0773614bfe9450811e341782000;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h546117eb11675d2982d4723df953c2398c10;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h84cc25399b54d168408df0f55fb2a0a09a1f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h131980aab2399d6d202c7ca958790ec85bce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58bc48180674c55624e5455be27a3689e6d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd4ac4dbfab4c950989f9a170e931828eadaf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9dd1efe1fae45cf777943c0c137457ed93d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ba406808810e63b751394850f6db5f9a4b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha980c583a84b45c50f1f86935c0f7d15c381;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h474fd5085544adcdbc50f37d6d5002f1055a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbd626b1d7ad78ef162f05c5026f2cd5caecd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc063a54ea9a5e8a1df8806ebe33aa4531b4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c654b6cc9797f75260b4d5371059312c939;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1f5f9266e3b76f3631993210c85652fbed3c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf59c828b85dafdcf21e6e915aad903a7ed48;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h618f79347605b41cd0ef4ed840b84ab20a4a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8c5851dcb12c05b62b8db945c0c8d32b8869;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h182711d5b3f59e9899bbbe9d1de136b82823;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h18ba9b654141786696d3eb74ebdbc059d179;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfea20cadc46cee83e0f0e229f84f224bf40c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h262719d2ad1cb3254b49bd95853f6f2b5706;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73122065b957f82cdde901e65fa81e4bc663;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5212c4d1e02d2d3f5017e0018bf2bcf2214c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a0fe3afc03dd253e162d41b3e913de91b81;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5224e60267359729b140bea554e9bf417a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb4031e8f758db9091b6a487d6fa52b41f25;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9be456e1826f4f31f1e5bcddb8145d5fb9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5812def349e8f06ccdff6481197543645c43;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h736c0328b7809d1883d8fc0465e821de5c75;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7daf5147df2722ccaf45cca3ed738a80091e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h949d7d08a365289cc76c83563da70621ac09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h532462bcd72444a372b90f3e5f7cd238cc13;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h681a2114c80e3cd2cb99d8f622f23cf22062;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha0bcef26a8b4e36dba28577e09e7319f5ea5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf7f163884234957400310e2c804d2fe3f47;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h322ac667d8480a73060b83401ad55c571487;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3b1ad850d5b012babbfe0cb78c2d08cab7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb34091954fe78c12e67b3d4b1f2ccf18e68f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc09b102234fa2bf6c30bfe1fdd266c35014c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8fcf4e3bbb1846449f5d36e22af4ac3514e8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdcf1cc2e8072adde4cc86ae298b369be8516;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h455e55cd3331c6f10e5a52b884336958ff20;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h955130358179296ac85f8797cb5ff15f8788;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9fb52410577f77aaaf6cf829d5e59f3958f7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a56bf74ed887a58f4b02ce4bfef96c84485;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h58a15bd03c2d74d4508d9789925c8303cb8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e49329755d24e06a3442a37447c27e8ec1a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdf5662187b58e0bcf5afd392d4c42f2a04be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfafe45962c5a0c16b06584147caab955ae66;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c425435fc68b93955ffea1441f0abf06c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfda8d9f1808f60e6e2ecc0f25c23a282b58;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1010c7451009145d45e25ee8f2a5719febcc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5af59489d56ba931aeb0b05b60f4978c9d83;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h916aa53633db1a26ab127a93e410a077f6cf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'had2deec8b4afabc2dd044f48af6da1af03be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec67280e7a0e0f3b197b7ccb5231052f9bba;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd341c6df80a9d821d16d674fceadf89c42b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7ede32573e197c360edb0bb713ac0d9c0e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ae598d0ce6b7ae1b23b5b5070a2f0634b8e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h164bb35af6073aaa048234b23a2f362a253f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7754694962bef7562f35858683aded8ba25a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd5970939c89c162094b2fa1968c50d663a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc88fd6b487c3114dd4753324d08e6d8fddcf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d1647402aa82f04ddf483f1930dd301cee6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h46320be7af4de46b8fc1117742fcd68f6c7f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4c9493cff01e98a755e50c80c39eea641ec4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h32427eb62167ec8e032788b06276a991fd53;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9fdf21ceb000de39b198920ed55bf5b8a256;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f171bb26ad8fc086a9b71f125b65c486a85;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8207e0be8cce88924e87ec345599d88acff9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h904dd655990dc0200a7af66fca62ab709cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h37ab622f47425b3e91693baaf402b2c36d13;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1ee49d4da26146f41b3c539378997de19618;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h88d2faa062fe25c07a9b0baadf1926253316;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f5780ac5a19039e0e1316406733a9828de5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h988640f79dc1cd9d6af39b1f94417e4938be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h52deee9e8937c4307a66e6db2fcf8a86b0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbfb773bf308f68da85a6eb47a591244d69cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h66ecf3ed1809893b55b11cc8f3f9ab480c16;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hec1a18c09f00bb27261a2a78be56cd88ce37;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h784f360874263400ac55734371ea8b5708d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f22bba7a0a58705a9025fb34f8c8c7327e1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2ab8e86fd12c741f9736990c1ea7b2f5b836;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'habe3e7e128f8ed40f41bff8509e3580a0a17;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h57e40e13a79ce3f1cc0a6d37a9cd4bc88f05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4338a6e0561a119121aec0b9004d95fd78a2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6657578b48f54ca06bdab071df8d043fc27c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9c795a12b2d8dd18eea9aa7cb409017be01a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha3a49096a52d657fe92a4e91c668ea160f80;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd77088392494cd3e5be3715bb14f04e6fef1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6d56c38c12df34742fc240f82fd858f5f05b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he3f852df807305d75b71a8feb309e76fe3dd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haeaf77a27d7b059228002bda835fdc3e780b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h90b55863a9fa2de7a7a381818d341cf7edbe;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he011c823d5c657e4a53eb0840bdcd33d953d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfb93798e54da90bea379b645398bde27ae98;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h107a27e231e9f0cbfe082d7762e00bb5e76e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha4dcf68d92bc2e3ccbb6be3cee54f4f01401;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd97296829f409b79ceffb60c6b1e702f91d4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc460f2d9bf67a6407fe2300bb1a8abc38cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2bc80b240031ebe8caf07c4f23c67eb5c52;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef3f1cedebab4cd21f509be7f0beca71f88;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9076c7271c4523f89acdebecfe0ca793d4e5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h598b583340c8bef21bfa2f2856e6c7a4f523;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca45f87b6b5a89afe74ff33db69cac08614d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h91a1bbc5c9cba5d77d1e1e84a9490c94cb7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7a3b0e0e7a1025099003e1467ea55f072201;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb73bf2a56446adbad7d0173bc3feb4715854;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b956c7671350e10b204e91562b7d57d07e3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1701a90b0cf1d0c822fedcf22a999d5e26e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb5540a5fb71701e9ea6f01d6dcfe15e2880f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25949eb3d48159d0045ad5d855f80f92f73;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3473a537667f38d58558312ac90105a6a900;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h841d268f31f9022de8d5d859a2d0c31b995b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e0fb0668a2e87bb74541f6c61fe84eb75eb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87abcda8e17d1886050cbfffff742b219c0f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2aa2c95e96dd3b15ca3bd0f87f3efa8acd9e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h80a775fe6887761944a2908293f67ea0e785;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h60027907235773026b64e7708dfa2f6c031f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbb0de2d20d0431423bfa272c940f6762fd77;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44bd5c9eb6867fdb94429d4cdfeafbd04a70;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4ad1c280890bba7b351c633287152731f5ed;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae1ac9f5a0c8c0c9d7daf95ae40354b7e1c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha0fb319aa5d2f58db07fa280bae72a14c316;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44ef1edd25bf53484ff9eac03415e9ffa59a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h14166d048cf1752f3b96693c4326b077249e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3c66ee35f2fe4017d5ee1e5c22966d9c19da;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hef74bb50f3700ea8420a30bb596a83d3d9cd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h544e8f3f6c8561be8ef830c6e81210e96769;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4de50a7d6c41ebbf8b4336bac7b75a1acf45;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he5f8a1c6e8bb5f073bf3547b917b5c7570fb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfef50dcd210c95ddf3078ba83e9ca1007863;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e502aad9720293835f2f7032445cc89d341;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hadc66c6b6471f8049f881bd7164fa89ef8c9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hba8037d1a72ff9160731233f727abbbe274;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he87267d3e6945b582b03e8ea800389d0d5c2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34a28ebe5bde7bcb169043b8acaab1bb83f4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6cd35bcb5b9bc47a2ffa05fecbb6a7e62a59;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf11ef434fbb4ba15ff85e0837ee8e51f97a4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h87fe9090419b74cde2b9b8d3bdf35e26b8b7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf065d6f0787c16ce7510563b48b5dad9d804;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hae361ac591ecdf7d8eb813bb5f100af3af70;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he298f03ff1ea4f581ad2684a34305bd118ab;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd43454fabacea1ac1f7f3c6e59ddc79ebd4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd2161e49683ed2f9cac5ce08fdd2e7f23257;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcd40109acb1f2887316df482adc155964710;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c5eeb4b3bd7ad698607400517f12da5b391;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e7e2a0feb25e1aa5c62523949c981fa8cb9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h518483b4ee1cbd7ec46447539258bd9c41b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce2b9f97ef04a9ad8a30946a2a6d84cfc9b7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h938def5adafcf7744a1fe32e57c86b0864b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc9a6b0ef2cf62076db96c1e6119c8eee061a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h569123328cdfdf41a0ead40a7e50dab76e8c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6747b1631438fb5f18c64d7ae4a70252bdec;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h62763f3499f87bbb9918bfa1941ecc40fc28;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6accd9958c0d481851f97d29eb8f5ae9e092;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7961823f69853638fd193c5d2b4c543e15a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5b40400de38017d4ee27b0146809ae464c73;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf67a7493d6475b87066bf4f36fb4df3a0352;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc29a1b3b47e7a71d9ea73676077f521b3fd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9f12fe91732184c7cb24c94caf8bf96e4271;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7b6fbcbce150a0491525c0be01c00085f8b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h66604690cd0b278fdb9768826bd3e2bb52e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h20dfb2672dab67590b62ae154fb6f75a2beb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h294f406fd2b590d7c32a5419856461908da5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h909914c470810b8050715d72c8597b90b3df;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3efa0ef8ee41f77a405a821627357203a37c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'headea767686b0eeba3ff3230854ef1c799cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ad60ac957bf8f49f6352f224517fca4ead2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc4e4e83250246dc4e5ca4f222846a26b8195;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b960578053cf3cf5896c90baf107561e15f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfc1c070d64b646eb1e156afdcf7e60a2a57a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2173c27badd9d0832139251beac791ba90a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5dea18bb5df3e1057fb58604c66612bf86d9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb5bcac8f4608b3c81ce3eebb3cffe8c4f30c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcffc88b9a4ce50d97195d7fb1dd4905f816a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9bc0cb1a56a9f5ba92f1f2477223c1d0d45c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbec918dc23b5c8d77b464c70ba3568f7d8d9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc81e138962783d0af98ffa35973543362035;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc82fadfed54a7d0f2a56e094e5980843282c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf9d41a61ceed2a9553c7966769b9acc9f2ac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d130eb68dd886411a86bca9941a5afda066;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf6388695ff7e38f5c7ec11cd1bd22a0473f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a8801e7dd3014b6ee1bf84cc701084b6488;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h30067142063c585f7831c7e9a0a14db088b8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h98903061043c80a913a64e9ea03af3d607ce;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h538ab68d0e2c6407c08172274f919288e6de;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha70dae5b73e9e452605bd7edf7a9cb8e6122;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha84a48ac08cc206798df2a3ac26941149d7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4eb5af2925aedcb03ec8221992d7876d3584;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f90b575c34b77dec6f9a3ec7abc82e8dcd0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13f98ee473c6609b6982a3dad365d8a98548;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f7041b71f954fe20c14906639be43076530;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1adc166340d830f9b5606847db11beb69cc0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h185af34e62c353acac492c608e2278937abb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf9339c7123aafd011edc8c8d945766043f00;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b06b18fc088afbf916167bff79dd228a0e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hab643c3bcff7b9b37061d9afe3b1b19e19be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h25fbc71bf90fcdc8b704649ce86b0fcdc54a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb9e297f9d4c4bb23e78e99d7a633dc154085;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h80562e56a392fd108659e902d8d4524e9eee;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf7112fcae76ab818f538c8c280abfd89bc20;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7cf48aa044b99cd9b6843bd9bce7a7617fbd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd610f5dca1931e207204150dda7f0018dfc3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb19f107271e435a4b0339bd39c0fce58ab5d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4100777067dfe1843315824a00869919dd3e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hced7ed8395447f621de80556506ec756bc69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h369f14731f7e5ea12de28d0781b3ba57467b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb5c4b6e1c302be9fee86f13bc19353454888;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h987c133fc33055083e127ea76139fe0f80d6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6b4f888ded149b15a94bdc7b6450134eef82;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e27be7a760927290db3caa6392af896f548;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h74670f837e4d0113aa42b887e1d44cbf103c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haaeb9a46f40554fbd8d01def2500ea32e4a8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd8cb6b4336f83d48187379f4ccce3a524427;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d0744b9ce563b207ab444f5bc504d81983e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h81da8e9b73792151fb4f413456bed94bd59f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8fe5a67ed94c23219f39aecb866880941e0e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3ced6c853cbf6fd0047ca81c1b53bdf29873;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa19d9c068ccc408bfd7eaf0f1400eb82ce7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42cfb5086e4fa67606d51c67e1b6d962c1c4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9183a6fabd7bedce250dbf55a99bfcfa6c2c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7f21277091645658591e63969e4eeab41c3e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc713a2c61c528f0f8bc97473f2e2cb0f610f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2a699037eda95df3632a34015faf81c7c460;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb8ce8b350ef5f6fd09555a0b727a91bf7a8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf476fe672c0fcc91659102dfa7c8a6b4b2cc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f3bb9c6649d10440eaecf5755551003f28e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h665f74d248cce6ea7ba8403958c75d4be6cb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb9cfad82336437e3f17f3f1b14dc0d0499cf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h447f8035f1631ed981819ca6fd923b0ea511;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8d7a72ccdef387b0f2f4bf7c29f0f0003471;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8675238eeb2f8c886b7e6b042f883af28115;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h293218d8ac879452ea008faf09aca285b4f9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3a5d27042e5e4a3148c6f40be14c1336facd;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3e4b4b8cc3079c8749890745f80162cf9cae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd226c69e83d1fb90da83fbca107fee51e1b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'habb3a8823accfbfb32cb5548283c9077fc8d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc4750d745d8782a743ecdeb9d2ed817309d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4e11d44df49bfb627d56453a8a81f090e363;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7c0249670059dff1e7a6e3543ed5e513a08;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha8e96270360da2fdeda637e914eadc6f9537;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2bc2e3c19b9c64854836ecbeaac165871f39;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdc52dbf617385b7258f0286ebd9c071edc12;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc4a58dcb94a05434b3d9f83c308825c43db5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7675889c80d4d9d606f32e19dfb19ec1fb67;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7374f68cf4180ee9e36a5264c7af07f807b4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6bba3187547c6624f1d46c7a0300bb1fdf2e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb6ac8899fe6317a041a7a6e9aa70d88b027c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6ec84b68ddaa2346779d103515d56f064676;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6adeff2b92e01b755d6af35e0228a1b4eb22;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h299287a8a69a7d1ce6afe339470bc35e2dfb;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc03d82f64938e907c207a9209e215aa99e27;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7d995b97ad9e8800cd2e114cf13cb7a12a9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he607336c92defdd1a88a04eff97d3f0bdb6c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e42c86d03b2f15e6399f4742cbfd3823f7d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf602acaae8fa9f992f4f971a31fa41eea594;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b4294c5370a06943615c3d3ba24a4268cd5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h293dd0d2c67994271e52954f3db8152a5a21;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c5b3568d730c43551885b0e5bdc5b2fffc6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7e43fafde35a1ea0d1550fad76847988536b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdaee84b67e6b142d34405f6045130e9e830;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7320969e83502d889e40c77a85759e5d0ece;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ef19c23c163c2938c610153c0ff53c9c3e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6e5a2c6ebb828649352828cf2fa27f2f5670;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hce4a404c5d6398953461d90e90258dc88c5d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hdd4b2f4d83d1b4d9beb07d9e13d7779f5bb6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf1a340e9464c93a6d1532138cc61c35ae4be;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha9c44f82892feb294d66fd7410ffa1e46579;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf7def255c43748a35cd785099867bb6df60d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha93fc28f2901e66937ac9780192b0f8e7fbf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbbb0f2d4ec67fcdef75af0869f1e9f88b205;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb987552f1d79b5a8902e1e7d5cbe6adfd112;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4d434d5c0d4b6cdbc81146ff72619384f24c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h19df62cee51da04b0c4b32796aba01ea9c99;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hebd98898d02c110607e6accaadcd2df5aad8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5a60ef44ecc87e5fb60cefb0a3b760f76831;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h5cc4d92d1046022be39a7a59212123e2222d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3747aadb7e61caee076bb5379c8a7abf34e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf2c0ea488c6c6e43da30c575349e69d6614f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h273d53a4612be7f479c7191f1f178196bfac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc097e2d6bcb9250b5691077973fa1df23c4b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc6963755889db3a8412573398863c07e58c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbc4e836cfc5841218bb86da1837e3b018f92;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6faffa1f39b45fbdc318ce8026113fce9604;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf058d3e406aa6a8db5b04e090944ca7c2ed3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8bcdced6fe732e877004d6a1c653474292d7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9da440c1130eee877779f2b48f439fb0c21e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8e3f0e9eae4d83788fe8977a193fe600b91d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59fa28a5494ce4292d2c3d1cfb1acddf95c1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1e9eb3e41c5fccf53e5cbf37e9c20fa866a6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4bf5d6c39c3804232092522cc528ecff9717;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3af6f06c7cf1840af815fa29b437c9d5591;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h424cbfe51145e3916f153c17295811c90d82;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h158eb0f9ed049eda7cfdcc1901a302275120;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4431b4b780d62e0acfd58afdf5e590d15d78;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he422a90476aaad10e4d56b78198d6990e01f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h356031db7161f80ec483ca5435b3fac876c6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h63eb55f00a8c7d50c2767d846ee85bd93ec5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb796ec21296a5077f81c010e4ab86eac85e6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h96311f83df192e5ec521efdfd892c28b027d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f3e191a0c7abf789e7eda32fa5f98c49f68;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c17f29c46da3fcf3ca11bfa74c106ed26b3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9d87f2876b3ae6f9ddaf53628c0b48aa7364;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h973fe2587180896f3e4ee56dd7d501209e3e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he7b61f5ac3b2cf0727c22b27debe409c958a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfde0d2976eadbead87af4cd64269b51951b6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h80b5a10c1504c41b957ff43d9cece5aa2668;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8490be26597c0d9469cc6ecdd501019c5312;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3547597dac4b86964ef4948b26c2aa370634;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h10b035e7a541a18f499aab11efb36b1e2c1e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf32bbec5652a98b4c12265beb2575cdfa450;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'he9fc3d2ebe04cb9c264189ee8b2c14157d90;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hc7ed923c21b37c11c2373fff29ae0fb7794b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h491e27191725910f644bad387fb640894e7b;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h797560bd343033e14748e8a629d32a98981e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3f7b97978c17bd9968e9749b65004b338fac;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbce9afc6457a3df3d8897841cbd697ebdde8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h47944716ea4820702834289aca41c287f3fc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7daeaf0d0475f86088805ff9691f96c19940;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h256c5c70f74642153b1725cdf71308cdae64;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hace4242b8c300ac1092553f3846f8f21796;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h77a89f5f40c0a94af6fcd0bae230b29addf1;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3358424b97c2ef9d786606e74d89444db89c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h34ef39a792eca83c357652180fdc434553ae;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7c6aae65b03f38434636572e0ea79d625d30;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4f0ecdc6d48860d8e478504fc9f109a0a231;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h416f7505823a499b1d30edfa6d708198d09c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h27cdf52ec7c24738b9bd514fef00292b80bc;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9721d7ebc1794daf69a73882de641346774d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf392a4e5fefacd1ed1ebaee944429633184a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbaeecb9b5011c928e044881894c146ab47e4;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h835445aa8f8c921c44de04fb38674fb464d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h245a862d73ba6bceb58a59bf434da8173306;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8ffd89cac69279790cb2d3662fd187756538;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbf7b0aa2ba860a5a1ac890cf277b07a5df09;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcb7b786ba47e39600cab50e8db9c19f1e01e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94c77ea46f576c97b7e594d0467af47d046f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h26950318fb7202766b4785126865ab7c7e93;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd634760a609220c455f89d7213a0ea344ab0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h31d25ee5d6e43847b365e0af6442835337d3;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hbe4a07657d331fd932767ecc652f980bce85;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hacabf385afb9cfa8a14c4dfaab02f927c0cf;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h9e85b959271c8b34fda438ab84d71cb7d3ad;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3513f97b8ed2646bbb0525ed111a7ce2a825;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h75d61689da798ee1754a7e62f0e1aaf9c852;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h361cd9a1882041df8954e9899b474f7a6d5a;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haf175a2dceaabc45b3723f190aefd1d3c1d2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h73db5806a607cdb10e089979a4b75add1965;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h2cb9a26fc2f32308c663d5b3cd5ba13568d8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haced6e116e85743e0dbe73a2ff3657a518db;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6fa184bfee4dd21ea2dd7582749e73e96fa6;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h7d7fa9ebe28b2d829a0ff7368c16cedb747c;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7862fc4b24c3506b9fd5b282ebf448677a7;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4702211d86f7fd6d53480e3daf2b45ee4c72;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb431d3a32df206c4f26dc4f726c2f02ac6a2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf9ee791e2650d746456ea49da59004cdbe0e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h82899b31c195c33af366fd66a453a8e7ab28;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb16f30a0c181ced255efb803d3a348049d0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h13ad6cee90a8a8f62a0ae526beec25707b19;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf3271f93e7564257e0e2815221402d8ca3c5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hca1dcf972b88166ac6a36201398da8643e25;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha166d2dc51e4915fd26e691cfeb7e5acff98;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h35f9dad2323a6ac52e098a4035c4c558bfd8;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha271492296d44032f43b6f7fdcf13f9b9063;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfeeec428d8075cfb4daf4291848ee3d12e1e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h485df55a6997587e3420ef86d8b635a89021;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hfa274efa390c14fe01f4afc3054f8382b57;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb3ccff520b07279bb2f0b80d10aa663aa30e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h99e89854027cb9b93c16f97b019bf380ff05;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8a230f71ed93d5543ad04dfac183f0517da5;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb316cf025b4bb8593b728ae785f1ed672427;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haefbb53f87c7009b9ec34e38428c59e83199;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb82828302e95d073c2c30d234093715f9cb0;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6dcfba6f25ff7cc6ec7c5cf85c75b188f939;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h1d0d327a9f881e0af8f54930f141c728baf9;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h70a84188bce9cbf1616bc4bf703254586e5f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h94d8aea03a0091bd7714f485231272c43f6f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h59e47cc483db917a2f44eb3ad11667e456de;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h6f3024886c579ce7e256698fcb4f8f984d19;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8adc4ee2667cbb1af085ee982ee13e6cbd18;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h4bdd21d0620c633104b817f1c86ca87d012d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h3b70ff21f53b1789007a428e3699222e0a3e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'heaffddca9bbaa1752dcd0b54a7b12fb8472f;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hf9d83ce9164cb45708a09a460ffba6a82601;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha1be5f3c72fd64b0938a7389e2f514941751;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb517f217373644a189f635034ee341cc5f20;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'ha7e47637feaa6d33fc22207773c2c399278;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hcca3e118d5ee026d1b825e9a1e35a092f2ef;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hb920b0911de0bd938ea9b7959e2ee44a9f00;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd07ae4b8c28c659ba74297f93859beccaf2;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h8826ccf9f5cda5c8fe22a40a52518e8d0b40;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h42d3fab5f370126e4e5dbf24a69ad9dd7a69;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h44d686956e0464ea0be3c4050c7c36d7ae4e;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'hd7053d73580456418fd855b4b6fc94fa9d75;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'h53c7fa1df4e6308f6d2909e12c5c5a07f34d;
        #1
        {src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 144'haa6feb3ff42331a067a72c317d74b205307c;
        #1
        $finish();
    end
endmodule
