module testbench();
    reg [20:0] src0;
    reg [20:0] src1;
    reg [20:0] src2;
    reg [20:0] src3;
    reg [20:0] src4;
    reg [20:0] src5;
    reg [20:0] src6;
    reg [20:0] src7;
    reg [20:0] src8;
    reg [20:0] src9;
    reg [20:0] src10;
    reg [20:0] src11;
    reg [20:0] src12;
    reg [20:0] src13;
    reg [20:0] src14;
    reg [20:0] src15;
    reg [20:0] src16;
    reg [20:0] src17;
    reg [20:0] src18;
    reg [20:0] src19;
    reg [20:0] src20;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [25:0] srcsum;
    wire [25:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h920256b86b792ed8356732f02a0f3549023e4c3fc5b1e6dab411e1c70def21c41a57a3c335fbc5f98c823eb9c6aadf333a08a1f80300f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12f3ce8df20640eafa5f8d3274831dec4d132d3fa6b5a0f66745d786585681a60739bf988507e743510c07af649d77fb3fdcf592ff5ae93;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdb01a216fb6c34e13c4ded17d5a5cf97fac73975ff13dbb3a3882cbededf2c3a0372e15eb87a40d4e82625a26085929d11d6c8e9974727;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'habbe5fb218e478ef96aad853fb0923f1b200e3b922cb551cf86d33f0e627ff9d59d9095294e6be6b888b2ac37965d4ec9be9de5238eceb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fe181b230b348c38d5d38b0b68a6b4f9023e49edcda69b43ab8fb43cf7c703b117e8dabf159c1a800348a82776a0bc428fb00c9fe076a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9ddf5883b6a48e20d9ffc7c25889f6c416e57c468bf8bb9ac0d724f4b57ba05dc8f0c4f2d00705cc21b52ef629610d2fa3a55ef527f9e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10877cca3f4d8b7207885ae487bfa47308bdfa36ad59749212f56a8568bd5a02fe10e3ab38418589599aecd9c34fb76f01587145b8104ca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18d503e77f936e3a501d0fec2ca5fc56f22306f0a5cb7af44c09c39bb1fcd07fb02046fe2e9b7c5f7d07aa48e3bcbb5fd666e0263e43592;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc7388ff1deb17e7ef42b3d7de29c001f72b38f2bcc945022f95e32480530f94e5722902be7d835476f95686e462e21516be899f130a10a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2bca066a32c34111e6384a1d48d24b50fbedf1eda03750b0ddafa77b7e13389a99137795ed86222dbd002cecbf21fa6d2c387938eaff3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17e9b6555f835dea7aedbc10f3b437a6062a4a1effeb0dd1396662c4b036a5df69c4522f442252dad9f026bff177f9c81cbaabd4794a424;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1298b34e5248f837110fcacb0c7a94e1e8fcd3b0cd92318158c131df6ec048ab70385ccfbd9a9ce51614bce8b0deac7aa0fb22c989551ab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4c699a99df3872080cc00258a686fdd8a2cf110217af7f0aff6872ea2cbe51a745bf1dfd16a96038b42468838affa68613252732a24fa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c5fc6db9a7c903c384a593040028147ed8a3117fd56fe4623649866f52ab5f6e7b9731ca47e777b5eb79c352d7f622fbc55b90d76b6dea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4acc1a2d78f48df3f3d744406d773e26aecabe95ea54237579270973857b49022aed28d9a5162806cf2bf36bee8249ab4c40621bcfafe8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11b9c70aa8663bd5b24603b418ed544cff8a23d47120fcdd4661134d0990b75ad3265226fa63206ecb182ae7d72ea32d93fd6b70ca31251;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h109480997d3448ce2b7ffda8c8e54eb950c1da08e09365491bea29d6205eeccfd62a4088cb62bcb3da3c63163f56b08294e6ab32ff60d30;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2a8743197cf5aa9937e09defa7c9577beb5bb75dbebc185fc7f8ff045c36adc0d6bb75a05af771408ab0d49c1cc449f8303b36e7968029;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2152493adc6a252325a3c263ff6b8d03774f829d3d76294428570b6dc94bd2c4929cc711970bd7b03ba7e5ae2fa7e5d21111e363213979;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h67d25f07df87440bb38bf2a66218c8cd45b49deb87a46366f4c6eb456e4d0fd9d11efeb54e05d2ca27ab9d795bb4838628fc3b32729d46;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15f5d7c4b1064a31a29ee35a7966e0c6962751411eee0f219adf22eb7a7b07472d8ecc1e72145249568b674df7deca68f0d943dbac8a4a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1be3599e68d3507414917b6ed92321d3c45405547ee3e920f4548f66e5350d71579d2b870db80b41e28b016ae585c274f65d47de3adb89;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7c11c586aaf02ea6d29c8bd165d4ed1e5d1e63e0f70456ae3b2dc07361e53c5e68f0c53701289c72db6661dbc02a197b61e3ad5cdafed2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1232295bbc05f9103b863bc3d7977ade2b225c897282781a46eddc2ba90dfc298eb6be41f7d125de39cbdb9da6568b0f6f43e448a5c4e0e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb6a6ee881adb01ffdd3e634e88429badbf2710a8f12920721b9ebd585bb08ddf93d647d61984f68e9647c573a8b212e1cdc07142ded0f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd96a0416b7d776511da0e3f59ff553c4bdc4a3b626c431aecd66e9a7fa06265fe576d346ac353c15f3ae3bb57f5761ddb68e5533cd47f8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h240639d9907f08ada031923dde8e3949641f1b9908cfda80ba6c05f9d735bd825dbf6be5d2d3a82d87cea4773d90f5c94218ec140c7b85;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h520d79f768fee79689c1a286e6a2f8290e2bfcdbc0f13f18dce23893b13d1d7ae3e5f2582b67fcbc3a75b04273ab839af81cd34c2ca790;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc9f8de84aad7737d686550ccef3bd58532edd1b370f9d32f8bb4badc360715f238f1851a50c2274c24ede4e24952823263473d92fba66a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h39f66f3f1197aee4362f0b54b727d6ff1d5cdf98870e9ecb795f2d9dcb7fddaa2e8122b6cd322a9080e93638115b0b36896fcd39187fdf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h270d5db14645df76055aee0ed1321a65ba92945c6a60852c16f99498d2da1357880c9174f23b9562f74f0645514a065e7453a971535445;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b1a8f372504a43f1daf2dccb3b717ed3d174adbf4d92cf418d1cbcedc31fad1e5137572a19380d4c34fbba95efecb910fbe2952f44fea4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6f127982efc08d6f85ffecf4df20a9abfea5c36707103fde65d8af84a2d19f66b420c387ae4dc1a4e75fefcf32d47dc312594203517d26;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2521bb0c959ea57f358ba4c6e85333030d6483b8b63d101ef65ca05d3f6b8770698a023caf194e81aef55dc56dd11b5a46990d5e7a3dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8cfdb14248617a24c5060f0ef0303b44217372dd0124d0a9eca7b0396f23a9b05dc6f77f05acb1d97eb9a9ff24f69af708032d2f7dca17;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fa84379a7a39a3ee0e44f27c8b1b671335c8257192f99b97bb17cf961d88eca52895a841536f5d54f9b6d6373d312dfca8657c26e6fd64;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h49b878346dd35a406c2cd31617edeb6e4a572c41d00238e5ec40448521b437b50c446914946793a9f11b91a573b4a9f75d0abc4989b35e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1545daae875f432450ab425dd59a2a504d89d0ac7f533ed2d3eccac60c7698c56050817df4c69f4c8bfa8a7c37c54c4fb158241567bc326;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf33d15dd6502c3747622a2f8a2ea7d22dac3b6dfd0f73479806425032990f78cb46117284353de731690c7657c963f1e35c1512ba726bf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2937e97839c212fa934fa0c477a449b140b0359af66d50baaf00eca7a95499af1f65a570a1e533878c0196af70044d00802fdbbafa5f91;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15eb57a0aa7e9639da4b5dbd67db1fc1cc1b53b2ad6dc1b5bc6f13c22cc6c2f54ab3497232fd5ecbef78e69bdb766148501eb54c2117e39;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h39320951b67068879bd82d4ef061a4cbdd1cd0dbb6b28f795d44ce4ff2dbd111732db0e7819673aba500c2754baa220e605a0b22ddb18e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a52721e5ccfd981f8b9d4fc45052f19980c90ea27d54cb1d25137c8d8dcb06158bcea39558d13ca863b88e3dd4b8643853c9f571972e24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f23df97e3e7325bbd5d449717aa74345433eb0f1f5f83a38b885c2ad889aeb3c99542f8bed09bbf922ac235c837da358cf12c34af27fd8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a13b0b9ee1bc543e4e54598462fb73a7dd05dabd50752915ba992df816b0230d812552e5013750bfc442cdbccf70baa5fcf41901bbe2e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1adf77ece89a9f13b70cb62c7ac5ea3050d66ca760556a47e359911c1aa055743c1950221acce10e96b9ea09e264b7dc9158cead424186c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11deef310a5df2dcc2c744fe6ac0ffd87aec8a1ae04e4e10f5ae6bf3f9d4220acdc48abbb54ddb145780f5c9e82ef02a73ef8f98a4aa648;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd8585fc26897a8b0c0a62abb24617920c4f9f84d86016bdb0d0b9efdd22722969e17755e5bdda79225c43377ab3fd7cdf20a46d7dd58a8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f10e2e14957fbe926c17c869146ecf5710d7afa972c5a859ed423bff035ddc21204b1a6d2ae2b4bb40ef6e7653c3c3c3afc18e394587a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b608afda9396549f6e9314e5afa72229d1cbc35890f62ec5fcc15182642a6be0bac617168285e92ce83521504f42887a4b3dd1066eea3f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9b3dd996f6cc964596d6e184b3866671bf4502bf01089350b8142ec0b88fa4542814ee4873f41c4e0f36958021a8dc6d4b066ba650f7a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a5b013d349d3ef8dbd2ca4fd1842e8785eb190cc0335b7b85579d965182bb0b7e5dd5f6e2122fddfe1322253d870b95b1dd96b1477c155;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1acc43b00d412081cd989a7d437efa9bc9ed0ef3de14b75921107a78873c9c3d06895650fea9177470ecc82dc9a07e49604d5dbfeb5c8a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18fb0f131e84173647f9788ed96d3a959442c55020126ede22db3afb2cde688a4ae3f457513f4d202c1a9742ab692d8380df6c3a2efae61;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h513ddeface43416113575e0f39233a2b8e29d56f9ef30fa0743a6255f0a870f8844dbe2637b2113ad107724d2ddc9d00fd6313bc3550a8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f12e1a9022cb31c12ed57ff241180190d3f863a3a532e103e15391172bfd31502cbda52edb964c53dd6464c9f2a5794662bd1ea0d9216;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffe9bdd277dd6dd528a2f8a3fafa9178261636c5e6d055b3e5762c323894df9ce3cbe98fd8edef19ddfd757ecf1bc0b2ae2df60df06fe9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16d392f77929f7829a471ebc8ede76ba757d2a14590f67de4cd56c9509dd42c56b56da31d1bc73aeac1d87547e421168c8d55642474680;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a827c0ea98e8f3a9bc664cd5ef859042e7e4d6efe899a2e269fcf58e623ca6155c2e0baeef25db82ca94ccac430e9b38588a96164b7902;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10320dbfdeaf8d9f6e65086b66edcf614262d8b8d8f9619d1b212f3a86a41d0160b26240ac3ad1c499cd45a4eacb6bfa0fcac8141830944;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8cbd57908749c41d606cacac452a1fcbaab058767311de6950c17e57e5976f84512829bffea05ae24328e5ddfc0a403c3bba743d3337ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h763f58865520908a533d43548096874f9b10a7566284243240e18b724dfd6deb8aecd16ccc058893dedcec1a0efdd23285cb3fce919d80;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h108ab41850eaf4f89efc60c2b11d697c0dddb4ee4ddd222a5c98b5cffa0af98f2e6b3fa9bdd211454f84554bbb974cdc22752f8ef0bafa4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b39e7b11d3bca3b026db4fd5f6d6ee726cf617e560936af43ad2ab53ca74606f22a806d3b4d7c5aaa6031a8a66d7d060e302461e3bfd9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'had78a7121d0a43e65466817c717f259e40f8776b4e9468bb4bbbffa3c32a3850f8d26c5baf98b2d770580b226311c8d6a4653e401d993c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h155039aff3437a2b9be9a805e781f1b99aea8aa9b0d23d249521b2c94fe746a1c216b810dcfc0191b473490d11b0b0a4ef5e307c4df5d89;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b07e90b01dfa44fdf1a68fc7e5513a6334b9fd0a1241a72520d57a60b4b7e7ad7ab5c8eb8ab8f66d42a2dfb172afff63713e2eb8e47232;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd67ec78c85f6ca0d1c29f9bea6df3f59425927141c382c7d9b503933fd2550b2ccc7fcaa01f82d79156dd8d82ded095de1d95e387f88ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h23b9c00920d0da426560df72cc07c5d8e8d4232307502494d81ce0730b036dc008024f4f5803c3ad200649df837a8aefb264ffe13c2402;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a56640d6a12c733bc81832e38224e79da766b630f3bce02f616773ea8550f08979b35d5b0c8b211b8e3174cb6bf5a570b993b0a850ef25;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h163b9aa02d6cde53a08117225a7ecef7c276cbb08fc080dc6044835da662545b41c10095dc684ee6e8556c813228ef80e223819e9e1e126;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11ee86fac6a374c26613db6e3f055d803baae73563ce13b6533c4a9a182e7d7f641ad4824a07185ad54d702b32efd411abbfdb12ff73b74;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e14525ff5adf233369e9641a6102137634f7c541076c39a434ec1b4cfba3a0748d82e8ea68ea3e6272a9a52e25ac7d0eaa9339d02be8e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8b679901c81b67868eb3890b6902c3fbf0234aaa089289eca0f46e4f15d576e5de554b9f13a5ddbee951b9f9d4bc4056d966941e34bef0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140f0dfa0c10f5ce73bf0c444bdb8e158cc0193c9f8a8e1b6bbc1a92dde48e6eba28980dfd635fbb869c9cad7a6a553e77d432807599538;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1380cb92005d668ec31cb1ef5c279c30cfdde8f9d1bab7a419720e78dd834758ceb8475e16184f2e05aaf519520be37802eacc8212335b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h197921756a621ef5fc0c2b6cb2f75f271c5eda4498a2fe1060439c330a132b0ed5e493a2be76d871b4ec2cc8d3cb27855e33a2952c550f0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h178d88de62d787073cb814e0ed5a1b5c376b0d67b6c0a7064fcbc3889f74f7b68859c8717d4212eade8241cc676205efd173833260b8361;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10e62cbca9be5de2ecb98aeb0129a10678446fd78dac18dbc2f8022ff88ecd560a473591eb52194938edfe07560ae329901760dd5fef2cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6b86d7e849e7867fa95fb9f880f5f9facd2646615e757e9b45183e3ce9a5c834659dce9b7ba59fd13277994ade018b5efc86ae66b84415;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h31e6755f988e01be5fe50adbf7803c25a7967e6914e66c788bd0042e406a29c6d432a68ebe16efbf41e1728282a0ebf56a6acc65def5fd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fe9fc31ecd051df31a841dec83c5f49330c3c58759e2c843d0321eb9f0afe200c86fdc96629277b45398212fdbe214123e7fdbcd481eca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdb3bb73e9cd9787e736d760f88738ea5c53ff90f7c1a29a90a4f35aeb9fecbf67da933f9634793eab4dd1c4c1002a18af8ebef39d9cbea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb01140c4f2eeaf03174c9a78e2915ffaf31d93d206841d2deeddaffb27ba515c2def56c99154af29c8fe2f2f55ce7bd170ba26d85129fc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2f5899437295ec3af897bc4e25720a567f5fe6ea3adae0c9223b1d4d0ec894b003b3aaa241b848157185b0e33488c8edb672c36d0854b7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h82f2519f781d3eb9828b809e81e04a311c1310329d6975e565e565de240d83437beecd8f47f0514f2b408ae3f63faf2c6509ab2ae204b6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf84277e32260030282849a2cf3f54746830342ebefc49c0d481a580ab50c37453eaa204a97d55697b1cc4a9f6482fa24e4cb6490123f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bcbf90ffc3dcb66fec632c3ac702d6fb6e483295bb771514c36f7dbd15a971554bb2f32e2a6676153f13f097978f5da4c756ea75d46be5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1969f9a21acc610f4f716b09caf1799b9f3e2265073add3c6f6274ab3e0228141a19ef5571f063dfde9fdc8f2fc8a0070206e72afeceefb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc9acd138beaa608d02a7b9f6243499a2766db9107c42b140ba1dc0cfa998a3bea4fe85954032f2efb05cd9eb620b77fd46f224d30b2ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6bde5c0e5a23039c749f3e60e9cb1b2aa6b748f310902eaf19c50a4eddea8043c2c6965c9dac94ece2f106506ae7e560f2bd0b3accc969;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e1678ccabf948c8ecb7a6a7d7272677711b34925110807a2c8692dab04105022f3420380eb8d8155782594c7a7d6d6ce304c852e5c06;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d94561e03f925b35707b33a945e22750a9b3fe0b33e2a7a3701057c03930aaed61471c949b7ff8f9dd2f14d5fe61344e5742221356a369;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e242e298e4e875973380c1c037aa89443b3ac81821fe1300118e5f64aa077a9d2259cc1fd0dcd7a03c1bf350f7c99dd0ea56823fd706c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he7352305d0b66225415af3d34fb6e4d07c906a4b704e807f4bc28a44d95e3c19b599bfb099527e2fc355c52e8e7a5e60d5fd7e29742f7d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8b8ab93319c6c441a54d2a6c01b9f589df9226d3817f8373fb4112aefe9257444ac6ed7450c5985e8fa311435efb497131037b125b811a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7d348195c4490f37c88b5224df18e03408e2a6403ac4532686b4fcf74b00449b1573c5700a67e5124f027fa5749084937a2508f7105880;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h148a4d4b25d1c5e3c3e3d657cb6958c6d614ff627fa4a625ea3bdbae2fb19177c4a870280fd2c1c34513d8ebc16d9483d6255f4e4cea606;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3fb0d8f40e3d65ee374044bead799e44da5fc7efd30b8d0a08e6e1c9b91c53174c19620b3234c5d7dbebc2c66a49327d20532091626d2e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf56575ae454bb2e1849954927ef147133688505b3aaaf2517345c1131d35e8e78980e246aede32c7e638474eb280a9b1234cc319417e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a92d4d5e7e83e7209c0fb4b0ef6c8929ec7a2bb4315aabd6c66896a49955680777c288575afd3a6b6e9cc010cfec920148eb81e9e9f528;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cd13e8e5b40bbbf61f3db42bd5cdb885277aa9379cc29d39a2d15017e5a9f52037a2c29154d87355d00b19cd89dbdf00804a5d0b1c6d44;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hda2ff1f1b7b5cc1e54dc1288cd960bc04d1e3c3d68f2367df726a25cda34504423a0f1a80fd4b7c415f7722315fde9f04ede194e710375;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fdbdab0df89891b869a1a254fc9654b295eec78ef3625540c966929a7b362e06147bdb5fdb1cd744f02e898cb42913ee45078fa05c3cdb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c15290a436a3e0e6eda74690f383f945658963174d1e98a7b8d18554cc4bbb18c8e1688a7d62e95bd9975757ab220c94a364b78d64f8ad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb7f633914aa37a84bbe45fd37ed307c8e8d54c35df568a543039414c8978807b2c756067b3b52ed644d5e4229c7cdf9e239a53d13603b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7b36f18814b59acbf8751879591cd7c318a6469cb5591c4d8b70558f446f61cb641b1156fa4cf4683cb9183046f36e08fbaad21b291374;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he917eb781e8c89d22c58546a638aceb60e0ad8d4e9c448abd1f46ff5d48e3379b7b93c886f24f0f9b59e0e8da1f791525b47c4ddd38b70;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2d6d3e0a2f8e30fb4134c7deb3c793c826dbe565898811b8153a6c6bea6b213f9841020467c3b03d2c1b3a87719a1d50e0e7df9f004704;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9597aa96e21a78bbda71edd136a4b9b3bb8310d044ec10ef5f6ccc22c6949cb342285dbe079eb0a6fe110a99730cb07a444e9781c3e855;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e2ec3663aa435e4abe3baaba44350f6fb0013ae91b860744cee47758c836bc98766b92d0b3af9e32b530072b12613fcfecd7e337625543;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140cca9305fba89a70bb200234b1f394b45379d0171daa2ce879dc305b24c96a7277c71bdf22e9fbea399016f63298110e4ef002b416ffb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha1fa6aac9ea409bfd3baea2c60d9d0994d737ef5c94bb01f53ce02bf47edecc296de52fdbafad3f513bb13394b2a2395acd0def40ac7e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h342419c94cb2be980f322cf58101149db5117d0e954157e8ffe762a279c58f8b32a79f2682f5f1c7d216a5f63e1ba9185514a66f02c913;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dfad8df2bb050c9c1fc1d94e3580cbed7b6d0be12521d373cc7b67e7eaa725c3062e37ad40f7a5240f3b98955de8c2fa20d256fd6ec7b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3bd52a40558dd79d7b9fd3cede77ad926a637ab9dac6381d740e232807fb277f606c2bfa118713a3e3e0c51f6cb0a8849bf82891a43996;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h67cc6d23836db72f8b93ea5aec67d40779adea93b5ce8b79ed1f3eeb1a95d0d21e7cdac82eab2f041fcaae87d995e43b9aab586b5f1712;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e7aa73df961e787ac3eaf9de7f5b43947825772898d03d7f20a7c81f60dacc7c5f9cf49de8075c438f4463aa934a0aacdc4595736c4aaf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16fa6d7c9aeb58ab32e55117554907b91f734ff1b3d9aa9eddd2f812c3aae8c7316dc367371d9476da085216783e744fa84f734a92ed183;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf3c7cb61adb98f0b3ae825ef49937619dfe883cb1dad3c7c202a32637c0be48cc4b34f0b1c9a701c156fa3a2e4baa0f534b43a509db64b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb18858217514e487865176c58dcfb3e2dafb2e916739625b1535bb8114f308496ecc7fb8a9f4c45a5a50586c82d586ec7ff36a2169068d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a8294790de814522513bdcf07f608e0a61b76967f611404cc02487ea5ebc11ba7f64282d063d922aa53f45c527a7dcaa5ec91b543a8fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11543c5ddde620de67471a0b8075542421aeb72bb51d9e9d31dd41e6b317f7eef06e4459e114ca7d6c17585c24775e432b96df42b236903;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5db743ebbb6b3c375ddf2830b25ff3d6904764387bddccd031964e1f736f10cc92ea18b7ccef8e56b250117e7103491abd7c708f2d25a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hefd246fb37fd51631c761088f68dea40653aa787e0f7b7386b264cab3a5c9d422c6412e8692a2d256266599fc9c351a1d560df95cf2e2b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8e3fe11b274aefea77181e66e2634dbe1ade1f8ba38f437ff49e89423734cf77c67bf642cb9ee3340a10ad24162d905fcb7c5885481ee6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c21d2c8278c278abc9de669eae6e848b89b05a1ab2235035530d7c8445c13a73c9e7863e0f6ede85061faaf0bcceb2ccc52255bc997ae0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fdf6f16d1b97edb56f9ccdb30d1817d2ebdce6bb9a11c5d88a718a0f08eb7bb4e7b51e3472e2d1e3ccc8c0786a5bf020f4b2a946821251;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b1323a4613d03da3d925cec339244b6efafe71b98687677a7e5f13123c1201ea831807507dd9feae99b3834a28c0e2531f73e31ed0d61d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h885049deb1a55e91d81cd82330eab57ffe3ca1e5d6f1e1c4a6405206489714d03f717e1999f70acc122eb951f6631aa0ca555d9ea2d882;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17456d1032672f7f79f0551e6d5bd001b973f243954badb63d4611726ff5f60c9dd918c2efe392dd53b55135aed5c0ac8625763f3d2a076;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h409b38808f1db26ad9022f14009e90efab4acc1a450f44a44d173f5c514c582720855b313c810d1b9f74e97c49d5644752452d371116dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8e5ad684c76e41087b1464e8f2b46d93aea290893f7031e83056d0b27ad82eada8823fea3e5d24d07bd29302500654437da195ce724ea0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b0cc777d77207c886aa8a50e91ba5fe2fdff080762b96574afb2de35d66dc5f787c69635bd3047dfe43c3710fddcfe4b9c220519d0b3b6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha76f36744c45d82fb28725b8ce6186669acabce7375e734cb382e4c5097760059bf980aef2ca727e160c291a678b679768af64843785fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h193a78829164eb2d49a714bae8b3a9074d88422f32d3b75c7da48b02ce84ebbbed16c560d2c4b87e8e26203e615cf5b15f37e73dab179da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h60ff7bb5f9774320ce8eab309d6e091805bef78d48366f5235699039d5c4a8dcd21b933d40d5155a0ac1575049a1424d739a41aa5181fa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1680ab9008a1187ac6190b60845eee77cf12a306f601d46ce72524e901d0a3b03cefbeb948b2ed31dfaae2758641a945372cf4ccf2605fc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h155ac8e40ead6f3c0d8bf555a0b9d26087548804ccd1c3c406014c6ea34f389cf0ccd0c990c50eab8c1b8359a24a23bdf554d6a51137a20;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h110814beb1f1268857745083ade0f88c1e86d6511524db935fae84e8e9056f92e022a198a5c9aeaeef654fb5d91d065de264afbe53b205c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h32f0994627047ea384a384dc2152849379faebd5e2da7b0aacf1dec57ebee4d470c758a07bbbac361f445d470ae3b9c6a545f524fc98ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfaa19ba7f1d33e3d442e6b10da178ec83810ec4c6a4e8c1b2b6c85f86d78fe70cba2e48758c9edb03e55dbc9b54b245dee4834a030b334;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf318ac995143ce057ab9ca829bab23d3cbcaa61c1df701bc23ece9e609a86bf32595609653af44b042471cac953e8fbda562e337e8ac7b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12ab59b40f9b19b917d48150263bd8a805c0e747188eb262866a59a8a417a666ba5be93b044a40fd9f0aba5acdbdebea220024ec3138956;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11d098de3925d065c27702382ba9b836c8d2a956c90f7a850c82a15daa46a83cdfb3c9c1d56b06020f767a368d21902fc853714c1ad76eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cf634efd4c9f614dee387001212c5c6765f6ae2e34e367c53556bc7917832cc343c550becb35d26e3999c9e8d09046e033416bc8491aad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ab96744110ef791701b1ea37adc76f0696c839dd7838ffcb609871a0f3fd62cf3d37ccafbc469ba8e4ac40534dda0f778e8d6b827cfb21;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17d4d1b2b89a32a049114b73b16846b3c87e1569abc7ad085c2023929990314ac1ae8d5c78e5b274ba5ffcc2c52f03d0c5f4f5162d8c582;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf3cba0e55bf5a0d7aefcc958dd771c4cd88b8779e8e4227177287ce9409133228bab5e8dcba0ccc640a26be95de7db4e4a742b7f9d5b43;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1724371d0ebb662597f5b6eb6dd95040a2e3860153fbf620beae4eb97e750226c62188b9ba23d6f00f6bb3f382d17d243ab4e415fcc5465;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1380e5c4fd1b582826f2a21d1c2aecfa6a5f70f2cc13bc4340ed5743566dc1bde8722336449f518974ce8b10ef5d77258a49170af27edb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c59830744303e9df22e62ad0e4cf638f9c21640d570a2cafa1fe4e9838570709487da0f1a8f1dd447d488e93415d3483cd5f5c210f9d12;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16f6f569b25cc2f8d5c092d649f7e54b8cc8278e8f4993c663fa8b3018855fcea453c7f83d1930f39f4adc0bd71abbe292dafe3d3b91202;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1726d5a63d4aadfd89ca2ee2c228b730f77426e653483715fb3e1aa59db5c364b0f920607d48034522ed571b5e1f2752a4de65684d750d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he78ffa42af070f578697f4a1dd1541869900b36c099fb5b5cc6d20b00735aef599ed281f1a0407344a21d6791d31a8244f7231c5b6ef1c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8aaebd1b9c4afc3b23e0d38ec6b4ac67ded5d27a65d1686ed2d6c781f450cc086f747608b91611536fe2657240d42f0c545da3941d4007;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h63b61b0d2f50c991e655602399fb96ed6ebc71ef6ee8d70c66dcc3d9232d3c672523802b1ab228883cdb67658f141164428e00a28e3c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f8a549d8b6890e5a805c1363321cdf2cc67e1953e4d4a56c7c7e96a4536f6f2f16cc0f4461deddb735d98b9bb0dcaeab7fa134ad99796a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13d62061d173aa603b68b014eaa4e6ca731d580b91fe893a052e36f18d23dcdd6773e43caf07cd3fd4183287d75779c1e35afa234d83582;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h415e7f727d261e74cfceb753a47b19fe2a493f1fac8d3474daa5b0e7fe185ced9ca1493faf3dfcde7bcc3ba2ac3821c38dc4d8c7096f8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4bee070516f5f8f220a32532c81ded4f9d72bc1aa3e6a7dc247350091c330d15fd5067107938eb5b16869cdfaddd43779d17e312f81c1b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ef8aa40810e9ed73544aa2b76660e8ca1950faccc51753be310e852276b500e8e4894c62d28c96a497cc3814c701b7f7eb0b01b24463a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a71bd66c6fda0a6c81a71fb027c4a5fc1cf78515cc36710b5b3e8744902d264ef8d6e214316bd9fa509c458f96db996c8ad4a2dea8620b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h174e805315506f445cdc3ed62e25e8d410bc19b8e94a676b86d955dffcda23188ae5b0cf13e359c27ca2381d067b76c6234ceb0177d6c3d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14e86fdebc32b37d0ceaa4dfc059d849c2c7181770aea0f15aee1fa8481191425b0beeab67431f3717c51ef278623740a9c7fba1943271f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a7b05f5e10eacfc4c7c41016e0e81a73a3b61c5c8f16ca5c42d41ad583442e829ce8b5435304ac18c88344d0e674d6d7639095ae52c6a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfe04580dadddec4ca38e4045655b1b39baa6689129d210fd03aa77781289d3dcfa05684962b4d98bccfc5332aa85c070a2ae6b7e968e33;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h372750efd62470c3ef43bcc58784035c81eb19d22a659d7891d2347dee6ce0832311b7137f0272c6e30c2d18260402ff008192549a03c8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cacf3ae1b4e9fb7741125d491a2e77317b7351f403fa09901fd8a0e7c6290fcf60030deb3013aced42e73e55a9ee0f31c2179fb8ca1a65;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1866e658916769d45e73700427f73960d3c4f80499254dc762f901683ac1f41f3a371b9f0ddaeb655a618755d431aa3a274fe927fa3e70b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10e58daa95c59be692da5ff08305fd53936c81220a8cbc734d591e06d2abbc4363b652aae939c1ae3f8d0d374b436898350ce1a46da8d51;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h181b79ea8fc9c142c467e6fb2812bfd2f9ab8aa6a1ef2eadc8c3166918b2eca8a95be1e2e9ead75e03062cf67782f034c5cd66a299a0055;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15d61214612082401b1f687b21fd9e2c6dc563acdcd110d197d5d7321d1c8d5736bf69236867407841acd4f06ba6a5ee649fefed3cfe9b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19da758c1fe9270ba2039f6490753cb7d201f622ccf3c9b3acb2f81b86f710e712f2cf95cfc726a42013f46f59d35a9944ca1a85728aa54;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h193035b491a447e94f529af593d1b1d5c33c5b603e9831279730a1380ece4fa517a678c7f200cd17a5bcb2a61d0a6fc03b49bc796a18164;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h76a0f825c10858f99b9271e4bdc16535cc6d45213c8fdfb7e2047cc1ae0ff2cd2b498231fa1daedd9c8a8b776250b1919b8a8530fec9f0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b6bad50acdf5079dcb7200efaf50d1222df37f4a77c9ef2964cb1a6a7a1bd9b9a330bcc6b9ac35eedf6229b0cea81e96a4e5ed664cebec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3aa27c3353f0ce2f6db6b0b5e7e60b35e5553d49db8cae451d8206495893c18e265d76006c137d76a059c06c19da8df881ef8cb8365492;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19003fd53809a140074ce464e86afd6c3fe0391da08422ed2589263c6a366aa3f74b498c8eeac21148287c6e49c4545d3092d6db8a2e94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h73d918f5093d59016e10dc47a60b45ea2f4f4de88737faa17641d595f157a6ea72a47237c09cb6734f9119ff724f4b9eace7f5ee24a537;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10928fb320d461bdcc0f1246ef71fb1d49594de04c84656769cb6909346a095c6eac2010645f10de9c487bc85d04a9861e7636bf4940bdf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e7cd6c4a4efbec4efa136ca2db95dc6230011992280613317f1a5422f2a9f8742e2d758661d7a3b890802490ebcca79521b991c4a8d771;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h22e5863401c82fec4f02b190c45527d683be9461ab08f42d09fe50c4c89ee6951d5938445a161fedee675709dddcab23355a7b9e74e82a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2e6f643711db5abf21ebfcfcb2b8c4ce173b29c4305f0dd8e6aef2b46f3bbbe55f63f9cc145d40ce7b07674d9cd1bcfbe77a866dd86f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h367a404f5026b11fd205040d4ed6679020a76b9483ccff74b115c4242a6edaa0f1e19de9a46755236e1042ca58c40683e4dc66a77e2bdd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1214f98fcf0981afd439cc73aa3066717a8ed246dcfa50a9d8b3d0331b8978c6bc350782733315a1d3e69a98a4202fe247f5db865cd0d8c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bdadbba4020b16d8d96b0d8417725fa552e16ffd9d9d1bf2b8593704f0b5b531ca2bb7b25899925d007f95f8fd4aa9b087fb4a2c28e18d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h179d33034e4c639aa21f69da7fb401b0a36cf71238ef5b7c3ad1eb48060e75623a3222b183280c9f837ef6ab7714f94bca9ec98ac6b7112;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc72f0369703bd92bd7c7a2644c252cacb7f5ae66676cc10279490d64b456aff43344d2d64dc00a6c7f91c6c1caf9396be1d23798224c1b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h46ad9c031612aec48c4ec80caf1b403f60b65a57a4e52d9239c2ec8c8e9cc85dd9c867296ec393a62db094ce7c655f6a8ff5da46516a6b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17bf4ad4f525f6ab8611152c91f4f32f70446cce0944471f7a60c698f326a67367433a3eca50361a324ea2446701b8d6a001a82c1e25d65;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h381f25756273f062012994b80649e532768b8200d78e4cd411f0391b55b04f98b0dcc59ebdc06302bde64fa3d2b978b19686b7ff45d609;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h122ef397a18826619afa455acfc36c5cace4600dd1654c4d3491a021d30bfc5daae39e87b92fde6ac9a169f205b647c2193fd19b288285c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de90e337ee88552beb7d49cd2928a20fb5b37f9ed791e0199cda2347c21429fedf9c4f81d7d6446a1fa660bedd449ed0adbc72778fc36a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8f6432b733440fb86e52dacceab3e130a709d3e6fe582a9d2e8f55db242cd51eb37fe3e6708d191098ba448c22c4866731311826fd6fda;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h107827b5ef5a26603c21b39de808e204ffcef7b552ecd6abf53c1c3881bb4c2cd7721d24efc8632d69f7aa3e3ae9d276a9f654e932b3f63;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h155840abf2b8f70c39ab59c813f30ac7264fe2f49547127b60bc36bb7683ee19de0060d3224190b531500dec6d47b263f79e4d020322522;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h106f62c32ee9f51427cdd424ed9ddfb20d1edbbea149307b293ef127c40b04dd4467d68e81565e162a15344b5d1f4c0fe16f74cdd950e28;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h67fdb34650f84cd0772924bcc3c78f361801bbf25921c0606e13199087132a30f560501cd5a9b85a9e61c36681c5a5819cb81688b7549d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h48edafb4aece3983528a9e681918ae35ab2732f969baed2af1274ea358d29ba512f2f6d65ec0ca7b554656321927b8d51c6f3945f50c17;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a3e7a61533f32516d50509ea7b2ce8a09eea3191ec00bdb09cf201e781432ca8f858cd7cb49c37a33f453d47bfe4ec5534bbff2d50c039;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15aac46382709b7815e2f7ba7c156362376aba58d7db148929321d41009fe4a4a7734fef729e40c0bd5e69970409e65b464def6e51b7ba3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfe9e0f4d985c480d10fb4b20d512088aa0cbe88e80c0c2312f579e962e9549d2f43e00b2a8db71947a08a97d70a8899ebf914865f23935;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h479c0a278611ed17a7134caa43d4a2867fc2de4534d144ef5626e5ca8cb9e19b70c69cff8f96e28c984124587847dcb7d9693ac637a430;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h113dd0cb10359d60b286754eaca8f924a859ade891f8e898e061558e0ba2b115afcdd60adbb7323bd575434b0ad12b213b0517d8183d289;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h46787b5a03f6b0a24056cfd96677a668a2447bfc4f780fa5bae42ec8a86e63c29dfc673da51fb6b0c19ab39b26867c800efd3eef9cdee4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1149c3969d995b4e3e4466bd10a185631f93452dc950adaa3b0ac7a8aa28ab75ed61786ee15971d2f30fb49bb1d2952a2d6ae530a13649c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16100c2215473112120048d5e7b920b5e152c9e679b04fed91a5cbb90788c9ae5e74c59f75e46b15e55a2bd2d863c20dbe7a7a77887bd11;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h99563583fc4e7968b6883ca28dfe899ca902ae345d046b825c7745632ee032a28af61c9215a0d696727f4e692be5da7c37556f0c36e681;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c9b5c385753f380396be6481bd8c0c73db70d33d14d8c67facdb13a7b872a2d418410d262153b4321e97c55f345634e1e109f34401ab5c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15cca02ce7b4d35d11219ed260fa635f535124448c05eb1d170624de89bedb5d5eec5f9a303f493dea06fd16e6b8d365d023a778ab6cd03;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd52d88f477f680115801d38de35e29be11d812f859727e967081dc22556a62c30d9d77d5da8ee5329abf30177f146bf57bbe4e197888dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ccb09bac19e4b97895016cf9e83e156442ae2b42d324297aa18b21fe448aa1330d977ad38151b85d532994b53c512e2df47c416f03f037;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f4c5f18f97a185f58bfad5733ea3514442a6a47ee1c6d61e5fd5530d27355122b5dc4ce212108112aee1e6b6eee4cee6aeb24642ec0692;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h182f3537488c8949373081ee6dd722469456ea3bc8810cb7c070a463509711653d8f30f2b7e10ec7cca1e0ad4d49ef854efbfd6f55b81ea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h45654f8068ba0ca1ebb04b3a3dd7a91aef0148d1630c979f65e293c1e3b0723a7edb96724a1e7c13d177df747889d086f190e54e1bc3a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb8661a809346ddcd8912fe26016f38ee32869621ee565ecc221068d1c7b29558c257e5cf29721aca8e9decb741cbf0581fcad42285b799;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc4f800cef0a95c02d0f517d58d7b8caa0bcdbcefbcf0b19d5af99c871bba054769cbff681bfdeb0c0e451fc0cdd7657021e6fb979a06f0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ec3eeef67c72d2ddac3b9577c41eb2de55313f4725434dd2bb728027f1248c6599d4eefbdb659a0b26fb6a7a50227db949e05743fa3436;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2a43143ee861c68dcd07704497915988386398487a46df39c7dccdd6da99b4b9053d5d9dd7bb639100a40032bfc06eeeac5f831e104cb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6fa69b678b6393fbf7fcdee3c90e4a3712a83de3aa343407a530085af0471a4d57a00c2a17afae22cc6d8d9768dd05d361d80d3627ef29;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14f8eed5103b4d7957acf9d071260d297470e1924d5b6061eadd4e52fdd1b4501fa776b54ce98d8cfdaaf51324ebc8d102c8fe4964c3d58;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5156e43077b5daa0a9c131277cc06e2671215b9bd66061e6afce7ec0883a782e0289d9dece83632a242684594e299a70f6262d908bd9e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ce32178754935716ca8ee7f6e2ca931844293a0e9b15d28cc06b66524e2b09847643d1888042a1d6c4df9b41f2e914d27c1896d9e365f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9a6187f41cd3165e461ee0fc9cf2010705f805c7e92f64c19bd50a105a2ef4eaaf7c648caf89041b8aceffea9ebf8466a3f2d8bf331a77;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1882403ec1a1cb8592cebcba2e99a587c129117be59eddee8601918a54511c49ce982c350b20608f162ba081f8ea87b5b21bf4e0319d03e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13857161f37645c5a9241999ea31e55cf5ccb145d65c811844514ea47f7e62186a7772fd2280adb7ab1c30a7dcab8af50529e1437510726;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6908a5b9ef8210ccf8f32efd04ef796bc44f97f779463d6cc26dee59b04f0cad6b35b89508aaff388b155120c66a0d18b34d96eb18668d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1003993aaf202be0657bd0a01eeffca1a51da71bd2f823ac85ffad8004b8915118eaf1e8a0f2381b54c88bf2e9cefa5f5bdf31fcdc0a24a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd296334636281dd75b4f5d53c6c04c6d8c856a01810a96bb4d31851c50690c3be97bbd1df3f442739d55d5be9189cf2f782ef8ba878628;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e99e86e74b4176aaae4ef270b51d529426da3eb45de781477ebc6c3d25b44b70ecb024f0857f49b0fc3b7802ab055ff095b56274d98600;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb2149fc9e7cd058cff91621c405c6d7c0b0661e582a8c35d4015bc6adcc4d43bf20f68eb6bb1db874ef802a00c46e8760e8901ba7eaa82;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10814795512b855993dde7d521f8bc2d8c61aa36cdffe2fe066ef445877c132a73a0c63b2b9511526db23acbf8f47c0480a92de8c344e1f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14565ba99e01ebe3464487d8815618539cf920ba805e3bcb3374bbefc06e69c8c093ac2c8a186b10c1261fa6f4d44dd224facc5501697f0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d5c7fc32f935fa5ecaf2660e1c59462d18b238241d09664e4603d063b2053e665553813db22720a199119b105235b4a29293c29c790452;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h116ed027e61cc8305d1e7ecd0473bc67a9059d3905ff1af17a73ef325380ea423ee60d3c8fd79a5d71256714ab80d80cd1a25ac1a7a07ad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19d33207e7a6b75429d15f10ce66d72619e19f984d76684caad7d837212391c6c2ffd240d7e49b62fecd36bf455514f1ed87ce7974f5f3b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h88e7c8e612a68c2bc5620f7afa1bb01ac94d4559388747b3b26ac37bd7c7745a7b163a7a4f9792a3a2b205e80cdbec06b347d3069f634b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8ca6c06fbc0e37e20b6140251975a2270bba2c6d56b62404822db48856d671e51eba42ea5ce066e0913a900cf9a5771c24c5d1f5dc4a5b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c7b77e9eef05bc29d25374e5207a773f4163802b49d033f19192802c08f51af04415a5dca3662cd1d06384eb2263402f6f06bab36d21d6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h54469aa1c9e08a4eed7845cecbf81773faa038555c3eb01678741c3e0d33562b43900fd44999be67de3ab58ed1367d2b388c0268483bc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15a11cbdcb788329a7c2a09253a4fdaa50e6c8d2f6f9b10d1852cf289dd08af9dccce283619448bf0ece675828002cae0c5f4a23e0d7d6e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16a3fc7d7b7f75faba8fd6293190426815b710d83c3f04e4eedbb871464a1454c0e717eb0bbbc98929831bb03baea16880e0ab07a141d35;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd0c75f92672b1bef64ce3f8d64e3a4d3c4470c1e92b198e9da307e7e1b04fbe698f9adbf82208e1268a3fac1df7a17cf6b6d0c474bec91;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h80ba5c795c9202b2a51a721e45e22afc46c1254230ee3412d8b98e45847ae465feaac30bd4cbc91a9106f957f6e6d83a01262aa9b1f14b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e4f263e86a92a5423f6feb85a3e9350218110155c94e0687ea20a6c76a99a8dfb95446a22116006f392c1cd2d56fcd28c4ab3a795562e6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb1b7231395af48ee38bd6e7bbda7ede82ccde8535776f86f23f1a36e6759fd31df041bc726def2ac1510b5ff53d6512cc58ec10036d94c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f2b5ed6ebb4fcf8000745e5c3749449cb1f73d7d12839e3b9fdbef8b6d507c23d028bd232ae00865f40725851323ce821c5220e412dfd8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc81b68f378a9987d6e426493023ec658c6923168fb8ce3cd45d8403cf031ce4962901729d3c16ee0a3f27c2b3bc2f4482a30a75b80ab1f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h111743b45636961da76bfe1fcbc243139f8b962748cae180ef8e37c23c84e6fbd13ee09e816e98d0f181bd473c3659d81777a96b60e1337;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c584d79d035e6dd2075c060959508430037745f50d91c8d112c45e8898e143f988fbc3f5cc022c749759df6f8e2c55358fe04e667916e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15fa530802308003642bbbe7150943d88420aa1b65b58dec9953c3edbb48e18904da888d57cfe6e06217c8764af1476f483e0292a16f01b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2754ff5c433fbf1dc2bc42aef2a99da6e04af0c9c3e57d8961c84f98d631349174607afefe54a5172b577aeb56df50362615d12c35a8e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc167369e95d2a611a945eaf241b6939384c0c37c1b2bd1a8ac3a68fa8e48a0d05405d99844c535e62e460460a28ddf192550055292d7e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10657acbfa5f50dce5209b6f2ed00b765c58fbfced3de46587f29da4dce06149a6e69622220720c41345f6635e0b77ee5a131c15a0555c2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a6f1375f5d0e517eab628724e72ef5a5ab0fed82d7ca59df3eb77d88e2169a9ac910730a93b594f56fd594cec8da5071d50c31e5de9c38;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ab511818235d4bae220a85562a7d5db0989c9418cca855be0b6ddc5102447be9c293ee578943372aaefbdc183b608c3b359a241aeb008a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16f623a76f2c22aa746985882ee5a277ffdbddcce6d11f36f087798a49e4098ac7f419b18e0c8fb05303904e972aa47a8ba7e5e6191744c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9ece63a920241aabe77633ecc262103309c48b58375f3fb1c0dcbd36d965e7e17c19ecf05829152a508099ea0c0ba8533ce24ce5f87aaf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1608bab68665d481e82bf2f522e980bf5106d7f7a6a3d87ca2d618d73c569ed07f9fbea6e6ff15c13dae3e39f2924a3a2baf4f910c5850d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h67bde60933029528f8168ba70940904a03cbec775cf83c5c2e00479dfd8a6032f8df8f60b2a688ce9ef7924af3b01be5a0c6994e8d7760;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f8a4ed65c6989243511415be58a0b24beb83383046cb3ca805bc0f3704913b36f5f71c3c88050097300dfe0700824c1751ee36a1949bb8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h130df7ae3185b5475d2bbbee09664a04bbf12184faaae8a629bb5ce71db5b440b4b054a1f525c2cfa259326e6ab84ed2f2dc0e2cb7cfffe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c3dd70fe15576ec2e2fe2cc3d027695882df7b76bff833e0686c4d64c24e558d8139cd4db3c69c445e586250dfc75e5cd533158d9d48f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12dd1b852635cae14ff9dfa7bb35184d0eaf59d61127fe61edad773b1048f8233de37ff00a32b8041305383fcc55a99e35ccac7677c5e59;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he6a403aee25cbfe36adf74da05267c229668af0a438a9d45d77f80d1db88a96435d29127122f2bfa26ff352c3da851b91247400902bcd6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1292b67f91c2f39ea28432aa106620b35822c4dc10adc21c6f19c2e8cc93b1f29a0810c20e208398957b287592108379712f7be257de516;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bfd028d4298cdb108beab63afc87725bf21ff88412ef61761bb29e0ecf7b2b4e6b77eb71059556690a9f5b88d26f6c7b0cd54e97b6a039;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1595fbda8bec2f14a7ffc085b767a52618baaeb7b938bb787ee0426e9850566bfaf1b1873f4a59da59b2453f446d7e4ff49e86145d98c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9e21eedc7ade2164e0b8450f9c4c9c092c21a287fe0bc102a0467fd1ef11f7d889ac94894ea84aa6be0b7405b48e97f85f39daa08d9848;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12fb8977c5144c933ecfebcbf105aed46b90facd8f224ef73caaeadcd4143b0d472c568726bf66ddd416c4ad01c6d389c4235166f9d7ff7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1feaf97ce64626ec7cf5062946b8b7b3eb854d193bab099f82a23b2181cb9c5b48d4643c23a51772fcb99c3952cd922397463c134e9a57d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hec7b635beb57235462fa9f43adc5dd53c4a7a93c07e28c12f68a17512bcb1517948fd790a5468bd16a0613a273214bd403b33cbb1f73be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17e3347f072d038ef2e698af64600bda4464e9e2ccb9666036b20c6eea1d180d72f574e5af5f9067d0252402dcd360307ff497d8b14d11c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c282ce083f10469718aa04a719e42327643093c506a4e0ae9d2374787f1e11ab34aed4f71593b6fd7e29a5b7a775320e7ee05811fc24d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12626deb2c857860a8a15ddada238bf9a83ec97632d7c4b391da6af4b43cd09a2be428fa1298f4b938f07d837bf877e5b4c611cf74cb137;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf0df59b4ba72270dd06606cdcf58416c04072cdcbbf162622e99218316dcae39310c17cd6d63b4c64c4b53bc392da40227235fe3a3bf53;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1617923f9bce181c355ed35f22f70d2f92abb0ca741f99372e4d85e5be42594d57d38942b7f73e4be8fc118e968f4a631f80bdeaaa12f0b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha9e94e5bf609181d7f7618f269d9aab6b58f8b8e61de1b38a5dce5f9755f27893cbf1fef6c3230f665269e187ddf4a9f9ce92c867e73dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f2aff4c443cb92f1f458f6c1ec71af4be75e7b047a3c46ac433b01d767038e099c97d4deaccbaead92d6070fa40f3b3ae230eced22e460;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6dc445515ebe1dbf8949fe22abdd04447efa8ae098a32d7725aefbf5e97aac1c7f4de0714c090511047aff693987b6c10da5b607ec06c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e7e6054b107ad177c4cbe118aa824afeb0ae56a0c9e372673293ff10c5546edf53e40269fd77beda228ea8da060617178c8c371c84faba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1944b13177382702e0d86f8b22ca01076b3635b9b6e9813b4afff9d949b0a69a3fbb1a87e08ab93eacb69d9a6079649a1727892e961aa71;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6e44ca397d7f2cb1a39376adc2f4d652d3a35cfe6950599ef7d5ee10b39459b5905dc1db8ad838e9885bf2a04ecae7bdd5bb911003031;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19fb6e5b911b2a79cd3ebcf452f4876716d641fe2b49a3d50333e28b4e0bf560f416d95892d768fc2106574ab18a8475ac381a6f5026390;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h180cbc3636e8f51a33fada92929b96f0acf92bd146fce5d8323e45b974b282fd2f22d61ba8a0a2429e5afead391c68ec8dba32931ecb69b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13f0832810162302fe4430b3ebb480d609da127b7b352455a736ea6e3fa5b9fb3b38140da5add85356db13a0c9c3cb963a1064bd5d46a04;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16df0d6a9532dd9e2a2ff3f8fea8c5dc87d7168cab5266eac4913ebe19bda43e0c7b034ca150ec24d6f6c5a9a6c9e703b29babade8406d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2db3ac449b9df6c9e85e80997d67a7be6778988ecbe34f0df2b651af7b9008883f06ad80965ce557db0e1c10077f3f70686c3d294d451f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18b6ea4b5942637cf98020010506c772bee3d72d1a7f1fb4ce658b963e74cabd9235a8e5bdc60268b13ce18f253ddcdb47a57b680d961e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha7dae58a77d786b5629113bfb67d6c488418817be0691800bc729cf58ccb4e1a736061942c72bf135609b22a24ba958284baf87b148c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18c738d56784a48d3c49d859d8ece37ae61c70c0492126c8854dfeccfb0dceab1600798a0aa6d1d1c6586a3c34ff623fd7a16a3db010361;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h347059575ef1d3f13f174b3fb98d3e47c1c7c2c646e059fa968ebb2d2177aaa38d2ccfe4e085362bed12214b3996f840998c018005a7d1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17ce6bae47d7ecc14f7d35cff11417cb91e7ef48b48ec231c8cf72413614b8036823a3debd81ee47a6a4f8feb949f2857909ba4bc5f060d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c3933a5c1104e265911935f48f92136666c038cee57dff03360fc74ce8e36bc56b93e456f3673064996e29be7556e131bd4034860cfc11;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb8e1dba481279447dc31955d41cd60e622cbd5503356f0a622dba506ffa4e065756ff11c7ab0a5cb1f745e25f401e39bf1e1394157a3d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h161f4934fafc99ca0b147f0ceed0f1ef6f2e897eaa3962f4806e5f1a67edf3eec911dbe9d0e61e3f4ea84533a9be7f3897910ad8b3d2dd5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4ea22a97e0302a635a38efda13ba348aa2a83587fcbbad0f6dc4e11e88e0abf7959eab7f6f28ffab726bd456aca63460c5cd6103923e0f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h51ef11d7068392da0957da7552a38366a204ff880a1556a7ed4775ab57e13e89767e45e8280931430be7dc4d12042ee059e02efea3a493;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h787e2a5ef4d956b10425d8dd3304331e0a0faea9167a910b7f971388b2aa4f0b57487f70ecaa666873d69faefae1dd820c93606e933ac2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h635808a71251589264ae90ffaf80a3b2ab8f3e9ec52ba30dcda697a10028d4f1253f6b59a4598ffa8afc65c5f3b95ec8ef02293d68be82;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c1a05c077f35ac524d7e87142675af706409cc441486616803d69c8cbc8222e1c628d340b650a007f822728f22430c516a981e4526b466;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13c2430591fe12bff6e5f6cd753113f7e2bb7dfa69b71b850a6d0e7b6c2c0a88658696450c819583c58774b93124c16afdca11d54371661;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15e1e34570cdc5b40e775c9462930f8f3f8dc4279d2300e8e50e7d2cb761ccad51381c3d7d901f7fcaa4c003387f8e36c084aa6c358720b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e6a527de5a73c99a236c5fa2195669f463ee20918a86370eae42bf00ac292829b900e38b91da352d8e6c26d81a80f722b3276b7005b0c7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h833d5fde1e96f1a71b25111799747a857bc501c6661c772f5da7040c12c112b3cbde22c4d5439bf6284d3c2112078351fae320eaf62e05;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h584eb6364c3cf848f27525d31f243cf1c8f7295ebf1532ae3fd2f25de27c3a0ccc59b532e97334b18bdb92b475f5ca90f0b42d0779b334;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h90bff841e0b2f97656eec195f678cad26e853f53531a14d253811e106b181c7a16a240983066e30df17c2298fe47649bb6e0a1ad025476;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13f00b6c44509364a4feda4ffdda0b206c6cd6716e7892b032d072389924140b6665ac2b70f5390d53eff38f288b40fdafaa230b9eeffbe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7c48ba43e028bf77095192e1105990b57e200590aa6d047efe0484ddbe947f4f9af92596f45ab33b4753ee465f6dbc57d61b42d2cb294;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1930fbdca3c9e5c2cc802994b9b660a649601ea8b785bd52e6e164e2cb52a54b641dc0bb3bf66e08743c142616cfa756ea817af75b4ee32;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd8e488829afa085e76efe2299af8b649073a748f2a1ac240acc9715b0a913c33a79ed825f05b029817c45bf857679bb08328e3324cb91c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h101d186f721c11acd0946f5aa6f590983796536eea4079a048df2a1b6637ce1fbc7f0de83e0bf44db91dec824b0dbc09d5991bc8449f767;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11bcab4f75b1d126e763b4696b96066e67b81f9a405e18a65e29b961a626ced8374cece9ef7fa603e3a6608072c265540b7d8ef1e00f2bc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12e55a37de01d02255aa2325350b8e3ec9fee3eee8e41718f018a0b103c6712b23ac2f78273ef6a29e581ac20b3a62fdb8d5e2cffce7a56;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13a9536187fb4d8a38517be904dba1297dc987064817bd3abd7669682d57e81b1e56f7a3d8e153f82e0f66bd76d72722d20a375b6ced5ad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h196fc69b98480b56b4b57a4420ec467785e8bbeed5b43689eea53029d12e2bba7e0fc759bd1d0d1bfc62fcc1f4f79f0f2f0a91d2466261b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h36dffb2db3b5378a3d51dd9c579b6ccc10ca936c8c0be6ba86ad5c54772bd53eec66322df65a5d54738ce22e59fb2c4c78c7f62d8a549f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b50868bc5d87afb587bdb83ee5ee0654738c9c06431e293702748ef3e3e2c1a0f519f9e7f0c97b058968f9d88a3003fe8c6f1fdec813fd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf047720a0588181216bfdacf5d890e07a7d416fd3fa93ffcc5cd7d6d7cbf12498ad576e8e3571c9bc29b7ed185605f0ea7a32fef31690e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6ea9495eac5d1a7a9af9b776fc3558b3e02aec8de0e1b9bfbf6bd50a1d23babffe58688bb6831e10d74e2412bf4ccd219e1aab16419cd9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hae4e3ef17c8fc3d068e000bb73d246841dc470de47604a487b3c3578179b807b9993b3581ed6794911b362a8a007ff1097dc41e7661317;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8252f498dae3f9100d3febca3b74c1e37075aa9c0682cfec5c7657cec5e6b34d196ecf09b13eaa230accae0fce6dbedc70dd75bf5a9fc1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c7c9ebf72c8b3584d940dc00c1a0a7b4b9ddfe2da5547209b93fa699501114b6d0254ebebcf76a42ab91951cab7e783df6663db43676cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1966ad7f1094c75b4af11ed8963b21cc8b26cf1d1c6dfce7914dcafb657b21ac51f9268bd33da376002a278a3bdf46f7c024d277de4bcb0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1afc886f321d9d5c2c3c9b89580bbbe76ea62a5bf252dbb7a94e4a3a234d3ddc171ecc9ac2d567872b86c50b407924f2772c7ddfd808691;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7691727c503d005f78bd5b7b0bec2ad64cf1da5456e807aff09bbb0e6bf83b7b017f1669b18d308595c2b2b2a0a8f8d4dbf08166b178b6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c7e7d2121c520771fabb9d582e2488e660568129bb2511c948168f9002126b9baa99764b54cef720fa01e1bbdfe1bd84b82e7c66a3d4fc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10460cccfeaa706c38e9e232e8214514ca83f83155514948d55fe66d7011206d19e65ee0b203920d1d41d764b0a9d0c126db9bf05c7f621;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcffaa634ef7ed67560654e8111664c5c0a61e719614dcb2203174e09ccd711c043b490214cfae4233f9391ca89439967205809b6b597bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdf822d6344a8835c7d1f80093af45a29f6644fd124838eaa1faf5b5b38d4f6af4356fbc6958e055ffd7a9c1bd7db06236ff89c05a2ba31;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1794339cc09982afc8017ce7895705c18b3d47c1101a686b0394462511e4fe295ff1f4fed2184bc3cbf32eab84a79b8e8b28b2bec09f413;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12f168423236de79a6fb1bd1dba42cbbf6aad01d424f1c85eebf6950b673eba7007119147453db36521e0c7ba00af4c1a143bee9080774e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1397bc889039a9193e20d2dcef4cef4c22155def0d972d44ee855e9979af770a4891e2d339af51523088b45ca9ba1b32f31a0d426e0f897;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf94767a3af42a900a938457b08a35c4221682d63c4b4dd522d1c58637abda25514a134cfd1c4018ab872f1f768524f86557d049eeeb8cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1165bddbe16133c656dd2be924047b72901e54913c753102b818868d2c219aaa5271d6b8e348473b8eb15eecddb9a82216156dd774cb3af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h417eff293fc8ca7797d3dc4a6f7626262b1b5336f9cf52b14df739dc7f71bc197eee0beabe8162b2dae74a73d2d6975c2373ed2ad7e04;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b81fd0172bec535f57830439b67ff3d176a130373b66b3ff61d4641b7ec13e64d99f3d9584686db0bc1aabd1988c09cbabf85e112ce1f0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbf0deef1561daf70bc27e4fcc1addb1f8d521fe3334a8698a2261ab92a5453f21e122bdd255b899b2cd6366ba8c299bfdb48ba08d2dd20;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h171e9120c296833071a69cd8ecee7d8d92df431b5f3f0fbbf702059f7fba3a0a82f402aac56fb57338a68b96b982f6d6766abd3194e3203;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a347c09e677aae270249e9bf6b9b6f1000f5f5bd469153e8a58acc26045abefa571bc25de62a257957a67be569f9680245fd2514e1869c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha314595d28d38e0464f91b23bdf1512839f43b73a2b0f70b64d8ec3b0453be1b7093e670bef96e08a4a3d1b1ada024cee7739fc6d96345;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hed4692875f8c29f98e024af280abc3ac4414410f20a679dbe7ae74ad8d65daea1ed84f4ef6dc0712e609b89979bb47be5be501fd598213;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h114a89e8e985b0b0f8b8efb550af53f604cf101dc215110404026c19e6ddaaca7bbfe32273538a1bbd428ff722d27392da723d1de511ca4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb6b25c1fb296540bb226d210e7d8498215f0b55b69154184f40a1c1c57bd307a7cc19a2eeca7b4685608a9b9458194a8c6097e351d1a69;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b94020cbce9d5bb6ff503965e616a75f181b8d559cdbaddfd3f6e05ba56c31a32515814c06d678e748aea0b9ae2ba9e8dc01ce475c11de;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he81b3dcd43b0e3495d9e0fe79a313e30c1b6460fceaf36ab0da4e7fcc8a52898de6b573642bfe14c8f3a9b6952c4fa7025eadd2feee1be;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fb692f51657ff3eef453362ac232a7115c4101843a731e20a3c7f131f80f616cf051311c379163e3300f75d8d2620c729578fa1349d800;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cbbe953a0491db3536fba70853be3c031b57b6d0b07bbe7ecca182f8223311ebfa293952eda9f2983b4222054b477fe5563411cd4bff0d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc82e748296c52944174b284571f7ddefc711b3b9022e2fa5e356bd98d3535e3dc71e7478e882cfb85f0b40e95496287bf9247ce0d89bc7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e4e5053da262ea0397ac1b984ada62276e65222e57481f4d42041568710cffba505b7d696b6afc6b7927c2db9c1e15b89c092218bf13dc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbe29b289902bb49aabd431fb946991b0c0e14eb51238e04f5aeb2505a652ad7014ef0d12682c21f7434e52099e0a5857e9bab6a7fbf9d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11b4f7ca44ebfa2c208f969e543426d2452620cec6d39b3ed76a4fd264a4c4e07145383284d944d732657bb5523add120d029048e28207e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13b3ce53b84234fe7a3508325ea5fe795d69cd93603bd8d39c0f92fb00dc9c9826dd16d02b0f5db76c825c011acfe176e0282901d339f52;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16c049c54fd9c178cb3b4652bbbb9e1b3950515145c9c6c37f259f2be0ccf06e8d84f3940a46e439c2a2cce0824b59b0c637a444fcf6d1f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18d61ea44ee447542d5947da4fdd3a18af03799c1ff55d6cd9387b0e8abea8088bfff737868344b40819bd2ff886b682482c80e6783a6ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18b5dfbb30eb5daf3512f26533f05841bd2fb0907ca61e219b76cfe30581bfc7bcceda16b0728562bc86a9bef3284d64057c5618285eef7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h70e93f950511d0461fb54678aac97f9ea2556d26b929d0bd9fe25f646f05261c295895d5bd1c9ab6475cb9fbe88e94ff214bbcd951c4cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7f5bb0cd15590ecb779791a99fa9c2480a2e348bdb64ff3d6c329eeee65c8a943ba55ee0b1d7a6ac032dd75f5ee250c094749513d43a0f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1abf0db169ee89fa34fbcc9c264a25aa836e8f28449cb6cc17f1b6141ab8a28ffaa0f398710b7572a8a2d8f87c194c0cc2cb5b4e5a8a852;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc9f7e671527e0323cf503ec0c7b2f33f6c1e0763b5d5be968a825094e1ea5fd2c3fd143b3641c5a468b1ce46ea839e043548270268d581;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h172b487889bcf9ee4d4a0e9c2340275444758c8ade488cf2b4bb95ceced73afdee3ebad0cb1ab64bc0ea48207510035e1f10658922869a2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2005c746ff1f7765cfb76f7cc4699535137ac6ddf7ab9d89d6286021ae046d7d5aba49289ed4962146456523125551239b3619f2a3335a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1959a11f9c21ac6711aaa6f51aedfe3b21a01cffb649ba6d96089a6886357f897f5f4dd19e5882938302ad5f9b3fa426387acf0370178d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14ccb75466cae56f5368f4b2aad962755f10db551e55eec46ba7d4dc4b6e1ade5c8ab6220f94b8822d1e55757f02ae2b97da1b55d40200d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb8450d5023d592c379c2edc2f401e4731ebcf7942c040692dcadebd44558594375e76ab23d535e496df4b6ea09c82252b080385e798f05;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ffa91f4dbe67e92cfc7b407933eb21c7568fe33c67229d671b9ea54cb606f7ef429e50a6ebef3e439fb9897f40dd2ec65131cc14ecb434;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he9c8024e30163e48894cb63c25eb8de9f6749109ec048d31a52230bbf1d1f877810d1c8ca985cc093acc5b915b7c11fcea871732704ab7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h914e16d20e859022c581a3b3b1ec71cb2eb5fc1d282b58647560a0785707ded9441e1b5e6c16c816d8b608fb9b090b1be00cfab85d2dfa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6d11fe55fabdc26b6bb70ff2f2fe5b3d4eaaddd5dc38a4721ece02fe5d0457aa23cdadcb3ab17744fcabb7f7994667fdee1da3c38d650b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b60a0ec17b9e3f75accd72e181f13052122a9e13968d58aef71dfe1772d8960101dbffe5fbde917fcc163fccb48d69cb96de9c77f40db9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc54b2c3171d127f7f86977f8879de27e4dc49c419ba67acebe81a44a3b5a8d65d80bd757e81f6f65888bc6d58b0950ec171b7352b74be9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f10e5825c5bb8e09fe029f2f5b06b2d56631ab5f4424f298012bd9c319551ff5497d1bfc667c862297c4bf3c07402530b6fe8d129de0f9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h808eaa214f1d224b173663d06df67b5cad7bd1d612d46de2052aa43895aeea344780c9779a0cc9a330656d2503559636ade9581337872a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14ae7ed9935e42fb2a48c8a322cce15e68bf1540017db3619ee270ce159dd00d013239420a9c070cbb70907da1b908ea8b8b15320272810;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bb6cf87e24f2be9228b4e95f2d8121f9016baeea7d351e65eed5cf4db95b429888a9193f2649c61ba6a09041e0c02bdacdfe5b8f128b07;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ce9e380c5cfaf7bee4629a19b88037cae1a4a7d987daae6d582bab3e7120d1e84df17673e8eb5f067a66dedb3d5a5153d1586f38baa720;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h511a83994b577bf1c9310d45237edbccdddbc6c8b35638255fa8bb09f28f11a67ada000de2b570785775101d85a19e1635d00cc3cb3a00;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11862caf74b448f80b5c0743a81eee1253b8bc46f00800c36f393d3682bb7b30a1126e257878aa6ec861c9393f7dcedb276cf05f3a67d7d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h140370123f0d121c5db94dc8792203be1f163431970770fc934b1385575af96914dd1c841114578e1115d7ea8996aacda69eb9710c7b41b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbe28a70610d0d70605fddf4356def1d99e2e78594c3ad894ca9af8426a81aad4199da1177e9c7ee91ee74e3bbedfa8e08d3f4b81f83993;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d9b19b439a2b52392a219a512d3c4f131bf5e11cc4e042330d67984d263451d7d92cd0c3260c9ba8fb81827931910ce7b3280841499e23;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2b4a7ede148f574e00652c6ee19f3690746a986bb64c248799c67de4c66963f2a5fe778222065b6f585392f1ab9d4771d42335da1849b3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18613488bb2e6b353db804c9fa5a9012202ae07e448601d3759c110748702e8e9d319990735cc5f4169b8d1337668b3e32aaeff31826764;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ac9751cd8ac7052588f16af4185729ef2737fa226825022bff3f70fc76681f8161f2361102f039d0264e94a7781f75d6e3d86edd44349;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de9ca1a7609333e1a9c8f06d8d5c5e3c0af953e7fc7b3eec05565c83d0941f6ef607a1c2e33b9d2ae45d535b584ea77190633ad52e5f18;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd4ed6749b9b33e73c1466e996c7d3cb0d8bdb857f0896fb74f210fbb4cca22b5f6db3f363badb2710b457928b2d03011f5962b566ad7a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1313809b4067b2f4f7c28c402418556d587620fcdb81c2cf3120540a0a4531c4bdfd625f97539d2e0802080fd51a38ed4aaeff3160fbda3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1417160c287386ae5f2030e4f61a28e159586aa360c78d7a49b7a4cfedf5eb7ec33572e58000a4fdca98207cf6af17d43aa63e63d7a085d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1163ff7197f9e9a106137506c32cc9e769d32e1834a14f2d56ec022455b4415021456ae114388bdb204fc843227ad6f4f6d6e08268373f5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c475071612ef00d6acb9bf7de78ebb7c549c49dd0787937c6279f95ee64143c9de813088613a3c66fb693266440905c7abf2a78ff2d531;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11ed4a9e62a2ad3df66c24412a55dc59a07e91ce037641201c9a5e589b53bf7843b1a7931407e2abd61c798d1125f63c633f895b01325cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d23718fe931454848b9c1d2737f74e300f8d4ee547e7977fcce8a2af5a50f468905bee7188087932e6d477ebea444c097e1f1c967d8196;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c81a05ac6f71031bf7c1cef23a5da45d773b4974f3fc3e40f688caf5563aab13e570b8ece05467ae3f4a35f7fa2a3c4706942e5992f05;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h21302d0b12eae59f9da9e4c55f43020da2f87724d7e9b5897c03cd444b7fd5e199c0fd885e84c281a941188ae8498cab1aa1229cb43116;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13a96538d30b667c192d89e917e1cdcf1281a0d2944f9927cabb2e9b00a56c6174679db09f00022be49af60a6232d2bc3d44e3187dfa250;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f9876b0892e1d5c4a46a4b7d65dca997501b4db9aeb73c7442697b7703409a5be12e958ab6ca37c3ba6a303f644cae435704406203f167;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d0de57f628e7fb0ff5c0e14887705187ac9e55e181093863addf33f1f0bad91aef5f00147244bbb7c5ac11bf998dc9ed5c8978f3d08619;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1999d457726eff295b831bd5c56416c8ddf4154663b3478c38600328fbdbcccc6f0a32aaa864e2057d78db8c997b619a0ff43e2e98edb0c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbd9e349a3d8c9f508a1d6a48345f6983c6073a226b406dd95cb3a48e34f2d2d88a6e6b19ca92daeffef8424973b4662c5474e5198b0feb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a00cd579ad05d46bb4c77f59300ac559b3fb125fcf95ef8f8aa2ac2d1341c069c5a193133ea11d2b4c3aa853509c17a4027fab0381d965;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2e34af66b7c0dde38c730b1d4d3df84410474f1ede687d79f70982cc58df6cb003637b095d84b33d4e555344a3c0d22f65355194efaaa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f5b87f40e08008079a56653e0c0362b26b9628a78b4134fce80569dc8cdc85443f51db3518e44d8904c2a146b007956634ecc4f0bff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h152546ddb3d6312ae335545bd9ea5119ab02e7a6c6979f8e4a2d46e0fda44351cd158e4abbe2f5f55f4e9b39350c4f1bedd61ace8e9a9f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2a46c90d1f17c87fcbfaa35da64cf64d0f87455b4b728574025e3ce108f874ff65ced3fe859b8821a22590e704345497d1bbdea895bb65;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haa4544110b84adcf971b4809850c0cc40cf41f16263c75006732eca2c4fba202dafd212bcbaac92152353e416cc3e67be2d766a68ec779;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h369e234e24ad9176742b6c1b1af43c5e03fdbad407231ac4712261d222215867e3cb0d8077f1daebd2c052a24da7615c6868c380a7cfa5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2f9b6de1d0cb78e75b1412ebf52e82cf9d061ade0b9c05373414301fd35c06d341d9748ce9f33fd46214ade6186bbb68e0c7055ca82ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h32b202dbacfc018724baf78b150cc63f97bef2f4c2f3dd24743f9b4f34aedadd829d34c675cb32eaf0505a3dec89e1d626d96fb6b3c433;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb1bc029d4df830c6daecdf399efc8c3b211bc06da0acf826bbcb5213b7b56e28a72dfcf95ec8600dfaef172ad80bd7d1b33a9023d24a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h106618846756bd99ad8648755c943f78783cc0b2a03c94a4e543a117572a15ed167d81c43f821e25a0336bae37177eb7a7e9818531b0366;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11eb5c1a4071a06d95232ea53f51f7d0b1861749895f817adbc3c17cc7da79cc95385e8b41cc250b421b2100d93c84a9777f2e1c37785bf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a02aa72ec57fccfe28ab29852f735eb64ab1f7eeda4a70a0f98d7bc7c82640618e41b4863f29e679be374ea6ea0f693f35696d92535dc5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc7c9dc63bb58de5729d7b23848b44970410891c02066b77acd4cccc7380973a37253c4925b07cf6850d4319e9ae0a3a8cbb572a9f58d6e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h287c857bd928f3469f08bc418fbabe536af0e1ce57cae9c1c97c5f6746830481413cee8fdf8cd597c59472d8f56f44f57bb1cd20ea556f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h111bde9d473c3279ae5f7715a5bb39ea8e227779a9db569cfd1ac3efe9580960cd4b146164885e8fd28dbb239e70663d69b4ae5c6a3c22d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1150d2bd4bc3640fc20a9b4fa87af16ce0196954a28f06521a3164b9ee758ce2524c5da2fa5e5ffa4342f07bca0164156898006d2e4a0b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h62ba5cd37c48cf2cc80f4df35044fd43468118409b9e848a521bc9a299bc07ca963a2f59c26c49d45972de392675bcee061aaff1cb9151;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb5fda3f689616fbdf1f2656a9518ce61a2daa7233ce5f7ef0dbeb32a269deaaba1b0be4827b4f236a015f2bb196edc57b9a30639950ef1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dc8130074349ff2506c2cb38779c3f472b779d6af2d4e2e7ccf0f62fa5955ba258541295ada17e43acf617ee51c2defb2be3b400a86bda;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc5105dff831b0d1eb66a66ad9e7a778be079f5b2ec45fa20e4471cb0f3bc95940ea2254ada8aa9ef8669389abc403ee76e97c469889282;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f7d66df34f8a174a18dc036b2e299693d2a5107acfe1160e5cb6cec3307f3bcc895421c6b8b842127a10a7e0fa08b29ab76e7483624c92;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d59963dfca5bd0e8a71ddea3945e688ad475dfb37e2418b4b1b06f9d64415ab40daa23547aa970078107be332c6ef942b4ed7405675e0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ae6b9900e1b88fa9764ee7cf517ca0526d1802eda924d6b399145586ed98292bb2c4b3d53851d78f43b3f01cc7e23b6b426da271799730;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f0ca4079d7345d168bba5ba964008ad7b1e00562f573e9c5797e2b424f75f4baa99c248ed961d56727a33caad73683f9ac35d9cba8b9b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h134107c04f04619eeaf69fef6c47aed9851e7c5b0b94d10524bace0a6a7cf02dab2187e21006b2865935c0de20780e38483b4d290f25dbc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2899f1193f066d41998d7681bb2c09280720dce7dcbe32e17df44318ecb3d7c0cb32c2bd7552112f0b7e7284d76cc72ad11466a1af5466;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b9ff4c1d63e04d85ff5183a7dec8d0a51dbeae5782e478a1a92f257e8f1de69440dbec7216d4c0365b038f22cb8b2ecfd14ef2b9deda22;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h199cdcf5c11d96a8885bff7f868a8856a59edf2bddee7a201c3fc2931c9eb44db40d0158d9acebc8d1fb9ed29eb70faa3faf58d29c994a2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h268caaa8780e174d2ca79538920a2870fedae76b82aaef7cb06a93b2a5690688ad6355438a78351f5e9fef48efa54ca20475ec996f1405;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h39d5b98155b39a9ea950c82a992362a9587ab308e8f2f3a31a97b3eb06fca3af57f4678a6a15ceac44a19d67ad633e488f1fc41d9976cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb996a3c044b23a0d4c1a96952f09a355245813fc102360f1a6a56440a69145a2b5a5a3baaca6e8eb2e91082271f7da3119feaebf9641eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d7b4d4667378caf75d32ff09dd90e6ab5e6f84ea8384afafc1f5d6ab44ad2f023e3f17acceac4ce10afc48f82b5a5f3a00577863b7cc18;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbc56c3b18a30988386198146d7b37a3aada340c6875e73dac1263f7836f648765564c8b9770711abdb16001358a26d84310772f90a2893;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf1807c46f04f7351dc431400df4d98bf91f280f7d1bf9a6f8ce64ae53d68d2ee7513faf6ebb0d4fe7e2cfebeb40a0f929cd5d52c0dad89;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hea7d6bd44f69585cd90fe2fb48bf86a5079918bbb0ee95bc18dce985e8a6aacb9da778cef75f608a374c3a6ee328dd400f0093163be124;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a228d143c9d06970413a86a49e5554cdc1c8b83bde9632c7c0849348ba6d204c3ebe52548850b545d3c869fac2a022583eb5178c588d4b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ff7b67004fe20e777a69c4a9b48c363216fcd9156f1d32f8023dcff444d7f99dbd6b8321a8fc3b46f573aeff0034874043cda54c555c21;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7567ea01f26f7a67169a9fa0c3920125133df1473eb76a7f58bb80344e358c85b6c33fe1c0e3d1032fdb9ffcfca5741160a6368af172df;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1154efcc901252f06adb1c632c86a2c7467e0a111804a71d599f1f023ed7abc7f360edc225de7b192c0f1b6cfca254a63cffdbcbd6cddf6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cb8a19b1e2e731fbc07da0683e9c3502d5e05936be8368b8c95f018efcd07914c18a44ea111209ebae2332f1af7fde397e223ffe8eb84b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbb11d4c452891c1801c1482e5f69b7912c55dbd54436eff16af4b4016385fbb8fce2f667cbd9ef7cd3573859823db87167a7a7ffd9eba1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd00b150eb6e96aa51f1ed32444e8bb759f1f257b60aa494701bb0864d23798468ba9f15039b7f2b768a5f82e96bba0631bd8d4ede576e2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6c5507ec6d8021a06c640c1e70fdca41d3256b4a50be9c0cfa2fae2c0e89af66637fb4e14601e5bd758ca7c85fdb27850d4206e06906ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h150ea084b549e21dd909b302321d2932f822bb325f147568018860789ffd848b5eb26cc33af57e55edec7c72df67074f02033b6a4076487;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha368451e8f1e7c6057bb20fa847a81cde13ab5c2c15b3c5397af8be39c24dbc7b9d4a51865d1ff1ac9ffb398619de76138b0218dec1b15;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d2f1bccc49060f477ab49bd32110950a78e7a825eaeb26cf4e6ec2bd5db317266509839dbf4b0862c74a641f55ef15beef1cc44e22bd77;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dff1f7080b3337dc82860738ca672ff2f8334bc38ae16e5a816031543297e18e624004a4708b5e344ced19ba80de9fc7553b2ae539dcd9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h47161c1b554779ae15918f62272a341c3fba360d887a690ea14d0a9461e54b25d5d0fcd4105ee8b0348136628eae78ac71b85b68b96188;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha222d51d20a69636367069aae553e6343f6f51bb6349bbcd65f04221be17f2d85a34731824752adb594b11bf43670cb5e78f1fb6fabbb7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c04a5b39557038d8aa7d89d4d30a09c451b7b8832c34972693a379bb492ca824d4f920682dd81dbeb8ab8db245d268951c3f0930d34195;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f2047292d74e3af420267be4bd8bbcd31de24eb385c2f3bd1f8f0bacf2005f029d9e8e1ababc20746a5044a46281b9678ab10f529774f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1664940010e216034c672ccf0888e162da20417f3453d2f8f44bee07808c284e07aa3e55f0e6cba6c03cd5d074e08b58622e8aaa2d1f0d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10a0ee11443e619ae2f2df41aca7543e83dbb53e40adebd53f788a04e04a242e7d2b8a038236d15a252d8cb6a33130809c9105fec784df;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h53fcead6136a594fe6e3963e3905ef28ea6b65e582d6518756f32ff1289938134d8d68ab64381010243f619ee363d06d710c7087d1f48b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13a5d91fc859ebf20b8b483a42c111b6c16518262804f96b639594ae60ee41249f594c4a6d5756691c447968b97149837b1c21e0a195532;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b64122d1a46825c57872b605b6080280fff99e8e57925d9d58e7fc51344441064877e97641ec87476e68c597f47eef195e7ca7210566a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5c6977437daf39e95dee205e6f0bce5bdb79dee942c4fe942f1dc28f3320bd3d18ec4b384ecaddad898bd5a20c8861f1a13c9087c248c4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1089a5bb50bc306b44941e0ba779c265ba486725e8a9624ef71e97d29e826881ad9f2d8d689925818fce5b51fa140d4f1304350e5931e2b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb747f7bb53d6be18382f9b382f9ea2112b1737c0bcf6bd46c7b7b5f41d2acf072c3f4756f4b0e26a5ddfab2bb97321fd8989e33c236969;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ce0477b7b86ef55de3e6ff69b657220e56bf034a756ad64b010d6af0288faf24ba7502a2a66666a10c506e49db5574520e3291de658c61;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18d87c744c34586c221cdc673678f683560bbfbf322c24dd8f52da5db86264296178d3aaeb13f6e181e29ace2e94c03a77e77f58092574;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8274b75e516b25167556631c142c0bcd6dbec3bd8e7a3621ca722cfb59acc02a8ebb6401a307c8188b8c87376409eb661eb3885a643c73;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h26ff2badb76cde3c7b5d64a80e29cb4caf84756de9bd49483d005bf2d8391e36808ba1e885af426c310f4af2edb14ef24effac3ddb4760;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f5744e73cb8f0975e8d203f4dbdbc08b6a3ddb07d7285e8b663d0263118bcbf59d8de725cc3c25e0ad66d6bf8283e8c5801585394c98ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h57847b429546be8ef14676d70cf4cd9ebd30121865e8b1c2de61153c139480828700844b56a31d349ac1e5cc6a2203b56fbd79fba736ba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4eb43f12a8cad179111c864eab7272f623886f48ad5173899699f5a142a3572768b7b1a46ad15e7ef0e98fed2777a5118f337c052452fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6b196ce481124e7bb7aa2557b62cced7c821af5b50f2019f54262cdce00b84ece6b77dfbebfd324d8ef0e1344483c3730fecc0a39e901a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h150d49a25fdf7dfee1787884194991bfe23b705fa0e4013f41a1de12b69be6d9d43d4d5034057bbb37f4aae98d3d47dea10ac0a6e15c12c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcb0a7d518a1bcdccf71c6bf02c3a8bb662cb19a14cacc28570a34e18b04dfa36c9a1240120511750008aa263a4a2bc9e723e4b3f3c2871;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8a0f39ca43c3f5e924266d39bf51cb18eb49e363a5e1f7acc04678e4493b56ec9c38878f89751435a3562008741ff3dd22c01b02164cd9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cedc5c7fed347e7d4459e00ebb0a6d1e6417fe18b1bd9fcc2d60747b4e3c88c700e130160c00f977c8ee27152565d3513e73260b1a04c5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf9395c5c8b6140740ce5de25d6b35995cebfb4e98ccb18afd52f5e0636d3fe18bd592f113f54276fa3690202a359493f4ee0089e3e48e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7f3c2c6e12357fba204438cfad82561dc29dc939669d9af1b24967c054ed2b628ecc85798c256fee2cf2dc536fd7bd1a4460119a9648ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17535b4b67d8c4c485d7296dbec2a69dc9b0e05db11e12536a4c1777ead78a14bc5d1ecac974496b1d0fca10b43ef7f9a70cf89de264689;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b0f90e4f8631faa17445f4698966573eed6ab6b8b6b6ad1accad148bba8c2283bebdb7955575108da00b69390efa748ec436747aae4f2e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17c20c679fc87063df8b73a5b99fd18ac8e433570cfc4781b9283aa786e7ffd2a16956e8800dfe7ade86105cee8f2d5a7207f8003d6b369;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ae85b78152e0553e7fd81d5fde0facecc8f69b3319b16fc40a81f3d04d792cdea61b61e479fa636ebe2c3fb6e440da284a226115faa01;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7be150a9f32b5021d8ce0d0f8343b747a00c19ccb81d3519fcea9771f665288a76278850520e53da6c595b607215dceda8101a1e6f4fb5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdc41a2ed619ff5d24e69345ed7868d8afdb012917dba6e6c19e846ec61602c731b56e8fa5dff489e0a11ecdebc04b20ec57f863020efab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5742d1b4a30faa479364e112b4b2de5606e55a6c190c6b7c564a5d4ca535e8c7f7551821b562f39c1ac605b25e48eca72657a82d41f9ee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e058fcdee77a55cf3547f81d052484311514f090517c1636d9abca94f1a3ec5db0bfd3313f8e51193111d5144f2a742e047131deab40bc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h104f470ea00abefb8d8e87f1cc343c1e1bc586b07ea49fa658c93a6fcca116b8c5a37ad1d25153ae16994050ccf085d5725de6cafd2766;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he89fcc48cf7d54ea135a39b6f6bb869dea69526aabf4db132f0258cc45ee7019a4e17b60fd3aa7208020ee9745bbee6229308cb7fb0006;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd473466214a6e885f1f27346ea99832bbe00de10d7266f35a06fb8286b080501e930260ec3211b44fdf3a09bfc547d9c8ac5470daaf78d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12ee3732bccd7ea247006cffd4a57d7549bbbe19d536c3b5d6ee74a1b10745de8516025779c8984126f410e9e4fa9dd811dfa860f821f2c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bb0ebfe1e96e524007cd87088ab353b2834d3d43c8f632b6e32d114c634d7707dfe92aead7c9bf7c2dc89db14deb43aca7621ee1173be4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9bc1b014b399ecadf25b5aea9a2fad8b971a3428f691952d90e7ab204f1888e291f6e6b9dc50d2dd1f82f85fcb94d77ce178345fb1a33b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11b708c80b6f292b431376f8dcdd84b3c8979f4b09adc1869b0a3b144c90c183e5b8b6ba9ca666c4942748c313c35b75754604c795b1c2d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h69601953ab6fccff03ee0d7da0a87fee20d02209bab991113d70b51dc7328c08e45a5f72b89a37fd0045f471910557791304ca06de6e47;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4ec54f2403cc72f5ca41fac4667600d9440408e689661ffad752926c0d27b3ff9cd120eec55e5042df4eccf35e373a071d91dbf13142d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h525a5d8c89a83b9d01c06c3146d4697b39e47806e043964173ae965665967eb4c0ffa536f1a4aa01eeaa556021457d9669c04635cec29c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h773709c9657a92774dbdf9942c0caac4f36b7ce12ae0a1944e5b5151bed7182714d99b741b96a41e7ad6546ec4992072f5bddc31d289f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18966a946d20d96b482c74cb4dea82870114dcbe2ebcac74a965c6fece82436a9f3f63884b463a5c43ca0f87e2e4b4ba6048f13aaa2859a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cf7c549d255939ab3ed8051e766584456467b1d461e003116c91611a92edb983d2fe32ba1ad0a3128527d43ef2065d4b0fda03cc7c7350;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2b781adf2f05c98f709ce800f1bbcc17282870638a6ed18bc509b671c6826e2a7031497993e95c9411b1ae94562ddaa321b5120bd1ee5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3fdbce56beee0b356cf5861dbebb258a714cc6d5aebecd7a29e807b451a2aa00d1644cd692c10840bba132b3a3cdbd0e7fbd60d1143235;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10be059e79185458195597e4979404745c4731e8f24ebd731a294447d45dbf654006a352bd7ec0d5df81c7e07ced107d81174973eab0176;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h79c599446e62fca4dbd7915384f6fc41ee8036f383c8c97f267199a01c445ef3b8bc5dc0a3b942aca8518abf7b5610b4960333bfd10dbc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16917007fb5ce8af71f870038b653ca94f221f00776ac2da77bea1cc350d09fa7dc307e199f889c9d2621f5ac8484ec363c6d2feefd4e17;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he2627d2d673393d92c861f27577aa918789c8eb848c7a39f87b239d396fe41d01b2db3f4aa1ff0504394ca6d015db7cdc93a36f898b736;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b5053a44d06d045b178cc9c2cd9bcbb87697561c4704531db5333e8f390cbc95934240fd22d30b3e59026fe0914e99c793b351bd21db43;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7274bf0f454a7885a8e78509da1209fd27fde7166548171cf4871e16b2a06e46d05d3b9ff8b71ec67cf2e7c44858734a494d0a456e4df6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8139d8e852f7b766cdfc14d9c29e6cfe838ee1f9800795835f7a3ce589efe063f72da2400a32875d1a9d84ce372f1cbf3a67afed0a6028;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcdc8e85e32ca71bbd73fcb2c1ffd2fceead373a0afaab4b7beab29a3042f8626ea9e5afe82e970043592f0a24da904bbb9866a99a5fcca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h111af77c97a0c531e42647ce108a17a237f42043b8b2407c619d4fe7f90077cd57b095a49ed2d2d900c80799e2618462b5bbda6e26c9208;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7023b235289e1fcfb80e43cf5bdd98ceab50e08b5d376a57642584b16e414bbfd884e3dd1d33498d12aaf2349fb92ba2805f01ea210e0c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5e5f3124bbf5baeaaf6beef5a650d716acee03daa51c740c2cc42eea908644802cfe79eac0206fe065d5f7d1ef71b4db946901dd250e23;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha4a7d63ddf5624e9e40493ba12fdee921b9cae841905b4914eef4a4c6757be6d2b6e5d309873ebcc36d5d3833e5c9108550a2f3b1c3ecd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd7defe1c1af38500dc9de765dd50cb6e27541ab5e23028fb4c3768ec69eeb6c43c32e4128c87569ecd40c3c292ba4f164fc490e56dc3d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4c693ccc3a913d483434587bb40064084153b18d280777b10496dd8acd2954fddb15c603f7de473651deb517ffc29c0e4dffb3e24ec73a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h57665394f221af50960ee9c85f913954024d6da8ae434e1cecfa8bbc32c026febfda266f4c07ab18634abec7dc121756dcabce89d90646;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1194c15a5340891b87c39b13202aa11c7c303f5a226974036b35d3e85f37fcc23b6624100c021786847dddf7b65dc93d42d5e18e6f684a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13791f554b4ae1b6db20116705b4093882994748afebc25e77ba6a60d62b4171614816f3f83a48a975b050b69fbe1926b4d94ed84af740f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dc3a251478f16bd54c3da9c986099a11647f27e46caf38dce9b9ced183c00d34f0c2b4e747b3b7d81fe0812c3401a729f1d1be6e378bac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15089d0d1193f847edc04fcc370bd71986b3e0b6c80a339fee82fb133e727b6f6df5399a4233aaa949651300a4f41114913467b754cc7a1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a7f87bac0959d1ca987716a503b8a0bea951a209c6331ddebcc34c0d3ac1b1177f10f6455cfd34e4e84ee90933dfe1bc002fa98e8b344d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf70d7dd3039a4371c5ec416a57b532c6e5f5774f1a9bf641d7009f651cb1b76e37684b531ce53b2eed7dcb981429c61cca524d0e29b1fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10f4a578d7d035608c9a3f85925482836d5c64d9a533e42be27d220af5b8a18757f382ee0b93f28274b0aad846b93ff3cea6977a0951995;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h137a8a58ac638a7b2de07d1b62826cec47a0673a6e355879447689f3d2efd4f1751781228e8320a197264a6ecd40c84836b698eac8497c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18e52db2020f1f572ac6b22504c32c3cf73007024a230839618300d46ebc6d2c82ed5d1f8b09e066181a02cba9c78a8528b7421fb0db4e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf661407a529dd89801abaacf10ad70474b1a4ce6331e3b497d10120f402689b2a66c18d9f2baa76b3b2000676c540edca3d9dcf586859c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h192e45d6afedc11edf07abe04097e532d6354d9ba740bf12ed90cbeab87b8882b32d5a5e70f4e130c5725b8dc5eb91300d2144f47bf856b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13238aafaf4095ad040eb4f819fbbc3c44add515ae31ef2d730ebc7331ee4bafc6136eb10750792498f0f0e084b55e4a032b2897dd70e2c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18ec3562aa75e3c851697a8da59dd8aee31c32c9e7e84a8ed75fa2b56485df9a116debdc4a59385f83465f84b40ff2f4a8ee1cbc6d6cf2e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h390f78599c7cbc58f0d7f43d490f5c77cf61b78e90e32fe6a1000a0a4472cb94ab064bad86f588e3d3f3f4bc91e05e272aa1698a6adbca;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4fd02d56c0aacf2505e4bb9fb65de75b91663c57a4f2d45c99633ff5db4aceb8f4fa45a41eb49a389ed663d8438ebd8b3b688587500fc1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bd050d71f6ff34cef6cbfd7642e58f98ad176283aa4da9e210ee6e19ee53fe716a21814c755f2ddc690cd7992e5fe92cac3d7f0b2cc96a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b081975a8660c2ad1de2d98d8e10be0babf89e25629eaa1bb0c93f00fd5fb674fb434f77670123bda52b26bb066350d7c5897c2cc793d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17c699f61a764b2086cfc6aedcb420dfd9e81011f85ef412e9a068204f3eca402f752eb37f53f862bf99d250c37b115c2f8fe3d7cb18371;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd043117ae066cd2062a3e38a5463d93a44e539c39827684bdae7e866629bfe13ddf6d65b703947329daf8ac398bfb98a54fc0c484f9edf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h191b5351737d3e2486da837e14e04839005286fb15eb81da90ee462da637d7fb82d930bee0b13f711385bb08000714ad2cbe3d53d49176e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf95f72e87ac53ca66b08c84423dbf3b524254ff5214f4f99806e53430a401f96e0a69c0fcde5342746ac6080a07e1658b5fef18b9f7bc8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dff1560b48b237600d8dcd7b5468dd719aa65297c2acf659f25584883914b819cdaa31533021c87ce7194ad37d3dcd9b188ee048bcf81;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h152e193674112af017ffbb3f7c1f1261bc6c32ffb3c78905b4af05d0e6265d70e931f1e54d281f12833be02a87f82e6bd895d7f3c8987fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4f00d2115b759d703f9b5a6f4606945a84fce9e87f6b5ed9e2081d5c0e910fbe5d415141b7ebd91330eedde9bf0a30c7b2dc796c228d28;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha41a50096ace94f69d68f7006f1716e714c97460a9ced1fb0869409cb683406627e0ae0bc8683b301d83826c4ef0d25a5c4a0178507c9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1620d141653144edc3187d05a0d4bc0bc1a9321e036a0c4863bf06703612c651207063efcbf93fbff3cf49a71e12c655b14ddd42ee8a0bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cc0e141690c02f66ebb78d5215117b0ac7251a837d686107143f228fad0c0816b3e8d14da8b513e9b4b90f5a6ba02d5999d439c37f5d12;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1da8e8620955107bc3e4ea23f97b6bd04c3aa4b7b79de004d2b477899b40e9df571a6175e6bdec2e6e6980fea9246961d134b4346127fce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h261b0617e316bd3b75dc548dcc63116c240de622abe99e7c9cbb7e669fd27e563d2371299433b6ff6215f53a1e7ebcfd249f9df1fa1eb6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h149e8ef043e66ad7325898bc516089f00520bc0fecb13bd2ccba398ca5100d4d9fc8bdbb044c6380decb7bbe8ef9182b340a5f9fecabbf7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1160ec6d5235060ffb4c3d9656d47064f73900db76de9d236956b4acbb99f4011be31f4fa9ab3ef1789d3be00e9f78e2daae74c44385295;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15c87455958a22a7de2119ed16244270d18bf14575600b3e1a3addeb583f4c897568e8a601e58f74c2445b0e171a5330ff27a2ccef78720;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf3694c269ef459a1c0a67108fd9374cf90e78d7c1a5c67a1529665d8b5d18f9e16572fae2b7229e1b6d3289d06506d04ad4dee68bcc259;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13b9a9681bee9f41fe6f6c145e2a7f912ad302254df49aebde054e22df36018a91592f99c75f51ae956d47570cc8c55adfeac60efbf39eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcb9491de3af9be5b1ec698e2eddff2d767f8bcea3dfa8e67d6350d7ee99c71168ecb23f3327c8a0fb2bc885adf757338625f6afe3883ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18f072b9e3256d73f69ed49c9eff23bb2a8baba1868feb884d207f59ee6fe19a7e3d3a150f88bed1b635668086fe6d37f4916321acf03e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11c57f18ccd06baf3985a814c44552a8d56a7abfe41241219b325c4725a0b644d4363b7a5177c37d8f2a7edae157c9a1d79892a6dd5df84;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c8f5b55d5835c313998a88b7746230eb26412a059a48c0b734aad11afbb5c1666b651c82f4876b47c5933db6ca13a87a9eab84b2152521;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18a85ee52281f39e5422343e67aab9e40244c40f965195e9e731592e655b564cc9bae950f0996cd08979e9ca6518fcf6dfb91670acc730e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13cf98d170cd62eec0f0242e79f66bb3291e89f60f93cd1363b1b4bfd5c9b145a990a5ada335a1d5536eda19f3cb86b73a0d74b9ddd26c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf27263a7e3381cf1b9d5785e27d4955a469000464905bd4427e7cdb1be7671266d6955d77216dc3264ebd08d229fa23585fe660adfd830;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cc51d1dfcadf22ddd4d669b10937f3c014b9d36edee2c5cca8422167876da3b6c39cab4f86dc8b4f0590ccc06804d0ab38ad023a7bbd4c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10a8dc73e7498610fc881ac478bc2130951bc26f24211c9fa550b91e72680f9a3eb4c78fc8ea8d8d8c560fb03aef3f2a48eb4586fea61aa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f2acc37bc4ced016b29aba68ce5a5cdb4c58b2470a349dce1178673eb0f29b9434c0215a88736257969c35e4342c7e682d925addc96191;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h107756e968a3d8d423b8aba9fb75bf00784aa752564325734081a5158da92a108a8dc4d6a427a55a943775a05ae7f1f4d05ea983fc1f34c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h186faaee18d0849b108cc9ed3cfe19061abd33061eff68e4c5f35dfdc2450a5762af7a3ce618f8625b1a427f192b5165ef3c8cc1b60ea54;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h58c8849437e0e8d069b743af5a28d892cca37d610234f6fd9bee09c54fd65f46e368b7a25bb112007fe06b8beb19f4a788849b57b4d4d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c5d0f4dba01a84df970965d75e94bea36174cb4dfc8f305843d7a6d518ce888689e7ac7ac70efa511b9070f00d43404862aff3887961f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18ba27556e50517275783de85d2a7b64a271abcba638931fc5e073661643ae00755ba04437200eadc7d23657e835f04a989d1d6f6cdb4fa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ec71662ab576043961611f9f196e19dbcbaee7461ddc2320f00902481f6443f6fc5a7ba95cb47c86b33c391ad0e911d0c1c8e9f195d3ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f5efd5022d8d267655f826d81d9402f8bf1882dcc3278cca083e5f50e823c3f6c6e39e2925c68d35d27186403a6fce84860a575137529f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h78a745c46de4e950548056c740f28629faeffb43b81b95aaf4309b74e7f0d677a4d7f7d4459ea41acb9c0c863ab787ea010fd9c3001bf3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2cc10dee7ced12af65662a27aaf9a73b9f329958469627c8745d3b938ceebc0ef6d9a5cd6a16db54d7bb6d7e448038e67b315f114f687e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h402fdb65035f2191add067d4c18bc69128f93a3112fa24ce4af1267e39d43703d73ff745dbd964904e99171ba2e7dc36c3614508821b8b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15a51cf7c7a3f743e138ebf2bba048cc7b5b6a8479ece2678469972709eaca1237b8ac70c97c2db2a85287c5fda619bee615fe95f6a1911;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h102e5fd9be587322fa4e89da19396b6dff788512ed58016a0e4445259ad0064e785e62147c32c3d2ca9fb0350c951bb7acc5a0a2f45421f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde06f1205fb0fbfbdc4d6253e2db2f6370bee4213a5244312c9131ee98903b2b1db2ed2c55adf3db92878dbe68a277e12285102c855ed5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b1268de93bce793ee4be3bf1633c411c1955d6b066add7c0cafbc91dd2c8327b2ff21bd80cf6f54817189ef0b53ecd542cc58994c2ec6f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c102e8d3c54f9b037c19c103a0a39b0f201039ba9d2863bee15df7dc548f063b23d110b82b34b56737ce94aa7b933d0e0336d3f877d653;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfb4d651f62bd0fc6e4a4cd9ec835bf1546ac92ae98b6f4ea1bcc3da5021b6b0bdc483fed034622da5bf36b117a86f093a7892601fe6db1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h79de7f360389b08527f7c47fed9a9d1ea0b3889ef569c027619591662170bb1cec56cfd93c4230e2cb54dcdd67f8384e4c16346f956edb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h137131874704f4bb19ccae2b062e92449303eb3a75d2dc23c4ce8a6822a466cdd3bc3f1de3027c18aee048122108f9aabd05700339febed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h149f5b07a163e848ddb93d13351cc7b2fa6f60748cf1e57912de660d40238f994e3b4fcfd1bd5a5656e3db5b30db93a24e0bc9d7ba3d7c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1346f5f70d41bb0043d7f2ca99a43ef1b972b1dc30598c3802bc7bbf2eb900f47bc31980dfb6475ac0b4c1fa0c6d9f5cd5aa88816da4ecb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h427b412aa9dabf5bf4b7329114b47334c25a5b7fafa9f78b5b43ff48b30a60cde07526dcd783aba4a4b2e9c9e7f77935f2cef41946d6e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a579f3a9f8ce911f12b6c5a66b7733ab234277a90102084bcb130b087fff384d7f35ffa348663be890ea0f54f59ecba47614808863b75;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h183a89f1077849c147f976cb9d6099829a5bbfec15c24b183c87d8efd530b1ca2a49931dd8b7ce9428e9581585642e6e13403e68f291d43;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e5ab269a531d96ec1bb1695c197a5864e6e397706564acdd606312563538ae918633eeedef767392cb5dadae15bcfc80547b46a2f7bcaf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h104b794e8d52e97991b30a0b7b278bcae542f749b604677967ecfa0486005bf75d6c8eb6918c99679dded88e91daf102e4206e2be50b42b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17a32d8bd24050476ca90183b4c642fa2939cbfd01a3e346efaba86ed42e91c98ae6e35537536aebd918fbd894c602c8acc14a5f3cac207;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h185b9283491a63913c0fcffe75e15f9bcddd5bd69e0f659c66bdd6ece96af5da7010fb7f47bbf0df04eb0db7266c4534a1047a9200bbc89;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h23833be86c21005056c92ec49cbc4da055edd5036260205dca54f9b5496c5f4728d422c1f737a8cc26929c2ba0429593ef58fdc7142b42;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h74ac5e319080e2d981d0ef10f16a0a858cbb7cff296b2d10543d3e0fa500f03424e68169f06f71b6d5eb3fa53c465a99b30232df3659bc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h59b27d924bbe57a45512c38db53bfadf3b28ccd0b902ac5f0eb56d5adb97382d3f9ee42e4d104e76b92bd06bb85d5d87477226d460ae1a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb7f42d02d1376f911b7da7b5206eb9e71e892fbf7c48f84ef8cf0072a4eb50a9ea8b019827c5e4da85662da6962d2964cd4b97e482d4f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hff5f818a011abf8cbfe71bcb2d2c43ba2446da5f67369ba74003f6a2419d49cfc3979e0a18eccc164d267d08623e727072e7a0ef2eda9f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19fc97b02703232a14d732f5aed46641b2a2173f38325deba980d2351444fedbbc15c2790bec4b83614b26f8566b7f01c59c94a4a5d61fd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'haf7bd5e0f9510e28fca5e82ef0884657827723499d989a700713a9f0709c284c1a713afb936f323fd73ae8e4d0a6104ad7914ee6d64b0f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he86bd37c6eae3c5d4def66e553e6fd3052a5be9b55c8eea5c683f808930558a797e66d92ab4288e3f8864a9d946aaff387a2bdeba776e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hafb4c3e056e5026290955f573f77dbb762f800e439e53068ce725f82b1b9011672dc8f9979de83d2e09a91f7c82d478f0fa10b31b1a799;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1080b42710792701d0b71e0e6a86d048c393b385781a46028cbb8c20d45c3cdfbd44935c680821bf9424a55f81bc94d3e7dbd0078a3ed91;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he17e3ab8dc31f1bdf98b69850c4999e6f2a73290358c02112c91fdc018a46ee0f0aecf1affa894b3a3afd1f1fb7665664d90c1afb20ab4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15a339df99564450620aed6aa216c1e948253e0d6e50b0455a91291cafa4c107aca8b33538d11f1e19ce81815123082455350a01013c77a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ea6544458e2c6e5e3d989ed76dd82ca1441e9e07f71f3d701537090fd3b6f244b51144b1fa1973c8d805248b20b8420f487798d2e61542;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h96a28ef62d66cb2fb8fda908f9ee9f326c0d4a318d8cedffdd8db1201f4ec7566d71e921a0eea3035453c65cee02350091411b4e2c0ff1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ba9cd4262ad4e0c9658c691674f3f7c72edc7cbcf6271ef454e2eedc40518e5b044cdd66ef6bdc1ff350a400746fc67a48a814d516d09f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cc7ba6a26e5afb4a5b59a1d97404c571b65fd681c24e3b7adeece7193ec8715de2701aec95d0b6df0cda0ee8dbe8cae2a993083eee0d50;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h358d4c14ba1566de95e1665388959c2d119a846371118fa71e37bb15b8592d2fe95adba458c548acbc9df0e5be18322242c6eaf75079d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h26dd2f791cba6bc95b425b7409a6a427ba3f84cd869571cac5c65dc9e4f84c9fd2d151d5e45c7c284c24b84802ef1080820e35ff2cdb62;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bef92ce70e02bc2a2f804b4c60523cd757270e3d507db3e667caa14184411f17a731feed1468f0e531e92968c6ad9689e8926303a5823;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h45249335c0701876834a60396ca60d3fc4ec500b8995d505d1ea05ad7cb2f41627d859fe112107af52ab41fa771465627097657382d5da;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'habf0161b065bb2cde8423ac79d752a8b0667eb151d5ae5a5a8a21e1ec7aec8b8c262b012a78a713fae3719992da1d9eaafeb31cfa77a9e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h347df6f4b0fb433a8246f462a8403cb1a1f7536cfb35c66bdd23a77263cb64f177e578ba922ae88d06bb5b01c926816148d98d1dcfbcc0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dfc5bd898ac51a8b844e6e798d38bbdc2013ef3ba16dcbf6a91dafbe88af244014af5ea7924d978bd7d9fd4fb20be2740e5a8ecbb171e7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h116e0bf11dbd6d9cb803eb9ea4a81cddaac0aa51fb3cf70361969319f3fc54bda826ce1962dfd27ebfc363fefed86415f1976df828adf94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc1877ac58fbcf5b531ee1610a897a0510d4b74655197820f9739c80c2927f59c3633fd2e2e7a9bc7e30338874aac373f956fe14d4d7ae3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he8d74c6f07bef067f679b194fcc57ab976d8de20a20b1e6e413d5d378bce9da444b9db20faefc343d3c6af48d409586eecfeba75815faf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b5c30ea261c86391b47d5fffbdc778e487f8eaae35273aaf25b352b603dd5886448e2d2d5fc4d0dde3b8f2ae596e55f0fa7e0ea0c2ea9d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hafa0b80c1b1b0c2eee9455a28baf66aaf1ad40acf698656ac890100c025df53c29bbd5f181cfcb90b1c746aa37bcc317a2f0456580fa1f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17109fd537c2b84ca1a03382f2945c5590dccecf9c9f40d53f644decf67d0bf28fbf6694323b22993339b74228ecc9a12b0fe86d73fa042;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf28a05d04f4f449d2712ea5cfbaa4b6c4af8d314384ecd062431b893916fec760b7f5481895afb6ef0706101bb7238151dd684fc6bfa0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h149c5dca8cc20e35483e61e6bf92f97ffafb9aed7075454be0008c0545c9f24d164831c131625e1023b211f382496e3f6aaac0b4090f7ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fbb586d06643f783bffd6e80315ff96845a6b931665fde05e06c489ac346f085be42d7e888944f3088471e95c44910157ed4f1fe707e25;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14968d9e3413452d67cbab008a63250109d84d0e271a8b84c6a09be8cfe31533a52fd6e137e68455750ddc924684196c53a2efb0ee41d31;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b798a5c7978344f1641c8c935b2110904a18526b22777a79ca0dad97512fbe76d2b6a176e1628ec33ba70d3bd2aabd73e477306dff61b1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c712e82f838693b12a4cd9ceaf582f57aa48dbafdea32bf43d1d065eb50e22c780554b21c44eb8a868c3eedc3d3a4bb659ca299eafe53e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h78b3930286e692d9266c6a36028f13dd64ad42a93d12272048bd6927866cfacebe03ef6ac5fd89b3b9842fb3cf6504f2a7f60feeaa1c25;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4ad10652528bec857dff4f00e02ff8d192fa5a39f7f0aa26ee9a1f73f0ce657df95b2ebc768e5c91fac03544a70b42158b639652972e97;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he04a8d9cb4b8111ba3eba26a6a7ab60699c1159e083f02ba3203c03db9cb3c4858031da750e8f8397e7607a6ba68a82c08caf80ae15f6f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11c500b0d9f7cfeb9b4eada2557cea7e5323810d08832bc28a7216a0bcc4e8a0ca6456694c5b6b93764ff1f8ddd71e0a11fcae59ca6186d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h36919b901b47b64259aeff0c13f27e83b7546df13d43f524e7840aaa01299e82aeaf6f2af139e6a74a29bd5d63fcd93791743b19e95464;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heea853d276e6e104259d6bc430c78f05326e5c2bd95b808839dc69de7ada7fae9451818d9edbe315e45708689aefc0ef876ca8ccf3cc60;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7a6d376fab9865094b845f71e0a5a51e2441dbe613f1b8197f9e530c16f505e2f456ce46fb8eba94e6e9634cd201536fa198f5f0427f97;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16a56e51e091a7e917f39d1003b847c543263111ce94b2b3432c5eebca77f69d26d34009af6f244e027325f293bf508f9194243f32b51b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2d545802b6566b74d30e746df1c94767a7a387920c54558900be3634088391b33e46c64af77b00911fba5d6d6d0e19f5d71959889387d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13b715ae54be7929f90f6d437c8aee337c28e1130b69160f37ce90011c0e62f008a1bac0adc75f8435d847e702f4e0cf4abc3ff0d1119af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4fd293e55a6c2fb92cfaf65266af4d3c8b5f33bdb45b93587713735a9d858dd09458ae64cff42a1854656122c4faa4c7d6254a5bf3a163;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16f7b5093f138c09895e5edadf4e317abfb019324b14ee656e86160a932b5c5faac4380933124a08ac36fd14463b7cec1bba34a9071ad5d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19617885a796438d3361cfac4308c2073d0d2cbac70c8790fab68c8e30354e79cbc2517bb0305d22ecd7345be9e497bf44df205cf79099e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c9c85c49e10c1e443e473345c354ffe990be6a05a96e2f96de0f53dfb395e49a82af242aff0686f93cbd694cc63aaf1fbb094d9ad5d17b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2c6da3dcf2b45d5f2b8cf1ed4699f80ebc387d78e5320854b38445636e1529ed6fe3f7a668d9576a02a02f7bc7d845ae117146e987ade2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'had5fe846562f22bb6c1d10f1727bbd6bf84d41feaa4319b54a02f19d9e2ae89aca979e4a4524a133d9b37df3c1d859ae2b245892ab200a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cc49ff196bbfe80d79fe5a0b126313a35da230b4251e04e7c4343eb74fa33713c0c2423902c7153c354ebd7d747ce81f2e9e4c45d132d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf029fd5b776fd94a3100b1ef9795fe5a341d7130864e5d7fb1faf11d95d471aa869639196eb32709c27b84e6f028ab0649c48b9fde82e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h199149c5a575d0cd3c16ad70d320d3d6cbdeaef6455c2bc1a9c1d91c19b6c3b4b7c064cfa62539d9efd5b9e9ae8166d0de3f942cfa01428;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a4005fc934b5a94909fa462257ff1c2de73586972ae5a78d380235e10b1134903409aba80295eb07c580fc915b010c037076b40357e713;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h103e9a1a4c797c1a8bd9dff7d69dd985ef3c279e2a655c106b95991ada586cd2ab140737cd8b9066531d9c52602f847c1e81ea2660a96ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6a4aeebd178cbd10c62d8d062cc8869f45636186d25dc8e3a281511da2d0cab708ae27f781ca8278e1d675a325140c26d32718e8de508e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c35d66f99ca7251b28a2d86f4d0aab411b4b54abeb037c42d749690eceb0868144bbc9df1bf2d8b17d60805879f7fa022ca1fd777ba48e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8965c35935dd0fc2b6144c9cbbd80bdd838b48b511b8af45dcc0685f6661ddde6d9f08c9894365d119b8a1bcbfc88a5f7e6823cb7b1c5e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14f712d47407cfa88efb8e5aceed82b231c07a3c424eb73808ff219b6c80cd9b3fa049b750dac197e91af3b0430833603ef331499940525;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16d268364c28b918fded8be51894db16e1af22e398341c023702109381a237929a606cf85dc50adc6313032b72ba2da5cd1bd84a2ba17b1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11f63b442cf9cbee2d5210e2ec8c4a807c6c853b53097f2f358edf7b04ffbfe859bd4625134cb295bd143e954775aba79bd33fd714cfb18;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2cb0106537fa6af8054b0d88cd43fb3e861785ab995c5f09e6dd8fd561c849300af868cd194b61c74d9eb053daabf829d3aafb3158e604;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cbb77e66ac7f42c2963ea5c347b8b9e35de4ddccc58e65d74c781b9d6d33d2be34b23f123c29db0496101d4b189d7d4b9a707ec519594d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cbf9db8ab8a70cf9359949075a2aa7307e8fd92b36e0d26d546b010c16b56af95257882a884e2fe5ce96efdd787b3c889bbec757f83caf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9cb985d89962a9f14bb39877c592ba0fee867dfded4637ed0a0b0c2a04349cdce6c175c24d4ea2a7582835d9222575a6341f01445dd0b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h101a746084a0913485059a4d50dc6b9e4026d10bfa0b3708266442ca8265016e74c9cf437f346585fbe4265e4520f49fdd4399f7cb8e09f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14a940d462e19aad310453ef1d27210f77267b8845613f9cac534fcef17d1ef2ce1cdcc4b801e0108b903a677f1fc1a8b031efaee3bf941;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h149854c9b9f50e59538fb2c650a752b9988bae4e956cd9146867286e834be7be802e3ec0452ccbad189f6dee11dbd2a96db922f7fa42788;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11b29f9f8b82d7ea9c9d2abbadf264fa44bfcf86392d9d0858ecc06a5dcf9bd32c5a65ee2bcbaa20a1f0fc65829d34847609bf9dacd21e5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ec3ff107ab1633291a90ce13ce86462b3bf16abbbe568dfc7b512db81e401e0343a75ed473616a84032b1f08349b56d12edf9e38955371;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3a6e4782d5912eb8792af5cf2f86d9071bd2e53b98e5b49fa29ea7d882c2d49b967fcc3f80d42554cb05f87cd8ba77c5f16effbe85547;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h97a7dffa9bec63b8f24558986d7a64b662135251bbf1067b67e61be86828c80d5d63dba7f41084faa2f94508e8db14c68453d3ce7acb8b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bd1dcd7c4f90c351850a723d8528cd59a8b4976b4b4e689e8cdaae98fd640c129ef6c9b526cf21feea3a081d199903a63e737f93f229ad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcaeb52854ab903897dbf9ee04c8a872f44d5a8bfa2592a722f430e7d5cdc5aa5e83890e10b81bb0ade4255eda0a7714f72bd49dbc6e813;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1701d14851b04711a0ae612bd1e88cc68e1e37692de143e7be2907ae36532becf40d46ccf0140f05dcbe910c4eaecb0d70a431c7aa4bb39;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1272f077830e76cb3895177350e8e601de4aa2cf65f125e59e0e128acf07ec040097ad4d7f3a22e2a805c0c87b1b48c2e8d8fbd484fdadd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bc460c7958be1c2d30400e6606faaaf38da3bccb83e96e5592cecd12d209f86547e4fd2d5c641f0143f7aefd161627e3c1f50fc2236f35;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcea8017726347d8c5ff5b090659afb1c4e4bb61b1c7759f31d05d10a7880c5ddb70d708279c46c191c561770f9bab512b1023faf932438;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10014b03b6827b539e26843c4476fdb39e1574054beb2fbeaaf300eecac082b48a1afdfd82310beaaf8382ea8cab1bd4424adc00669e7c7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bb15fed36cca644841487bb0f7d3c02369e1c0255e8ee507a3e7ad1ac9371039abe8f4e4e9c358ba2fccb92f0e5852b8211d52cf92c79a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h60618494a320383ba58719f7825c5b484b282825252187d6da8df3eb44c17b3376ed5c7c6116aecfff6838329f80515bbbab7b64f2c764;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b70f742786f4fbf86a0c6f78b534d4ef6f1dcfcbd2f71e451c26dca14722f772184ccfbe171946cd89bc76d47dc6918765af81084157b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d2dde78aa235aad04c4b2d80442d04b15fd2254caa4b906ebcd52505c042c1a5d6213597a053d022ebfb3870c86872072c41cb6312477d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b33f0dc243dc98b74bcd627f167591b8cdb9a5257425b1dff0547fae30b6d04ca1fcad450ea78049be94f25907aa06a83ee1fd7f438c1a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1201f7a1611ca640f98b9fcf0abb142bdf66486e3be56f7ce21c5f355d58cb99df541917d98795559a635cdd7438c7462de919d97a08fe4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h638c41a401dd0ea189adedee7e9c059bf4fcfb15689e1fec5ed38174ae67bf4bcc29b7e72e02e835db4d8ffe605818c98583ad33d2372e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e83304c9d6bb64dbd2a6abd1cb08e4c383bf74b588b1ac5e6ebe9e906edd1cdcea4b52b3edb335ccdd290bc44c60c93d95232b1050f87a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11c6ccc27c675bb4d2a3a69f3788ad70918cd163e0323f09a70232e9dc7f06e3fb73392b02a0d0ed4afbb47c68c9593d7f9a3c4c131f2f0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15387e98b66cef0d313c9e1e949afd78dde4513571fb6a3028204a226967f5f00ae2409cf6350e1227e8883c38a8f13864240fe16f5e843;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2c066184db2032810a2423dff2b6cc5bd08acfb6db2261eb43fa9f8d4bde80ee9e272027d54947c7becc3825450144ccd3e7664854da1e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc6c0fba6e47298ec84a2c27465887a7c5c306a06b456316dbaa6cf056a0da5f62993f6f049d36d8fd7f973951e681db3e5ce5cde9326b8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16146ae1caf03871283b121ff5f2430b790f051fc64ae823b18165c5ec45325996db66e58cf283a1635ab88e4dd3a47e9b466fdb535d95d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h919987d21afcd68bcde9f8d944f8cce001fdbf0566cdcea0aa56f9854df8c4989a1492f0c61f6b0ae105cc0604256f3fa397e37bda9120;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9469c237222cd912859ee672b2d2cdbe9db3024f59aedadce8bbe20b78a6f912ad732056748c6e407c1bc5d626dfc9a0dec4792b0038ff;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1affeb0349cb202409769a086f73cfe2b21b79b13816a95ff9c9c5b833ceaa02eaac93b3b65332a1b55ebf681d5b3df2d9f04ab29b785f4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16180714b430aea347edc3b5bed89a2f8d1d79b3561a1037da4bd0078c3d62bdadffa0f3ec48f6a5abb3e15a1088c8f4468b3f8ae11396c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f0df8c17737d668e83755c6b9df9548ebe8e59d259cb1273b29c5466fc8b85d152ea3a9a521fbe6670b17871cae2ad9e31750b72aaa2a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h163e4fec6d4ff2d10e891302559354a2aa749d6d606fa6d564e0762eb32a35697dc8b650c6bd3e3c3c66dac95b5e555c5ed1b7f351c254;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1acef5895dc5c780cc73f3ffaf2ae5531cc0c8bfdae0a7a3658248741b8eca85232200cdc8ce25ce86419bd3c0815554fbac09543d2178d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h563785c6e1c189b4a2b589da278d00bf4e0257fc471630101802bf6d399fafd25ac69c5602cbcf867184720f5ed1fa83b1886ef7effd43;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6fea642e184439d38ae6b5d872af8809d7424e7ab955d0cc223c24254cc9f9fb1654deb5857e01cb028cfaa67d5a999c6b84c36b946039;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12ec8322a21b9c76281270d09074e723f14218995a57c2f703e8c10465556cbc2091b698414f79579582013ae31156a0124948d2ed78ad6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3f9c7bd72b31c726f55a677e26da71e4eebd80168fe69854dcdb1971d78b57b1a3c088cb29454a8c09dd9e5dc999de4ec3c93e2db8fd30;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7996f4f9bef9e96e047b26052e441ca377b1a58867dc530e0c32084726e6468acc8a5c4f4286985e4069f319884e78ccc06fb47dc59b94;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h103c665367e4f62d1742f0aeb0e4404bd11d421dc0a1d7319177c55165000eb8424a0e19de6e564a2a9714b40bd31b966014c7f615c87e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18c6a1f12d7e5d9ae644c1fe9919bfcd6884ea16ec7919dd2dabdd98d701fb9d11bf548c284ce7a615bb03f1fd0069ab683d7d6cb74f89e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2af29ce1489121474d48ba92291e7781df1571fe2cdd1a56c59e97a604760bb6e1644c2b189ca1b460a4cc18ad019decf2d3a91a869688;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11ad0ff1aad1bf534279290cc945244cf1718d54bff3dc887d205aee059b38b4699fe6a4519c1bb26bbadc577ae489dd62f8a7370832260;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b8f4db7f62d1e5e51e8d62c7e8f74ccc8c4efa6f83dcf78a2ba2c55b9015259c5febf625d3374356e191aea7ab75c6589529edaf6c8f72;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6cae4f9ed800f42e1d58058af39936ff52b2f43102e4972e0323555efdb0bbad51d8a76b6350bc5d39a23311aaab99e865c08cbf158dcf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1815c8d26eb1eafae155ac397bf9dcf5de85d92bc3795afb3338e9d7983ce4c0df48e4043126728ffe21b7c5bfb50c60797b8e9a7bdb13;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12eebc224d44c9ec9a52527db13b1d0c73760758124249b249f1feca741a22eae07902e4e5e9bd8aa4339745d484b2e99aebe9c43401e2e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9997dc0bbba327a8492ce769456d5cf35274324519fba85d5378036c101ddf2b5e80a4e6a9540e254e9ddb7d10695cb858e45954fd0ce9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18b7216e4603788539d7ee5f7ad82353b1939d6dc748b9714af4223cfee5df8be95c2b000eff098ce9583390c0f7563fa9ec7aed6335ef3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ecb3bcf205166cf5fabf6e59ca0a2d65e9132202be9b0eb1fc97e1a213c35ffdce66cae8d7d36216685721678674fb0fb9300ccea4c27;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcaf2c162d970ccfa68bc40ad22f5dfe90895b75da5eed2accd9f5f6f48ea54e9b16883ddd20bb7d0dbf8176f268564de3b7d5b7043ffc9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha2bfd20bd1169a95da917848023bc4369d34f126d89ebc88d0ebb4f55f509ae5c6c30d93b0ddfc0f3f2a71196365a63e39f188e1e74336;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc573e883b5077a36aae0a75e7f9ce992e50c9572ec8b79d54d5997706cb226f4c992b86a5570c324166e9f46cdab4ad9fc61fca476ef8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14b4e64c7da1d1363fe8f93b5e39e5aedc706a830d4aef3c6ebc7ef4f737d489e5771aa3b1bf8de38403acbbddf01b6c8565d07cac8f27d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h272c7c4afc2e2a82145c8868fa98f6eb14fe88a62692f011dcb885f95ea1920127b727d748b965227ebc89b460663ca3e50bf0183e3873;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12e49d37885d2be35177547cd17f402a5fbfc829c3e6c72e1164feb3e494c928dc503c950363cd3f83beeb85590e264623e48886660347a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fe5d9598d6830cafa8426953f830eed3630da2a190e8744da0b78ce8baf06fe67d77f825193a04286138128d817c1b128d76ac0fd8a885;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3df7fbedd82db35bf39e8a3363ed463ad0fd116c8c673935672ae84ba667996d016384e2b9af2ce6f9754f1bebb67de3e9df004ed4f83;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12bb1ce10d82cad410a76f8dd28781e71af5cecb0e086a1e755c8ab261e7821a4840fcd4590149b02266e4730f15dae1c19b0217c2670d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h137a33a0cd2c3d5dcd3e01f40811c684188814276f74a58dabc5e21554a916784dcd45396e04b56890c809ea880587db2451589afd70424;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcac4cbb239235cc607934c7f1efb0a437229254204d525dc09a360805ea8cf6403c91b9187a995e872c952886bd2b23b7331b12e0491a0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16054fba8ceb03525a1ca7ed9579890d5622c3d9bff81c3b0be90b62198464dccf1dcb82e6274a4bc3b2b5b4627bb6fc86a76ed987ade3d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10e7b726f52cbb0388ae8aac61ae62a68c754a7062aa08a9075251380932876ea7552afd4973e2ec0a263b69e04bcbb865ce5e432d61d57;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hada63cb46048523ca50ab40f54861a73680f61730e9e5fc4073d1ec3e3edd6cb75908e8997ac4e93d5e163f97037286a491f0f0d74f870;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e64317658b575c23fa2f9e56cbc67c27e072c9b7b4e4bfec9dd17282e3e66e668b85e35187a521e21b2bae482b7a438a879b366c1eef16;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc5cf6a8060dcc16963bf4ec11f0adb9e2554e4b7700b1b8c7f2b74e7e98bd6343f15109d9f2b03f5543d364478d478276dffe09fdb6adb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13adaac447c4e8eef2f1a12fc9c92db177dc45635f4ebd90c20a51ebafda534b1c4de7675d5ebd6d3b7acdb1f49a6b6674e4c15b4f24220;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf483d22633626f878fc36fac45912d2d1962e393846e1d92da39c24d35c055157c6b1012221ea27abe78758c9f77c835d658d7473400;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h43b809c881a63b406149f67cb1514b23d35cdd9a00d235d2992908b2723e5b90260a2aed6939f9325e55293fa5427430d227c95af2455c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a5d1a65e089c521dc38bb4ce4b098ba415d456197da531d6b430201a0b447908a8a7328277fa1bd4291db75931b3215dc419b016a410f8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2ff2a238a15886a04172a854e21a91d6d1d3456b9bdd6bb2dda457568bf6b1c91a80b5b3b4406e0bd392d6392d6eccbb511af38849309;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha038cdca6aa9176f6c0649e67e8d716cf84fa7f6aab8dc6a40af4f4b717a3456c167fff3feb94e049ab5b01f039876dc2a5e2a9614fe8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h105a404c68dd958d284d82b2d5dc905d774503b2666891c8a595ba97f43a9fc80f4f5eeabb00884ab8dc7b2bcfbed10401aaaa4915f119d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6adf2cfe5e6185742792393f3ae3ce75e47ee43e09848984516b8e602f16ac92162c7deceffc19ab81af265e21ec638498af788f2a31d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he279a12e642308c1d6543c14cd893768e702904bda5196531c04a3eacdc7e63716ea2cf3b049c1e83a292e17969995e34a9221edb00cd0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h79de6a48ee511db15953f765c7690b7557b541a8656540fc3c88f713212f09542f664460ff7fcf14aded63281334dd65962f1cd170097f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3329f8e9f341f0df4c6bb1f167e230064ec4480255d68406dd7fdf554a5b8f7637e8d5c4e548900f1d3c44af0ee301243e7be398ca37ba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1458828b917b61dfe52dc770b607c94cc43fdb3b17372b76c3c9eb0529867ae45d4d04f7e74fb202402d0703e39b6fb8333cbff3c1b4da8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c7e622c13e285ae8a1bcb73a0fbb9acc48dbc72b11632cc6cad3d69e7c88f6ad1e2044a3f20f3fefd3ec929777436e0df1b7222af83dde;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he9acaf57ceac3103fdf6d5627006e7afd2425de15acb595171e7aab91b942cdcc329af526df88f71fd4d010334001c15368fe867e84bc4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h129ab2f7e8d34e9f6428caed29b3652d72f1f792b4ad92f6b723ffe5c6a9d047fbe02e16a6977a4c600a4b150d13eac804e4b1f99a06e44;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17b5a75642f811de9d0f0cecd3f65265148c5f7836963a580307c5702c9e6a91752c6d598641a2cfa498b4a4f61babb436da14142ca858d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h59518e6cd5eb679f24e8c4fc2ba3c29c93a26cfe0f9cd6169668c648923983cdf22a19521b3e21f85c9110dc397a54d40dcdfdcc55477f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h27f717d33a51d6148a5ef5e0aafa0d9a36689428472ace9dd1da6e03dc93512cd92b4146679aa51d4c08acff2e89ccebc6a808e251a7c3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16896805b394d50c2bdc691a594590cbe631436d3630dcfb213f5db76b07f4c8db81a988ff1aa387a84eaf15fe2549d44da2988120e36ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h180794d6070c152f91b05a5a5c8c53270556add9f28198f5c8e9fa46423a89afda41d993eb429cf54c13e24171288885976c80be1173944;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a919538583c50a9d649510db1edec829e9c845cad90bc26cb14c60d444693d8cb69d7e4ec17117daa4e13815fe6300129811f5e53116c7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h49e57905f5e2223bb53a5804aebc665e3c57a41b7bc6d74867dbcf415bc4668e818fe2c95674a3504812713fbb9aa7ecdf38a61092d345;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b399e5eedb45832410e0cd20ad5405572f5662f9e3faea12115a1aad4231f3b1f4affbfd6788cb6b9bab61a31ab01666b4f8447188618d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10742eb42fae6ccbebed70458655c0bdf8dcdb45d6ba745faf10c70074e85284cb0ca49dd6dff538485094e50c1fa4369f09999c315073e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b605db867c990d9acccee91308c37b2b3de129683bb120e00012cef22b114ebf849ea8927df2e7d945a4d9293affcd1d7ae0aad869a329;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h46815556f12f7951b95e25a5d8f7c5a3daf333a8859cf1b43bfb5ebaf8a72c67d10fe1aa6c0afa3bb2db21b08d700e40d619681dd0838a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h100d9337d0fbe23b0a8720463cdd3c79219fc248988255e0c172799da3695e082be5001b405833a2d185fccc60df02d4c021f5d3e24c125;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h766635845f241f8117a64f15d526ee30c8698aa55776ad2ebefb3fabefbdbefdbe9efaf7e5f2698df19d6d07f3a1dc456f4008b064c3f2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d2e8be9bdd6afbcb12c6481a9e8e1b10a91474a3fb904e976633d4bd8880b83bb78de82c8f26eb5bc731d71801c7335bee3351f6b519d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17453bb1ab4039f1684dfe5ffd93af8f20af4575e18e1f0b0e041bde2e1db190d00e77cadcfe758bd19a8c50eeaf15f96af0a629a5ad32b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a43301e24e5400d199f986adc2767489012a8d629f73cba71c23a460b9719d914e768f12cb6e3b9ad96d30155ea1e03bf98adb1059faba;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ca214357bfea6f271746a97a01ccf5c36a0a4869019e95988583d5fa4bd42cca8a69fd1d229e5f22b6f432782bca601be54857bee2551;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13aa5d9b5b068ac4c999c147c58cd5eeb105dc5f3932dca68bac3cd919dfc7de501f2bfe952ecf77feecdeaa4cb5a721e8ab22256d6f27e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ac0cee3f21faf1dd8eaac92076f4c32f1a53a9e128f59fe004f599db545900acff2ca2daf19267f0074d7a61833eb9b21af148ddd2bb84;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha7e43abb8419fc8bb21d5d31bbab340aacad5939d7bf043b1f246fb865e72433b28d1d77bf9856308f0fea3c15ed33132807c7c0b9bcd0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17893d8cf893c7d6a00dd7d63b904057740382f80a951cf76a12f7b5ed9cbf8338684aea0d3324843066813ba2fdecd2865f1836eb659d1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbada613c88f15b3f51bd74c1d5a147b487cbe520f0550715ce25ae870c5dc433aa8afd4fd959be60ac43909667a3a4e5ba0abd418981d7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16380cadeb962e8fe57b28d0d11ff182a0aad7f8c8626600b8158590ea9aea8637f187909afa52cc600a5ad2b8e9ea0e404d55c8af81a96;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ae8ee108a29f7d5ad24ee1ce926296beceffab5f3f4ede8ca5c0b404c385384cbb869791b04e00af6738dbfdf786b99d24b6347608d8ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16e7f18eaaab8e17d3573d69590577b96b8e5b30c53148f4eeb3271ff673aadb42579fcd6909f37e15cf1b777a09eefdcd4468cef7c84;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18675d39bf3c978699dd463d78edd1ae43a2165e0cad072e97ff7205ca54ff15ffa0199e8f988ffff81d5e36249dafe137af5dd9e874fe4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8f1785838f6dbf33060d00673f01a33d8ab686193ef29528843ea607679f344111b56e3be59a4532815e39a59b5476b09274ac3725e8cf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c16066c41157c51f29f0f736827aafbfc08ed22eeb7c08b9cadf8ed7f0591f5a0b952f9ad2d7bd30f9f6ce5e3edb88b6bc520601653903;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b73f595808b6fab5f863f233b8a99f4fdbd7a0d0990b121855fdc0603ef57e98156b89dc4ef8780a6aaab26a838b809b41bf6fd0cfa1ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10438b3b771a5d81235fdf617606d349228574ef67635a7961b50d881589eb19518c160c1a110fa42134ba92b96a8f59aecb6b6e429b0af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h133a3c0dcf1ff7119b3456bbeb8a4008e8a31f0d531b7d87a28389e46789edb41d3cfc929ecb309b4aa0565b4cf04d5a65c6921f087127b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h198a30b6cafd73f0f006b5b07c774c0829b835bbef0843a3dcaaa79f24604ccf1c59515d5fcc95a1b2658c1402f9d01519380f4aca2cab3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14051d9427bd36ea6716e7678d1c6580831e9a965e79c015bceba26eb11e37aecc6684085a6d970c06ca0b2cf79db9acedaa74ab7165a7b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1175ac48635a7cee06bf884064250727fec1cd638f6289d58f60be961a2f1ca13e80dd6292372e32f037b996a62658806bf5cbebab132db;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'heca4928e62ee45019433a6bdd6372fc7af9b1f9780ee62b123f0d3d7c880fd6f512c00e9ea86d3a615d633e288e5bb6dcca4e685588c4c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h95aab20806182c9ae09c04cc4f61361d39dd3d3c82e824889b2018bea1ba9263d99e872c5622134f7a754985db98bab6a9d6b58a1600ae;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb647d33aef4af2a6abff054636cc4e3b22aa24f9219598a7ad1b0e5fd553edf43498dc098517fcd617712acb060276f9f8aec9492e2af1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c0de7818350965eec56473cf82f9ba9cbdcc9abf6008d2dd67b9af2f52266769c97bf53eac10af2ff51d3b5210715e61e61c7b977500fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha15617efa1f7647e5d510312e2812dde68616348373c2445f902af0e7f10a42d00db6a9df262d1775f39b98261f2efbd062141b880ef7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h121372c29b50eda35b161444c5bf7665482f7a1a748e742c1b1e8dba471fe283a0fd0ecc505ccff5352623958cc3e35c3d88d4b65fe5e68;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h71eb692b1d1889bf69f15e5a617b9948efc6afb62f263a00918e1eb8ebc99e445ca85e81f1cfe0e99f1165745a626c36e9bfed0e0e649;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5f48d5117ccdebe829ceeabccb3c3899c4346712179d93f5b6bb5a08ce4f21408b724a4acfd69145ee20363c8395a35def0c8defe117c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h116f2405a77aec9747a3852054ae213dca28fab602608577386f283035f855b1125776be4e58fdb7245ba8dec248b25af12d70a0decbb0b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b254bb4c8d8d71f5868a55fc0ab91de3bcfcffbe2a0209d56216627734bc611958c80b25068b92aa4c88985e99c351d5b0d5dda296435e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h21be761f3ce286a67ae82baa2660ae19f722a72333d1a4f5b12fbbafc783360feede5ac3b4a9d90c3f10427ceb9838447438276131e41f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he0521cf8165002d9afc09fa5e7e77d7518415dfaa64d0829989118efaf7ff1c84f6f92c8aa052b044b785ef5ad28f4ccd1bb348b9feaaf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb823557fff812d5a3500cf732b1dc759d854baa0878496f56450871ebb7f8fe5d5a468fa6f9d270a69c84a46823c7762589dfe4e059a09;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd1b8bbe8bae3ae24e7d37a870503be08b71226284d6fb346917bc915e7d19c14fb77eff1014d082fe84546716b95e0b43f87304e70492a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h198ccfdf6a4f4e78a737e719c573ca33b5f418e4eceb1023e64644aeb6c314d2295f071fba8918b338d6ac3ab045820e1d26a82c3912d0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h60d348cb57431f7a63ff4395393f335e979160debd7e721167643e6d797c11f90c1df5efaff3122a9edd28062a062b35c5cff3cbd33f88;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2e8d9529518868b5bb6b145014b2121632236c7663b54c6320386eb79854535af6cbc6002c6eaca2fd22ebbf37879b62708e538d567b4e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc65e45c78976aad89a0dc3d2b83c86aa1bcd1282c102367154eae9ba5fbae757678a0b68c9cc700662f1b0b36670f94f9b444c57bff95;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h135454da23c5395a297c7c47d673c9cbc3b8a75449a87ac69d2ddadb58141d4732e6a59176b4d411fda0a07759589e6fa0461856cb6fbd3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4640759b2ad82b163a363affdcc7c15685cb880c1a6b5d4bc371b5b386f5d74a06038f9acc38fd97fbe284ee123dc924e6093a48efd1b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h194c887a1fef76588296b081c18934f8c89c1cd665239037fd15e45ff71fd4743577abecabf1afa713e04bd83fa4d4c906df388c150cb99;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5024bcfa5b07237b453824680991a2d82f912dfe0da7e569526ce804d9f49f700882ebcc6c572fae53e5a358064ae17af58c60ccbefe70;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16ff4d10562eb3ba1ea7429df003c6e482204253682fc50d27eff8e6024a0971a01d7d8ba577c6b436ecb5ffc3838a06c2a88eb8ccfafea;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf298fce9c7b049cfa02f58717f8261e2ebb502759544ddd18fb2e0cc5c86435b73a303f618cc386882fac613b003d507e374b0c62cff0a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d6c84ff70dd1694c9c219e1e08842b7a55d1575716adfa205bc2de0cd64833629990831e1efc2de10fc1daadd1c6bc50c11c494697d744;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1a4a972651a157527251167bf4392bc80e558292a6a2a05e13df84f77004882bed929cb4f20ea79c08ce7b0c502e1f058e94d862ca42734;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d303fd94306aa76e2e716e008820caf7886362ecf739ea871c5cd36abc8273febee75b77bf6db322c11be6b54565a326223944294e78ce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha523a985d3e13487bd38048c846c211bcf16f1a8bdc71d4384d0e7e72256dc9dbbc0093746e0dc58c6e3312fc20d67212872f9d3864568;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13ea2878fbc57c1bf719272578e4f23360ad8027460d8ff5d79cd44d135db17f5465ae09ad1579daf82c61c5b568f16daf1e86b94ce57a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h42be80923349f7e7b74788dcd1c555d964e1f06fbcaa492e0f613e6d49af7f288adf0fbd1986bb039f1d4a411b273c4b15efa8cd935ad7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha9b158238fbd3fc4a8f0ef176e716fa108d528232c83ac1cae8149ae20576bad79a25a9ae4c945459c3b6063e74563216101c5524d12c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11118a768bada880de0767d68b3572c9b5986495e695b721f2778b5b59720ba5a486c84484065eecaaedac369aef4b799e9b94104a15486;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12ff54c0739671e95c8b03811cde4bcff6b3f4c693b53aa077021c8395152afd7da6be4853cb7b036f1404b95383930d58b4e0452c01511;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h164227bb945b1cb4156a2746720f3be0af8d19a2c894249a025273d5ce2ae2692413c45ac9b01feee27a7ea4770cd5b4bfbdab303e6bbb3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h33575e8d5e52702ca91b90b1825979dd8be8c7debfa140b717045888899bb7f3001c91ea452c1932ec7038be33f7da39b3919adb7b5a07;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h984afa3585e9720cc219d6a5b2683da1432c43c254a1fb5bb4bbac33a998470f81366779184f6175437a2caa36b1840cd17df8725fe799;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11085c277135a9115905e3e822726ef19707d0fd959120cb78203613da8775aed807e7bfd78617a4c3e5c6f9a07970bc53ea5affd899a4e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h15b4a6f49011f63b57bdcbdf29e490782c502c1158066b452399717b41576d5c295ee4a54d983a8d7066ef21c8800af507706dd8b9440ab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb218d03aff8c8bba9c368ff467054b513af8b5bb516bb9efb7ce60012928096553039c0863f9266584be3153ae809b647106f8b98d3af;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9a6e047b2201b528abbdb8e8e60408944464ba5c806550ae5b00801c9b7f06a6311eff5c5a5d382b6ba456875bf1812fe90b9e38ab42fe;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d9aab668da7ec53e770acbc328322aabf03a330c8aa336f2d195cfc6b2be6867fc4a1dc5fa4ee2e6cb720636ec60240b2c7cab8a4fb4eb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1633c6b69bf79661979044e9cbcd739797b18d53f9d3e06e5a4fdcd093c3f066eb112603fabcb6fde65f69032cf292b08ebe6b73f941ade;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1db31ccf104d3e232b2966d3a9708cd73c93e99235930b86cc3374a4d9b5865243995723e7e06f6d055d73413c227620e04a3179ba7e2d2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b4c8a8509114578021fd7b506a3427aed6ec172de738ae8e450ffbfee3fbbd4a87f0fd1cf8c73d62a4d2b3e7326fc83ed53c56f1d509e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c4e0c7f9d8721a15ce2f380323812764237aba79798c3308327704110c4c89165fc4d7200a1595f211ca349a3ef48f834257958ec8a027;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14c6288e1bcb62e4af94451fc6882f2b164a2e7ee8bc307c09b09fbd628fe12b2eff5b7fb39c82ba24c3da51ebe31ef6f46d63496d53456;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h499b9be1db3ff28ca4c0673263961dc0ecb4372c27425dff2833958b3a879515dc236656d44129a235d4b6af746c4ed3bc7622d5b64c3f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1221c847289391651b4bffed5b9f497dd547ae6863f72a4187f19f768ee7482ee8a047c21b73c17aba29297e1bde93dfad2319783e014a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc6e6a5eb5b75238015429e0f9545572d21574ec0898710c28937baca034fba288ed6c7af0497c336efc908096ffd74cbf3219eb1b7325f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf635f2e96fcddf6b30031f6640cca5646a21a03437cf6caf9b8e91d2fd604c525d11f45bec912bf6a4af14ffa2dedcb403e13af91d6ca2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1761be4ee1ab5b4e4fc78bd50c0bda65e4d697fa69abcc61aeb3081b39111edc4e9770bbc08ddcc04aaaf797338b9baaccebe748e896461;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6863e38ccd22784221602c1af27dd3e55ac486748caaec800ba7e20142df64b27c7fc1f083102752eeece56243e5e4a42440f82c50d1c9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha5f4d9ba9e0a3c243a4c8aa250986cd0927400dc1565d5ca4db9240eb8dfa543beb5f841c61d8dacb1b50072eff60d7eeb06e0b34200fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hec25e250e3713445fad2d792822d5e08c0cc6824687393fdab4c1a9c03ddfc6401b77c36446f676a658f2e3b4e4e294317e7c60f07ac95;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h92fb87f10ffa1cf46d3466ed684b499f64b74d1f4c4c97af191fc18282a1970a7dfc2735eab10317f1624e3ce2464e22b4aae67f64831d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9b91e708cb5f20cbab494507ae7689cafc4d30236af78ba99bf80fa429cc75406b60bfafed70bdbce8d12017b3eb04a7b2d12eff870dee;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4c23b7cca7b9190ce99949611b2451be04e8d30dbb93b0c644eb70997bce5c76c329e11f251b6d7b6ced26377fbbcabc68308b78ecda35;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12e85adcd5a6f4c9bbdafb0bc8e1a3aabf5ee3f0f0cf1986091388268ec3fbd85c1770247b2f4d24b9788b20e1328dcd953e55734e6b5bd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18b487ad274ddfc505c2124d1b9e2e608024427c4c7dc6f780ab07236638592fe4539157e4d74002f633d3c35f32be1592c2b4c76e0f349;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11e3775ec64f336b852fd20faa9d40aff1eb07282c12e4e55ec6c19746aee0f4f865796e5309e0e9a24f45651a7cf9f70b9600c7e6179ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h81af287d6e4ad2402db824634c7684fa0b798056aeb2ba85262faf2cfc433722990ff3bcd0d50ee8a208cc41a82b82eb066428014f6d3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h708a2089cefa251d7c337f191e2b4c63bf135c8cdd3d26b43614a5486face671ff58580f1fa0dc73988e8a2620c9d9e7a171aef65d7e2f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb81ea32e04b9b36cad144d731a6c8875ef3d94be00feae95c530f790e9e08674cc80dc410396a45dfba4f00dce0dd568a238b8bec5102;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d1789c67f7ee5a708e508c3551df33d32b030946f3b670b04b4ee94072a6d56c599706674cbd57facd2549b56b48f488a5cd28ebe578;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he4c22905cabda1cba2fad11194fe478b5cd9661de7f01b016cd2c8bc6c53fa8d9e378c04ce4dcf9c26c465656955ea50fc2c0391a4787d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7715e63f9a0fe615c241a1487ec953323d686eee62ba933619215adbf56dadcd4d596f24f8551f0ae6df2bb0c32446aa08f78ea5481afc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b0ca7bac74853a1d6b4e204f82e50d5898b46f72c37b95d199c49e0a2ab9f05f91330bcbbed8df9e2cc34edc633ef562cf3703358fc757;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d798d5ebd011dc60b86ff1abf901f92976fd679dbf907952f1e43e1531fa594d2c3a371cd9e7b85511c44895ee19ded58545602e9a8ee9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdb2e24ebbdea2a8dd1f669a7805ac46ea11be2c787311c2fcd0a6a939f95641075753dd98002b9c1466698aef26b98f85e8032ea3da42e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1bbf28c5728d0692cac7145fe4385f4c72ec3b6051277edacce2f535fd11bf125c2d282d42709edb398d8f9b53b9cdc897424021d449d41;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1040cfe0c2ab002da6061ff62b8b79390d108fb6698aa14a1591fc756d26049e0ca620f5adfb8004790298c7aec68b501d698a319111693;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf94542056abca1e8e1b732df030932f200a7227189502202039ae69813d72969689125652e6beeeff91bbf5dde261dc2b0e7954c4954c6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17efc67880410e60fc6084bc298a9e858db272085025c7e2ba127d65ea9a4b62b2f45ea943a8e859e975e468bfc3b1090c9c82f28db2c42;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h42a42bfe3f9bd3c617e195a20507207d84dd20342c9d48808860397da413732a6825eea02152ede3faaf68fcd7ca77a73a14f7e49646a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c05db4e96da93ae61272b1c6fbbab19c6a177b593773d0535c99d7c488a8d3cf130cc7ea3b6638566a8c1c2295e00c8dc9f9f7782139f8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hdce897ba982293505acc8e9181476dcef218be128d370d2c19b619361d38c251fdca48cfea65cd6fa8b9777e7949e480c06851d97f8fd8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1682eebc2fdc21b360c4b52627128ab0f1e34e7f03eb23861dd5c426f56f90047e7083c63e6a15663ea7ae39cf1d675a6f9ce594d3331f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b323a8cfeb55289c9326fb6b85520eb1cfb176c8700fddbb9aed773fd36612d182f4352f0e58c8f642e141bfa5a70e0244aba421b0c5a2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16c432bf54e1fb8698937d6aa81ce76764f84b46494d8275105e40ba5f58cd724a15f556fd88aa2cf514ecfbb74beedd175a6a353a8baa5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h603a4eb7cc335028a9001559823da6fa9329502a1a2fda93f55fb7733e8682aaef240e45a8bc2d0fa957ab9169f1032a6d934cb75c2138;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2827224845cb815ab0129398f2ea6447276305c4dea395999db1ad9d13c754684c1d69fc8767ba8a2d4e999cfc177b2838535850427ff8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h111c49b402b70d273904cfc6d12107c3d5c1f6c985be21ed2f6cdba568e353aac0b7d3da30d7d043c694a4e5f933f84887e877cc8b97415;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12efe07636d68274fb4565c66efed3b69590687732da0e6ab1cd4cd93912a68d8acda778386cee1736d89af5dad067f3ee62e735cbc529b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c814ea5e593bc50ee090119447b59290a387ffb3311071930601b3d7b0dd84cd8a0311665d991bac0339d17b01a798f055de77cc1a546;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h69b494336e0ba12b42e0c6c7c5b1b667b7a0263c8aebeba60f0015a892102a605609181b28627bcc51f6a1106d616a4789d29d44a640a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h75f1d8bc83f7e6f7f320d044f9be08d671343bd0944979c583d5772af5e35a5d8ca0c88d7ba2b73b0a92ae7b3a42c576191049f71d9cd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f6574c93c3ab6f1d988b2bacc60ad0d774b62660f414bbcf5a345789c564abf655274eb39289eae58c2ae50be489db3a7de2de81649cd1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'had945e9bfe07c64b7500c61e2f28c1e05304057f01b372960dc4809501ed18562ffa12ec8403e67a82e5131bcb5d5fa46f3a0afdc98e55;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d0e2cdcff68bb264806508e9be0add08950efb6331933b4f22b0575774e3a68c24f65080a75a9ffad00efd033e76fbf38f3e4da2baa674;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd1f34528b6e9086717c1efdfc4e0b0f027e611651f63729bb0a803fcca1e5864d619f5361db3a2965cc4835a7528c4104d23c11382c462;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h7a965942529c58097617920f47535096da123d275e12e1252ebaa274b04249e945b9ab6c15465baee90fb7682bf49f832d42c955317163;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb52fb9b6b73a4946df305099bcae55560ceb5e54d30528cbeefcaac6d734dbd440fb589ff5df78b1940f6af5f0aa9b02317be8b05a0f7d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hddb2850567f6f29a69a1cf038437f611f7e22d7dda28645d2439ba590d478383636d14c274b0d8f83bbf6b3f023d1125e65e7f5397dfb3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h270855ce6990b46cfeec1c550376a9c678334f1da8ab9a65e5d0aff73fad6da1a30d74b29d2bb3b7f65d3b1e8d8cba65ba659d70d64f45;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b00df5dda37606241b4d86c4c28dba38242781fb08eebcb7528f4ad9489de00c068745d218e229441ad5c9a27eb93f66b6dc28977e6f1e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13d416280f9ea048c335bc49d6bc22e35e4b09ee1e4f464917ea98305e3d7a725457d587395984e5ecd3a90a73711e286bf63ff79000da1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5c2c823a0a74a490bd157d4248689fd999652d3810d38c9f9f414aa1af8b94183b7f8b7f7cbd8cd1f1dd6e911cf1660eeb584c547bb2ac;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18059dabceaf4f2073128bfb89ac8b7432c1b7c636ebb96d38e3a77b59c4848cf2f57942397beecafb9d23986089000c07c4b5d52fa07f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h390b8212c625ebd97dce88e732d72e2f0273336f23399d81527e7f6cb3786aa4062a4023a8c860fbb5922bace545034f8740756d69151d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h94a02a4cae31b1d66063697700d1ff4880488ace18fede14b381067bf11c2c34e1cae532801961968b589db1803c6d29ab10ae56c1be24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16496409caf1cd9a1e20a7d615523ea345dd433ded90500f940220b96b0a797ca5d20b14133cf085b13eec869f83685bae2ab7112714170;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f6e451fea2c75fe1b7d977a1343bfd2e9c78bdd6e856232c727750076882b0047fd0fd197e2b539f8c07489b63d9feff87a291e98a326d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha31783f618858cc08c6a594ee38ef2311c537d4c432787ca14a654c741c663fa385f1da817341f6a91a6be3e8968aacd53b07b520c0b05;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h153fd760cd1a0c8fe229232148dc07dfca048f159d23e52f60c7391c01a0354fffaa9cfb0bd4175ce4c1d310257fd52ceae1cd67f9e2082;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h102951caee3c09023bc6a13e3bc3406482b586ab05b981259a7b46ad0fffb0a1a1aac857769194952fc67c0d6e0110ee26837ca8fd63b5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h102614cf61a3606c2025ed4eb7af5f1883039595ace02df80713e24650e2614fc11560e6e6375c455989a529fea68f26105fe2b3b205a62;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h68337903846be974182e8a8c73f72ea5c7154d7d750502d6735774ae0cb306b4877d7e080d376dbe845253f4d2ec6e365430f93e50dd90;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha84bc78d090ec7e1924e747a49b5b608ac1cbb1f74d736de7f05538bc991fd5c18a4ca8ee423c33956671db37c902dd2565550fb6e359e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d2d7a2eacdc78a42c620aa1531d41008a3873d861720a08171f7cbf3ee683dbdac768c099c99f1886481dc63b7fb9e64e15dcef7bf4b7c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfaf7b0ff2858fc5df21e75b53aa8ed17e885760c3fe23794833dafaf9b370d8f4bc411dd267a0d298ec759ba3ba51ebc447d1683742585;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9cf74d31bd98f042ffb4f3606ca4aedb43f779ad913769619c7590c0645f3c4dea08ae78bd30cd00460dfb7a89a81f136cbfe4e00f1918;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he582513c741ec65ec7aa97edfffa19ae12d8343f673cf89c30eddbc122a44d980be9d236c8849ba8377867c1982149fb6e54dd7f8c22ef;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13cd16ecf267b959692cf7a32c5d81f04039d40b7587a3ccaa6d9905f01f9c40ccfee1471c87476d1a41d8a5c10cc27298e44caa22cef10;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbd3b4607d54aed2894ed789877e1fb022a5f757e137e20e5f8656576ef8cc9e75d6c1df34f18c6be3437b6d035bcdfe552aaadeca277a6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he6010e964e2750ad3c768b25430e5fab3b6330513cd8b0b8feb6bf1c43e4926cf1f8e575f7694dc5d04e50088a658b82f713f227debc5a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h58461f68e0f2d9437a46c131855d079ec64417d16742d3f599bdbec9d1b867470d82a1f5f55e4cdbfb081e425041b3193e787f0a0c71d9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h108c34c9b38f0ae828f287145329006e774a28f29dff1065f916e433b3b9d67a92f9646102b0e5a16217ce335845e231b9a7f64009dd41c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1195db9fba45bf4a002706274d93c4acdb63006f4d5ac3005764aa2f10acdf074275cd4995188675efc06dd6d6e2f01ad7910f0743b4391;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1075e1c03e95b178613f71c8c3765e21a2cdc791721ab34781d61557766a5d0fbf8dc59c4ed6c5435bff4050ce1d2547b452661ff93e8bb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h62cc68ea2b61b69792765d63c2ee234d9175a908cd42689a8255d9e2d49f7971f2acf9c0e349244e4727175d8ccae7f8f73ca5594854b9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a24e7219cd3da5bac9654ad9cf7c5f26de3365c343fa82c48ec4fb2ee3c99ea7fe1f5bc5728867635f48b6e19ccca309b593c73b430fb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h668cb88523dfacd9db979b389cce0b2fa5028a4b1f7b11a4fbcd4019660078815184e3ea6f51f37d468e463b04239aaab90e6f6859d48e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h54f19778881ad096f53ffa45afddb5c6a0cba5a2f2e1f5aefaceaac79932818c5d6368479c6a67b873159aa25afd9d08206ab2efe2f36c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9f2fbbae3fc6d83937573e11777b3e876f79c45008ee58a28f3f39e56750afbb7cf665d1cf3bfeed635a6a15cd74036bfa11456fab5568;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h113dfdf481cf9fa76107ae9eaea77edd15e58971041fbe955672a2755d391d40081f4b4e06122bfd7a2fe5176339a368d452c554acb8e38;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aed6b44f8cb2c97647c70e5105c4e87f2c4f849e810e3ca721ce70ad210ad13dfbd8737ef6befeef77ecbe65a44d4b063ed2ba3b8a2812;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbe2b7075e1220a47def296ca9330492d6dcb0c2f24de6700dabf094bf898e02462556c48fa9b20e761c114b510ed11660fc443acf40d11;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h71bcaea2e9d304268705738f69835b9e09f80f5d021e522682835332e473ed55ff3a8395260267ae452b29ebcd3ae5410eecfe285f6365;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fcd8c0354cf6d6167b0ec9a3a173df31d066e7095afd9933a4c6027678a97f28567d940931fad98dee3cbdd1d7bb48f3510a4eeb03e00d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f0bcc03b48f071290a43b0585d62d08b3eaa24991f9d6ad87b5963cedf7c05d9cc95ba61589a41e1b41d7cf591066666129c3ee0602727;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h142ba44a89a919e85b12f79486ac61bbd9ff0bc35ee0789526b2fb0fa9f1e6dadfcb4509690a0f967a00255656085c21971e5f1866a8fb9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6f99b69b08d6de3a6098b3ed88bbb5ab8c07e5643b0ef363145171b7ccaeffe45b4749bc2ccaf4925f0860679c0cf8921cecfc172d3393;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8ad66f70ce3a14f616b6f27a87064d85a2a139a490f6eabbdf0c51335bca5ba2585c214b0a288f8af83a85bac3e26bab4bc29bf2543ae3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16985e95ab26aa67e1ee632e39c0fa48d99e109203bce1682e8c1bb4087992e144adca783fdcd8d873d5e1a921e5d3f9432328de5cd12d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h16ea99ac018a4cbfbe17e81fb21da426a13b3f2768965138644d3ad4e159a1caa43214e0316ddb89906b012ef531c39c62599423a721b92;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1450378ce2b29fc86a2bd363c57b36c1b8dc9969bf4b91bcec80df857f2761c352363f96fa9fed758f956800925cba7dabf145f60a744c1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14c94d693237b560ebbf546c6b839c5d8e1eb9df3ee3a6a389edfb94a208055b109eaaa7134363a7a6e4b928044d682ec126e773009be5c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17b001ea515976f88fd2b9b32a3f306f03845d878edc14239a69d98f02a1ab656899b2ec067393dbd2757f7c8530bdccd9166d457e897e4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1416737d10c41bc8bd1d3aad5769283adbf3606a0007da9097f47d44e7ed4feb4cf5d3fe1ed54b906501fe216b5017d96a6c9287a3c7fdd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h72318df6598611b85a9079807797ec0ded13ed4cbadec71ff809644c343c403b7c3dc639d769c754c4143764c8ac5e0ed88e6a0ace9558;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4ef399d754428fa363fc807b169f8e8ab211057fd3284cceff180f8abefbaba903662ffc474d0cbe6fbedc89f2ba7114437dd7b567303d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h28af2ca6701d15b9650b280b19d9f0fed8bc6aa23d3b8c1dff4e01e4ddfb758fec8fac17971d54a944d57bc33a26cbeea26fbcc31b3c27;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b7a2b0db5ffd6e5236af75ad58596e2f087979a452b8a45f4aa72b7731d50ea44838bb1a9a73618846650cfdf3a0060d9c8b7986daadce;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1246e49dc0a91de056b5fe33efd7dc42a2ae26a51dcc0bfa5170c7e77d071ba4b405e204df114ed1a3f27df81e4d22ea837423f18fb3ff9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b76c6a77a1af8632dbd21b9208416dcb1fe25d4997e034369a19d198d886329d9fdb37fbdab8e337ba66908b822ef7d84095f189d4343d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e1b50d3af2b4d90fd6011365aa682a6f9c137f40dadf2a7ae2f9566fa5034b76f9eb41586987692b8835e2102ad718632241b5cb744e79;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc1e856d0e1ac046567cd0351c723c54634c27a9bf8aeeda99a1a57804bd8ffc1c451e555c1191d04d3733f3c86ab726ec4a301590c5bf7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fc69f55d8db66c38d2cb3f64f6ee16102ac72c1cbc48ae5559f4945391e6f4c2f493c12e49af2c7524159c7fa05a49a13d47916db911a7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hec0e70ad4d423ff28414866b3aa8aed5a9b5ba75d4307003dd0ad1aa108076c77496f10f010718bb1bc21c4b1adce94774a78c474f9da6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1449f47a28ac828e899b26e8596b8e5f996449e144ec651e60a0dc35cd8fd79a94f1c576d2b7b0755a2ce347540b53cfb5ab9185f65627f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b089429ec6b404101989f4e04e6a6cada4ce263c5d53e28175c07366a45b8b8e5a6484fc44f63f6f359949494a1a206820679fc826cf05;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc1ef4d3ca2a3ea494e30d55372a359acc7ba0934f48412c9af0b21282635cfff63c8e694233efd7fccb38c8308d8ae15016bcc5ee9ad16;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'habe7dc2d2b5eb829703627e923de61f454fb4c55ddaa9c61ffdb3f60ea4e6096a70caff1ee15052a4dce38843499b6681b3ec46af030f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c2f8d1274b3d5522af0f7633716ead667b83887d50463db8b5dc9505bc49e29ac4f3af51778c36059672f19e6618386b64c7b54fe01291;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h166fcec00870684bc1fc8e0e35d95fd084cb071c4ab44e5c3006d1cce5f742c446f87fb74ac2f997c76548c4b549e1d40806e7a7fe50ba7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d40accbd68bc7e6509c6b3762c0a63fa4a21bccaaea78ffb532a62e323ae962c0bb04c97f691b92bcf84991fb8205573cd2bb9d80dd416;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11873a663d1ae4df25edd732fead9434451464baf4397eecf025eeb3c109652d4bd5dc7d842726f8d84510585ce88043829e40776082b14;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hef806ae3fb85a4dd9ce6fa6933ced98021d688f3bf50c415ce89c01c52fbef5c01f41ccf2471b4ad5e28f80518129d8bad8a41563f2b14;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcdb2471bfc051865985f56f0aa13911291e9739efc4e49943f9273f37f7ce7a07b7285a1ff9ea294d8bf998a17ee88c03c5ca940a676aa;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'he02a52ec393eef0ff6c6da5e735c47a969dad8831e587ab34f630a644bb9a7cc0190a21f25691b92c8772aaf7a7b8ddd7b8951d86dfce4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h81543ed86594b8f6b68abb5c1a3ace53cafe037bcf8b3755adb420953924eafa2e8693efa068e6fc2e26aea3c0fb326ffb0f9e0884adeb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f109d4636b1329876bb6292d20958988236145931b379d41a83ed361b7936dd0690774320318d5831dbd18065fa6fff2eb10637d1eb653;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h233600a2cd3460e9770d09c1b6054ee3d0c4417168b6a8a0d874c893c955caf8dd75a52d375eeecd9c9a58cb70f905e529831f017653fc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc2eaba69637d4fb398cb1987d441873812b928fc61e27b4a6330330fe690b9976e1c8d977f9cad7bd75e338b0c33cad062d45da06a54d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b1f90f3c9eb8c5f5636592663c8fafac5d02289457755f5488642e0fcf9588d7f6a32c30e418bd2f7e3361a344f2329cde94ec3fe55d8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fa894ccea08fb6af632cd3bae7bf51f134aa02dc42c78d0c618d2db0dfc804bb65ca30b253cf7cbfdbd6b174104d2fc3271aa1144b8fb0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19e3ad2f79e1e574507ac0d0296dcf0b5b9a12e02a00f06ed6ef862077753ca2395e2b90f0a25d9d7383085fa5dfdddcb4b4d027a9f4b71;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1656cfa9b8b8cb768f79831a46b7bc1f3bd8c05d699e3366cd2eaa4e4cfabf2574de0b669fa7f66e0d34b63b163917ec7d84da555b97ea2;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h448d485a18ff5bf81c27ec0aee1b338281c10a17f5b9bdff93fa0102b2eefd3e6579222b4654caec49d6879ff58587fc5c40d97f52e331;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12037bfedfc3483a58ed5b5f3974ec7402e9ec60bf2415b2cb883eff172d56c0f39d04ca77b80bb8d9b25c2212337534fdfed2f8e9b0a5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hb39b59271f6c24c8807ebbbc2eee0a74744e5e3284bfb0930738e553e9c4c1d8d1d332b5bd9fe9ff0076348ea0a82ae96328d380d91088;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h52632f8a2a9c874a256da1e1cf74f9984c5215e6cc54460c3c9471d5336ffa2b42d3c1c98d933312deadd02ee504bcb5649c27fff587f1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1fad65bfa93bda320092dad8bfb4104de1d6744217a04ec30abeffb8858c12fe7fae3c778f19e67188f12945d1a85550cfc3f63ca161045;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hfbbda7ac848a989d0e1e375350cccd6c976c05dc0f632c9a5b4d938d00a5fe3e07dfe8d7e485142cd0eb11bf47f0a6b08ed36736f5abfc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h13d980f9ec52785a74c39827eb5fca689f08c59e1a2067214ecc8a214889608e8572c84aa4e33b28526d222f78a08adb4b1a7b81d67aaa6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h9e42dcd355bbe4ba23f696cc9d1f29daa7eebbeb0cfca5bc4bf6cfe038e2957110a3370b7e777ee94fe1ca6ce36819fed0cf9b9c4cc40a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dedc7231e4c6c2a14c5cf4f708ddc231edff9bab5d647f5005646115622b3d18ee2e6c748f4f63cf56203ac42e8fd6de58fac12252f2ec;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f5616543a5027880e0b2e268d503c78c39b9932e9284a4efef31a0ecdee48df8fb1a998eda2f6049bf6ccb7c0d58208aaf9cfcc4d690db;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde93229cd643cf3c55c78b0e3b4ed8b5e8f15ae38c0bf0dffca70255dda5c01980b9456ed72e5557df24ad27334cbe78fc244f05d4a051;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd5a6259b8eb7b71e268c1eb9ee1e6018684d7b0409175b3b37c71fbd48552c39b7c3b28fe4a4c631cd61827f19891368ec495442cdc47f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1acc41e0f0a8d39cd394f9207710ebd238653fa9d0c9e41b2bb8f1bb435650a7dbafc56d60427692a1332ee4fec58d26af21840d7778101;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h153e55243156444c66d67d540deaf3165aa156059d820bebea874298b74955a95b35dbe5dc48d71cabff4ac9a87aeca6665bb8276581400;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cec114159b0feb5edcf4638c6f22f272268a0150644b254a1ed2256b4feb01622cf6afc07bb91b002f972f7a2f83ad75d97c59b9da0a38;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f33ad14d288ab98eda51420a4278b533ce6cfbae889a504c7a35891acb0c4126e2da96e630d8c36a42da3544c6f14eaee5135c9630750f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1351af03cf2a0ff64cd64b40db7a0beff9bb0686de17b58bb4bcb551478a9aef0bf1d9d66d0724e3e5e73174e9421f1124756d170d1a0d4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h183e4c5cdc370ae111e7aba5a03a11e933913e7c37c61dec7daed9abc97257b21357270e2a6935fd11ff322dbaf1c2b1c28599099bd6d2c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h43cb5692b340cab7a51d1fb622d61721e295e3a5349208e36c12abc70947542724559dcdea11d85a067f97ffbba8e3274b78141a02e88f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h10d585a4cff0ad45df8953573e8f697018c9606588584e1714030157044dc528f272564c004715f03b3b98ee3458a238621073420a94be5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11ef8315fc96f90518bd13bf07750dea138c429117e128008fb29a23b8b449e8358efe24f4a32ebbef57ca822a164cec244201dd431ca10;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h3579952b836f453136e32acbc358f89fed46a361859253ec9ea667bfe9761b1d71b65f4817e522d825a04e6c51fd5f50f043efdb8affa4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11a871e9cf8988a09023620071b74bd7248cc7e48bdf1e3f1e094eaf7c4d0708e28e6653ad32ddf985813c41ae737ccb66db5d2c7504e9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ad9df98f0a6971dace94cb02a462b7ce36b70d1016db78a828737804129165d70f20753e0e7647c421a558fd72907bc35b7076a8d12e36;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h2e237c9abb0dfb530c10e7ffddf94fe3bb0f8605d1722b74d27e348dddab73632ebab718d689ded892de69190878891cf5977b6ae2a995;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8d261f741469260a068358c2c8d5020025ea20790a2816582874ff505d880ad6016106bab752ea042f19c46eb41d19034794633a1d1642;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1491503e9441e6699d7a819a7c99855e6b2a99f4cd8e7e9b3b4d449ef5873effe968b2ad79a63db7aef3f260c8df6eb0ea64cdc41c193b0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c97207fa6b65bb797755d93042bf94ee70b8968a6aa59a5cddb576c7adfd9981aa329db53d010507a3bc3a4a2d22cb12566b5c9328619d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h193d1dcddf5d1d834e7fc19fdd73c76379b6a07d05cdb0b345041b418613fcc439d6108e1d0eca939f4f1e762ecf92ed73e71f4551b4b2d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcbd6c2d5e61afbd18858f202e20baace3074751ad95d5e48adcc7b0d3f4c3f25fd86a9a5b098653e3eb6c9f343846d320c5442fd68f01c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h101fd2f5947ba378e98b24ede62684d51fd81a8bd57f46b7180394b0265b809b550c34b864ab5fb8cf609f927d272af27f7be91e180b3a3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc823679564c8b169644a82029efa8b443e11affeb11f5a55d902a959181a4f07c41f2823d46438e9795da02c876f41b63100c28b9f00f3;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d6117866d213404c74847fdb86041db5b63df49be2b8fa33f06c79ef9a167d1fff5b4430950af8a34e7968100e350b9ecf1466975d8e24;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h993b1607b146f49a32f9e12166152014708f873f74c10b9da878a6056874239f6efef02cc8b595dcb8a05b2f859f6806c8e3aff4dca589;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1de7b11aebdc7cc1ed7fcc57eaf485e8aa73c7f17bf3a302cbe2f101780ac4b90afab5a4899e664dae5fe4f4f81bbe766736eeaf86bde72;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hcc9af46e99e765dddfac0e917443ff491339d48d3e586152dc563544f719792de360054daa5cfe64d897dff3d5990bb458e27e111295ad;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1f0f0c35a5fb80d4d0c7f2ff65ea6174703820b062cbae989c84663cae0e607edc00bc8d96e7d5433f44e26374ab964e53f5b27d9aef316;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h6de4ec5f94186d75ca25f9506253cb2b5881f5ef66cdd5a13e5dc3a77099c7471aad74d1e50112ad8f7528299aa01cf73eb8b88f43571d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1eb3f8245dfe9f0908390af22efe080a16dcd0f17e5e14414504d4f4edff371fa063a514c46e2d1fb440f3999c23fb23d0a49dcf86aebe0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1860947ab8087f39374e592b573fdb490bfeb8a87adba8c493a8519fcdeda8b741d82f55786f052bf73d436205783a152ebe58248fdf641;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d71b0a7be3c78cc28b537928ca0fc130dc2368a0cdf1ac90e4f172a907810b7183ac6fc596eb5c21d44167237a60e4460833361fa0e231;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h409126454211dde12b83b303040e75f396ac65fbdc8ccb97ed6b7b674d8a7a7005233bb4f0bf93b9855b9945b3581a927b0288abccb4a9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d6e4e298b83aaaeea1bcde5ead904fc06d4db3b8c3482a5d3de0e2ef594891e9a5d62317fe219ed611fb820da298a71cde3f4797c54b7d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h195a16b348cc08b17f861b326be725cb35a5ea79cad944b294a3e96e61cba1ec65e1a494e6d925929ffa82032d9f281125433b00b82bc1e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4a41ae33c3277a2159f42e103c4fb479a809308753bb0cf5c796149cb58810b16ff9ca04d509662d3761fe40bad443d795b6831481877f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14fe151b5cef5ff4df57beaf8cbe15040fd212660bd641651770e85dd2a8a4652e245501d468c55a238e9472d411570d4648753e97e9dda;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4b05260580d626a849834dba6cb8e83502069c8f0baf4232f1aab47a308854f77e74693a96c951c82f499aa517dcdcf26ccd0db8e515b6;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hba28b6513267238c798fff9ee75b3164d393e423fa33e0e4989c8d09dd4bb591977744bdbc338b547d82252fcf5ec87305c956af94247e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1af9a2bbb8cb9e14759808ec07f5dab7f608b4f133debc2c05795816421c984f6b64ce443c9a7422b1bb5243e4fe6bdabcdc45e6469153d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1578b131cd111bd4fb8d3c208f34a3be36f6c148974030df4ecb4d936704cd16a741b194f7a639e462d6ce1067b3e59c0ed37d02c7600bd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1ddacd3cc2db9d0751dc07ea4790023dfb6dcdcec4095a2b2fea7352dbeff4338e8c50d2046ef9bbfbafad168b5c2adfe704197b2edc83d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd2536ba5ca8020e95b0ee1a334ffe1565550e7050fd6e4cfad56eabcd918b13ea7a00b398f387b04c0fa31ad1f186734d2a0f6026ac567;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h12b7ce9e82bb576952ca162e9e31f21a505ea247bfe44f7d7b06d251d63e408665b35a7f34d551137699db520f493c82d45d7df3c4f160c;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c4b96cb4edbe7d4fcf0af43661f75850e07762819ad02c3a2218bfd7747c2fd2f1da12e0db1e983d328970947efb86a282ff63ac59cd84;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'ha63ef1c547a9e8cb9c723194df81ea981ac9f9e401774aadcb7ec93e7a7471b573cffb0af3800ea6b7bbfeadc306a889a5ab564fadeb5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1c25d2c5bb27fc31c0eb0f030f4a98b989e84a92de998745ee0084d09956bc4ea958492ca42eba24c81df68b9db7496599c02a64edaf4e8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1aba54575a492d2d7e4fdd2878e4a0861f262c0f77a5ef9cb83115ae7d4288433141898e6e852e934a5304765d8cb013150f2e54e2266e1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1488d47b5fd5c868d6b8189db380c0fe27ef921fb2cbfc6ed6fc1f0bc52d0cb3ce5f1be201f69f6781fcd5c2930675b2765bfedcb46ecf0;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf9ac312e135d418955c52ee158e16ae1a1c1406d99b96db7a21408315bd39fa4a3b3771446eb50e75456f523753456dd4010657b38eceb;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1cee305df08875220ba092288db4e1db83b6e987d3d4851d8d7eed5347483ac25eb8211dba60ddc69f419f4dd710e6bd1942bded2414757;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1e81d0895c4dddc0f26dffb5abaa406c4a36f0a3dc573147418e0272fd1ed38432bfc49070b44add30647fbaabf3b521c82f347eaacdad1;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8c8cd91e618a854193d0700ea5d4ca1fa5dec5e955ab63efa8a1d4abb8b146bcba5ce11c923b29ae6cb4b41a283b6ca3936106c110572b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5faa90c95dc3ff4fbba54e3e7137338d8790b4fb71c021b28cdb2745021c1a89360c7624d69385473a5bc3c4327fb8336f8cbdeb9177dd;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h4bff3952bca9e71c8e96c9d7b252770d68680c5c46c5de5395ce21bc7928339329e7720c7da16f5d9a43a275f3cccf77c161d483ad7398;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h18568298f12bf2ff4a8778e9b1d8e4a65ff2752c77948a822c031bed773ba3d6263a05c3e0d17d34a96d2b42322b1ad738c9f94de0a856b;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h952f45a27dc52e697c8f26d3675f6d8278390a3c743a49ca754a988b3380e108201b7aa4dc4b76d9db155eb2e16679a37ffda13df453cc;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hc6b5021d3691f0a6f14bfe1df982085e99c42b800928a9d0958540a43a62a48f21045dc1ed6cd1efbbebde69725f30942573348b1c0ef9;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1db2e6e7170220231cd238155d19cf525760025bd19a3f844a3476f281ee591a4cfa6cd44a5174d455c5cd70910cd3490be663a05e0de5;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h70fe824989a45f9c0ea71daf65401051cd9f6147cc78b28bfd22f4683b541282c04c5937e0e2e746135a05313384018e5ec4d166ea213e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hab08216266e061a9587dcb15f6465380b9955346b4aa0f61b824d9d315aa32146f5f7aca7401d5c597111e71cf975a048e63b03fc70380;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h99eaf40a31cc3beadf6be5eaf1d9469769385f804ded5ff8217c147c737af8c6c16f77d294fc9e228c5072a74453548389f50ffdd55d0d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1976a3690aabe404f9d0cd12236a7d259bd5b51a9dfd92fefe0f0ea1ea4594572d55987bd22cc2fa52e28aeb05ec246a8a295a277d05eab;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd7ada8d596c8f53b4f9316737a776e3b6079479d15666bc032861bcb95b922bf5c9721cf52eb8ef8421b3a41f769bd79e5c3bafa57505f;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h169ef582dbaff647d9c1056b75376217f17d83037d637598d8994bfecca107f03f725b5f46722005b82ffbcab8922cbced11dcc78a0e3b4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hf3f96beb34e934686c4febbffe6235ba69d3912157b0f1a2d5187b45f319391b94581b2f747a89c7a0532eb78517d4900a177399f3bad8;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h19af374f13d9e57c76429c7a64e9de5668050364f1ba84cd41aba8623eda84d87ecf84e2f3263570ea5f6f256385e5b16834fecf9f94674;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h17535564a5df6fdb118bbfce6a7c217bfffc04e9e206216acefd4d1530adfcf1d6462911a1069dce3fd751ed407e04cc912d87fc0bc058d;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h82045d1b0ab75c4b7b8fb489b739ce9bef778382911ad18b8a45416498a61a4fc8a7b5714c163d6dc11c47832e60f2e54968683c09b574;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1b6fce675df3fe5d563152c27fa4f8e4230fd1c05cc805f7b9ea01d6bc3835462ef40e5084dc808a49c7a9cc7b5f59f9869527f01e31e77;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h5f5f14dbe8f3bba7663db0bfc49588dd66a23cb7bcfe0a65c76cc515157c6c0c1a081682a185df25308a9facd1505af1ff115abbfc26a4;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h8514ca4c35d622d1b73ccb96ce7ce3c4e546eb4beab256204b0b414a05232a81954a8bcade459b80d95a73f15bba958f187cfce820768;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hde1d66184be185061d67cd290657d24bab37a64d91b7856c86873135b294973e4d4d0adfc6d6115e37d3dc1e2b5d60367defab0731fdf;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hd0cffa1dd10ff4d7f390d7b6ff3e453bb395f5acbd6b972d72771f9106c5c6a1c7e039f2186d67597292a87366a1b187c1bfa1e8534e75;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h77323e098ef201a0cb0b3af03fb554bf2a2a7de782ebcdfd47f73eb2ef8850ff2f501e4590cda3eb3702fc5652f54958676990a5f53e13;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'hbfd6620139734f30deeaaa9fdda83c6fcb23a6117465b26de1fd30bf4e33ce37ac8c33e8dda6a955e61bb80f24360e32690ed36fc165ed;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h11cdc15a6c2b77ff7f3c4c75c76679bfb9c739a6ea24391ab3c36dd424187abca97e1dee4e23e64bda67e439b44b067cb65228c3d7f9834;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h264134051ff79de3df15e81fe1be20b730c15e8ca82f23b572e6520c47efb770c721419c487edf75f25f55e32006e7837ea063af766a82;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h138532a0e8f2b8197f9711885dd311fa02666ead389354284952ddfa43cf87f0209c4ca5be6482ab06154d89d9e8d67fa4a2d76a555bbc7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h14dcf922c3c0f3057d88a7067d4cc9aadf17d748bb8fd453ad378733755d079ec73ac67521bc0fa6c02ca6c8e71292f3f9372e59a29b2f7;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1d5cfc34626928fc8840d526aa39cbc969ad04bd84fb36111b8aa6d1325d6a5593208458b9b00114ecd0fb7da54f0c342e49da7b352ce9a;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1dc0815cb1f46a8f5976454f68699b6ec936ff3ffa373277f616f6ced6fea1562169d8fe63868f9134b84ad7589caaa678b472cd54dbe2e;
        #1
        {src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 441'h1820ec3f6a1d43e1416bae86ea5822ce000f4861e19a2f90d69be327eddc0c9729b1ce6f8c49abf4912ac3752b077a615f425f48380f910;
        #1
        $finish();
    end
endmodule
