module testbench();
    reg [30:0] src0;
    reg [30:0] src1;
    reg [30:0] src2;
    reg [30:0] src3;
    reg [30:0] src4;
    reg [30:0] src5;
    reg [30:0] src6;
    reg [30:0] src7;
    reg [30:0] src8;
    reg [30:0] src9;
    reg [30:0] src10;
    reg [30:0] src11;
    reg [30:0] src12;
    reg [30:0] src13;
    reg [30:0] src14;
    reg [30:0] src15;
    reg [30:0] src16;
    reg [30:0] src17;
    reg [30:0] src18;
    reg [30:0] src19;
    reg [30:0] src20;
    reg [30:0] src21;
    reg [30:0] src22;
    reg [30:0] src23;
    reg [30:0] src24;
    reg [30:0] src25;
    reg [30:0] src26;
    reg [30:0] src27;
    reg [30:0] src28;
    reg [30:0] src29;
    reg [30:0] src30;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [35:0] srcsum;
    wire [35:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30])<<30);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9045c8643b7ffe5a657a689f4bff09ab00b236e11c5ce61c619b33f906607b7f440357b42c7299e0c2b03b57dcd1e239407ee7bdf7974a72c24a2c1a9064bfffe99d35acc9c1e4b50394ba28a71f6815400caaf9a56bc52890f535c85b8b74d3fbd68834c3fc38050ac9907f21c5036f32f651d519cec7e0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h720174bcd4029541d28541ef12d352abc649c38f89ebf030584bcff4b721e02af34cd3e904c30c4548bb76b4c9634baedf83a3f050ecd17f73faf25c98fab3080ff4a5ef4604ca89c40ff0d63046a94c8122ea50b0ecd822690b6d26e08c48efcc5f545cdf04b16084b187676ab3469ac803c0cbbdd7210c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13384a316f2c463c568be2be9d91b40acb25b0622fc5c4a8f31d6129acda9cb2273855af8b59344263bad01da27c72e3dfb4c089971fd0bf598a6c2b39ba6f5c59cb468ce57cc04fa97331ba5a51c6105e03c8de38e2dfb6483e2bc70a4c5db8a028a1a4e5287994d8ee9985844e5edf3530a273ea0d90cf6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc67433a5729971f5bf1182a402b2eeff1965fc059098346456fa5ad68b2206ff354a3bf7aaa8cb650783804f520f7bcff7f36ca871eb4c440036fd760cee336ea67f844a2420863d2c79f10d041601bc398e0d959c5ebb1ea03232a6589178af52a039660863f690cf66ef5ac96d4383d19e475833a418b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14fa3ae0c87d82030cadccbb0d93fb205e3a0326aba9c241dfdb1db6ff4e6a1d4f779e8faad1fed28dcf7f8cbf86270ec6ee0c53f13023f41bceca19bf7eeee6530b9ad81f8c1bb5e091bea840c24c5c713582e68fe238da6f63b4d1eb302ebde77b1b03687392fd7492f8ac6857d0c545602461ee9b4f351;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he749d012a7c2a8d4a241d85dc7ff86a8b7f3b38f9ac3ea95a986ec029c013b432c33573863f8c76a1db40e62f84a2a37893f85779818c68f989ac80270dd176b717a1244d6720ab46a48e4a275c5188edf9ea36f33103545a54f95531e9032765730835beb35c53d260d782c03dc797d28247eea8ddf35ea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc5b542336ca0b9f637ef759cc55f0aeed4c2e3c5309228a896fbdc97a5da2e8f01acbc7705d6c9c9ae41e8de9c8184c17471a2f501e6a0b395326c5291d14b3c308a89e10121a551673c526e36d71c60bcba8677add259a0edeb4a1305f355309c5572c14f69d48b47f18d61cf26fc307153d1c5b100c563;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15568866ef50affb31390df02f175c9159c8d31b26d71ae1c84d0fd11524b75f2262ec57ef87f705944b1d7490cc9227925bf9f879943449e5ddc043d7ebfa89655fd2d503d787a3caeeb7ca9467081762688460d5345608380a2bbdcfeaff97623d6779e1367957cc327e48218c13ce2d7841ab2f6826d2f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16844bae5ae1d80f01d2ead80166f58282d3d80d55af11d88e5bc5bd74bcc1fbc768492221e88da35ac2da4d61a470bbaa07abcece4dfd8f74a23a003e698760aea7d476a16dc3676b10a7ff10607d32e6458a67eedb23840e950c13e259e7cad8e05a867e37d84871a20375a7d3ecb20afad10f605ede0cf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h424eaba43058ce0a130608335855883bcd72de19562051e2d51ed0407395a3941c0fbe99b9ff8ca6586f1acd918d3f5e69d4a97b148b9187e68df913cf775a726f1c0a00dcc1a90967541576062170a9ed489d0cc505168e14543747f9079bbaf3bb830116ddc78f7a7618b5bf0e6a6ce4d946651c9fe799;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4c65b1a4af1d164add819e75e13f225267d767a4b06e33e71778cb9a3740f6ae8de00c892c12e5b9ee54edcfee6cb70f953dc7b3917c82292408e1796ec7aa91926628c7bec6d513bce4d9a356922b1a454e59dc641c4943c8a59abc7c86689b69e5f4fddafd23f75c51a0793440ef410c9b5dc2ca3f9f39;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc0e602c5e0a7f4e1c9b87b2876a0c5329e896b17c1edaf6c39c24eaad4d53c21e81d78b42ca005bf0f6ceb3044ad6150547cee70b35bdc289eaf06883008eee7399f25bd1c5ff185468dec71638dfc6f741f1d0605e6232a0ed418b5d12f3e2515310cdb590942c40cf9e7100abfe4184bad510d7faa3c52;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8e5dc8b111bbbf2a2e4c0006b986f257a6c34a2a6d1271b4c2d8365eb2972eff81473ff5b7e0fcf602d20839cae8e260ac72ddc6aeb30e1d4dc4712c6a02e9f07c7d3e8b4b82a3315c79c4c1927e9638ecf288bcbbde17e4b4ad8fafc54881ce956a8e903565977c4133abdb8e744775f59399248f8001cf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c6940807fab831e6cd36cc112e7c53afe3344ce85f31853976b0926c10f79fa65562a67b17e0e579f90dea266a098d0ee4b4d11cd15bac41253afc68ef4a30a16be4b10f395a02542a60ba438ca2c8ebc5e4c6643ee7bb8ea236ae58e760141347ca07057ad2b2b9eb5233700ac24da94709995c838ec857;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c7f281af07258f90c6bdb846aff24f870a089e47a3af36403e6b84f762756afb7b9b7e9337d6efa99a902988339efa826cb7404acc5a910d59e09515e83470d358c41c6ad23d082064b6c3a17579ee00fe66012d4f1794376675aeed0220ee2ca866a428ee0e032fa8c92ec76ef57cfcf5153d6537d14985;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e84a0c0eabc817b9ad6dcf103ea676d7ae4cd30d094a9f77aa4c19e38ae27507d2101f38ceeaa6d29053478719fd49edf0a9d3f6eeddd342083637f4e5b320f0e69e2d178f63aae97da65f386d966b55ff8079daeb61eb266cc06c30f35e8d69f53a47fbf5d1a0b159c5f1f2a661436e26c99724fbf94cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11277b6f2d0b07dad58a6d41ffa11de61430538eb8d2df5e79cbce48d186e9ef17ee8a9b78a2c6a26e9d4d0337e0b6a475b1f95d4ceb8fb9a80ac7731ed6bfeb7722a999955ac719d018d624856db29bb3eb4ecdc0e4e53c543d3d980b90e1235acf6d3f1f8a0d79466e50de59a6fbc349d9d08392a7adc4f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h142c426cd4dc125b1fccb1f99173655cf0110574c5addcf8c3d685aeea8dc61d22e068046d443a82a440366fd003e6dbd7559d5556661d7e917138fdac6a3f8bc6888f311cec47b1c1651c59c9754e854e3c2b0f5b3047b9477236ca029bfb8daa76f73539a0abdd694e1d2121c9643c7a205a8a534bb0ed1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h58c0004e0a5af9275cd566defff2c3a4e00f81b1992e4b5d44001fca379fca5949519cd17fa302b6e1a4676e7dfd3b6619fd8f2e7d686f707fee45a1ebabe584f7c3e43e0a900b70df406508a78aa28f4d9454a2089634a3c17aa13b2295d4a92cc10ef383fba07f0ced84beb70c576fac44ff934d7934ed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfd6c468efeaebbc9a5389fc95cf586ca239094f861321f1a1e7504b73d98572d94eb0790475dcfc6a94780419835a0a456b64c430cc954aa8db94103d643c25c08ffea38ab48a3b851e32b062b97507120dd3e6288b6cd9ec28b6e9576f9e49b39f024c7757eb3690677a06ac24a6420b884758f1ee86b3c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h961f909cd76e3c773c0025c6cf8ec3cbc4134e6bfc09edd46c13a3acd494552fa11d798cddc020949a7e87ff8321c21fe7877b93c715f07725b1a769601d794ddabb4036aa341a741274df7bfeb58a2c9ee09d33bf0c23fe8c3fc66f34ed6a2dcecd94cd42243241ee3c3ef7e9fd8df6dddd420bb061fb24;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10023f086e25388239400e1f16fa81a3b9ab511117f3a73f478419b05106f13a000e234d8bdb189ed5f6dfcee82386a459af0eef1de076a5345ad800d9af179e03551754755384689b4583076293b3c81546a7314411447beb8cf7be25512e58816c982d6032084e5fbd8585b931c068fb6de9a38963d2419;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dde42bbbb4b07ec8e19968f0209564c9de36c04d88cce664cae126f16e8a97ceafd348676c620e618b28ca072851e1c9c1364bc2a1fa249168b53c3e5a88d1f23a1e2aaa1eab6ad8652aefe4653850c361241e1bcb87005cd9b748fa53d30c2cb6e70225865fe7255ee0bea1c36fc38a7870798421949fb7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd22f4c1c5ceffc85374062b9deae64a9eeae9f0ba38d039415e9b3c91aef17ff1c34a4827cd488d81e7a8a6ca02c9fb2f204c5579027167d233c065f8fc6efd9a69e35b1fe059f6e370821f090ebb0c56cf3b1e2adba5320513c30dfbfdb279977f0f291b463bc699640796e60c31fde7efcfa0a32a9f6aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h114e56e931648f9c4339f2e47e4b18bc41741c7c37f68f67915926044cade4df47156d462f4926b239f3b0c4cff5671111d99b4d9a4672b6448da23941329fba5ea5b5795314eb651b7face7af58c75a08808deed728272974f770b4f97894c645b082c3f7d3a9df2aef3bf1bd9aae15fb936a568ad66b8e7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15e89ff647e54ed72c063c6e716c34f2b5cb6b050ed98d9b41a15c325cf643acf95c578aa4e78e454c5d0fd8dbfaadf14c6e49579e7f08a4b6cbd8b877349ea59acaeae72045fcd94251ab07c2c818731362dbc7dbea276c23a6812c0f2eabf24b21ae3b74ade831edafb21a68fee1a08e8607035140d8e82;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f0fd60dd24900ba4b6e6059c416969398c1057820eeea588ea232f9c83c37037253edb573c6872f4b884dbf3eac4d42f8939ac24377596a1ca7fb7f8b4485378644a5d6e906b54c7697e2af691a352ef7e6e9ad39a41d4794e99c02a6980c14a008aafd452758bc2101bc64bc49bffe697d96681f6d9e59a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17ea5197c6732fb0f4bdff7951c50910c5829eefc3b7816618377af4748ed7c883be04c9434cf695a6ef6619fd9c862bf54977e6a8c6cb525684aa8352a8bef66d59700eb61a195167f0bb69f997272b180e9fb341ba96f9d5551f8a940b7a937f251779d2391d5be970bcba3fb2aa2ac1ec3ebe11e83c336;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d6b97621c9a61c3ecbe7c1d299902fb7edc421a6a0cbfef9e50bcae7bd4753bd832d395fdd7e1200aa3384cdfb3b05242b1021361deb6afbb406dd4009151472b4c38ae734382354130edaf04ab6f6ee02eef6d3e5c6c240e243bbeef1d63d4ef6f0dc56a4032b92591e7909cbb06956948baa8998364642;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdfa64b6864b479360432ec3e10f921775a23a8fb065ead6bab575da5f3176315c4d509fce63804dfeeb16d11ce81672884f2f7229b7bce042245596f4631089bdbc262dc8ae2e86c57fb5175b1b71831804c0568950312bf278f112dd7c9ed0bda8c71c7a97fbe479d938856a575a770d17bd6e0d923ee28;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h76ecf67d5ae6d1422886ee84252f4e1c10709f96d522e52bbf89de87adf84547d09b27729e476c9c35e328c96484e6dcbc9f8f48e65f997ad09ea03d49303d9f51717224afcc49ded1cb0412bde8f1076c9ccd96729635cbe3c855d4503a07f0941d62b5fb7c67b0ab4402db14b7f7a833b58ed7e727f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h182a262d44e5d42eb02114fcacc5f248303e925ce535ef4f414dad8b2ee27d320683bc20df03184cbe4917672d9311c3fa76356c063f37bd2d9d3648402a6db024e061f369b3d9416d80579dca811ce15abbab553b38bb5a21a181a7185b0ffa3b78d5447475a4e8c28608ccba6e17a2a116d3f78f81332a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h169b4ff6b3f1bff4d2dd703c95fc46800f8907d74e6f1a74543e99110d08ef486f3c895a2467603a47e1b127dd936e99c23afc470337a92fc80d7349155a01908c10bacb6968f605ad44d8fc40a65832f2feffbfd6222e622539585dd0d618c472bdb9f716eb00591ab7207c18452c341440da6ea48f2a532;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9136dd9af463e8448e89c78df671781f47458ab3adf6b8f3d71d49cab4030e6670e9d521f9a0fae103d5f9d2a2a670c7af634e69068c53aaa534201633a8e8261e9125d72fbd9fa66253083c1cb471f487226671b00df737c55a58bd5351ec129f742d2898c95d2755f5d93c85d0d3449199150e4e5756a4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h678cb595ed471f37abb876d5e7e7f842d52260e7e634cfc0d377a34c287135d9f4ca17532c07e8d788c51365bcfbe489c9f68d89cd155fff7b266dcf6a4cc1fa7a0cd1d6148e9744991930d34f80be438974f8c16c0952a6b72da96a66774c16af467c7c4b45eefa91c5949b51faf51c5faa3c980c8321f9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h141fca44b027ed3837ed48eadd501e9684ab1339519ed34d8e46e91218425540ed676c67dab7eee05f83312101b35d2404e6de4a8204c0efa8b83a3a996249a7bdfe910b828a25d377978f1bd7ed0741be55fe75b190ef7e1ca01975cab427d9171c718af835de1e94bbb55ce518f3eca221f71419c94fdab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c50e0a1e0f6e20b1ed5a9f5edb70e5c1c3f8b368ee2cbdbe95cff6013ef57b75f5c44906e39e139a37ed5ebc057440b8e6a37d6839c1730cc91049545892712c22bc3d093998386c09660a190d85d9aae1b2cf2602bb530aeffbc9e524e321220f21e717c84c405e4cd11ee08194a85fef7063a737987d21;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1285b47a44358739692b6d51aa039916c4aeb30b4ccf1f36850ad827127a3562c13664eafef5b2015e87a73a8950a0ff171f05e43a104804986617ed5cb7316bd8ec6b8a9ec98825400180c5bbc931efbb12479b62a01edfde2ca0ae2b324052b64e03111bca1704d012f00eb1a5add9abde5528b228db6d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd24a6a18a42f45918196a7e5fcadaa860bd2186558fde7757122f6a0470a136d0d241262107c2f37a7d1f4247612cebafee565f486d4bdbc33f8a5d0f91c039c5dd26496a8db08439081d1b28a26a16549ca0d0601951f1fb82610f791f7baa2e17c25aa9e62d874fc563c4a6104f7a44403c809abf6b1a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10bbc1660bfbb0f4567310be77100023069e6488e192b47b776e4c6e552b38e3c3e9de7a14df3b8cd969442dd2586b7c13647dfd14a77baa565eb989e4ff37032f8c773b10b8d76777e47f0711af39e742da8a7bd5dbc799038cf771d0d24fcec0fc6b4a746a2f6ef970a27b709c9af94753230bd8c7fcbcd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha7781c3eed14811435c4048e86072184da56a78a0e97f7633cb116388fe98209a15ee69d0861db2dbe25468e54da6787068b835de5fd27de0edd6a0ad4f50dc206f93dfa7290cb3afc35301a00e52317f236d5a493c6a3a54de11e4d23c4cc2acb695e623af7684d5ca104493772b5f8ddbb13ecf35379;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ef1bf22f032ad0c9e3836ef7a640ec0cc1cbf4983e7130c93166b6e65dfd84e9e1445301b0f0d22f8b980250e202e5c71b03cc56c8b592fa93bc63c7e692ff31f0790376eff55d59fc446f642e49c5d9769794a40934371ac0d9550e44a40b77959e0f5330a5ff37d8845ac97362e5eb7279ea1fc1631e15;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1674349e0ba4605000665fb9efcfa084059235f9fed7e0d95010f2fc7d89b02a808580d084b61a1c1447161c66470078e5c85f82038a7893caebfb3d476335a9f1d642a00afece981239c50c55a28926d8660eda7d1d772c5bdd34e6dd9d1b2dd4eee2647601ec222de5a08042814e0af4e462a04ea6b79a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15e5b88ff7af32b0eb5a23a36d395a2d07e0c1fac6bc8d40b7a7a38056383d56a74376d393bef7e334ba3774e87a90140a4a2fa208cbc447de52f176291b0a499baf5617052649257ea764f4499a6da3d4b2506d26fd7f41d98e3d3ceaa159e3a15e88600b2db8804eeeea81a12db6c4837b974bd125406e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9912091d16566eec0be59c3fa51bf1767929d49dbebd10a0115f04c493fcfe51211e2cd5d199a95903c3d7e05ffad933dabcc3c3877f2c64bbe6072cf2bb8c48dd3fdc5990dcfd24304078e8d0cde8c9caecc80cde118085be5a1080fb065bd9cf3819a5f1033bb1cc8f17dd52c4571cc1ee1090742a8814;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cd5b89e23790265c8b85ce8742f4e1656510efe56570dd872815841fa165cf3ea168ac48ef47f37a3f15e0b7b3d2f85b2fb5d4b976e7a207038c243da05333ff78a42043295e7bce3d0ef28dd1d07bf888a467a51cc9a9884a4c30a6334d349b5d8f3719bc624c9d4e4daedfe87e0a3deebf1c705b408c1c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb83bb4a71002ba117cd7531d65db84855626ddd522206894263a26686e14a03da4718aeca83f1f036f4f603340d7d6c850a01466c8a0d69e18917e2a568cf415c9dd8ab18174786f9db084867b04ee87d260ca579555c28a230a5b05d728245db30853e1e8c7be8520777210e18944d80f05a2838b07ca6d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf5ed8091a5bec10d4087b7ddefb5a75b6b48e1c8f1494d84f679031e26b39ea3754d5d695abbeb9f013250d39181586ef837772afbee8ed5abc2741293a199f7b8012f251e57cf19c8d12530c334bdfcf19cb84da964e63dad40b61066a306728ae01ca3965cbc2707dfb458eb75f504fc09da0238acdc5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h137426134f79de040dd249571ccf4c1f7f1e010313c06a1f60d90609afd270171b5faf4af1f3e016c6263e619395ebdfa7f33a29de94c436a1b778adda2f9003b0b58522535146fddfbac1f40d0ac8c1818dd38b616a7a61cb6b72343cf1c977c6873582bd3e32c3afe88574287c1edae0444a6adb05534b7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h168b7265abbd5bff2cb9a73c82e284695c456885323a51cfc11f183007096879a731a5e9b6602b2176cbc451137412d14c659eff9b8b3e5512bd24b0f98f35da80e458e8a10b2bddd1b8caa9d4b7dc4ab002482bea840331fdbdc7b27630cc0a5c05a6b8a9c25937a430eaad23ad16d6f9d2eb8ed3e9e0551;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h75e6fe7b66393ebec55775504c17659198976b66dc4eee9a8042ea2679c0b10332bcbfb0bd887cec3f7a5758fd8b4881298a4cc023b04cc9ea8b0efb705def619ad477733b71f83c8854a71c9a3fb39ea46716ffa30d35b827ee5f3a9623335baef088610f0becaa9454e2eb619af2940040dc4c3d89e71b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12aaa2aec6bd94cdff139ab0d27c0759f464fe6866a33cc6dfe873cca0be243f4b1239da79ce15fa4e0ec577e240f5e7b092c07af47f10389e98bf053cc22a3209e48b352f47bc4e7c00ca8c627a40c9736eaf02bacb2388eafb74ba91e05bceb34e3765480f642d2e05b7dff9a34dd21ed336c878577b1c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2642ed9062308196ab358533b8825d856d1cd766f0a54cddfb6ca90d8bebe95a1a133342914209b13af1897b0b16837d491b38be43897749017d311f54c33a983844aec1bfac4a5c09babb634e58c7a388a8f23dd08533c33c96fe7aa3e58f479f4094267c4a7e41e8213f60756e9e656f9f309e45cfb328;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h64be9cb1212615cfc8713f794b7fdc58829a6f06e4340cf0f1b8c8acb022546066af96351cab2b0a1ec5e2e6508429ef6952e07c15fe0dace4cd611bbf51bd149f7cecee9a22035613a3e98a07119d1bd6e2325a2a64488c7643b2599e2c25ff9f7439ca53e534aaf770b1ad17dc35d31e2fc9eea79b26de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc60cfb2214ba5904052b5ccb9a1e49b00c645e94b2df63dd0ce7804e232d8b9ac28fd0c3f0e4f6bec777317d6f9d1b84fe87efaf644e23c9db0d197c55990f91ab845fb138db515191b6984b852d68e29b729e9c7fd6b8baf3331f26085df20e688a6791baac383bab42bdb3fce0da815e183bd4eaab125a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h268fc800fd5caa3322a0840e7b5225b7b8ec4a2a9e0c022e02a0a011133428286718ad21c8c0f219dabc29932ec1ae0c15c1166701aeec3304abb0e7719cbe65892d5cb1452b5f30f03ec8ee97552f72cd1956096ab6ff79e6f896a0cb7ee5e8088e7dedc21fa41162ce08270d1f49ca4087f9540c742d70;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h55b6221ee531dada6d19e0c333f645d382962204898cbdb6c5e639fe3336c4cd97bee465f254868b859263cf10d0fc9c683e2c5da65da037152cc78b1cb634ac46222934a95fdbebc6de01012db14bc9ca5ecfe1223b8dae4ce88213c012b72c3f8569701bfad39ae3bd5977fb1e0675c8f45881df946f3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5b779776b412ec417d2bd4ebdba2d40739a3e565c7b7b1fa65327b53221ea12261d78be4349e086698bf6581e94087cf918c4f24f5c2451647ccd7005ae1478915c0b86df8ca87499f26802aaa8bcbafa7bb54c9e8652a5db4fcc2a654cf87ea8c51518eb4f33203d6e6d8682df29479cb85ea77b6efdbe5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e9748946e1ad49d5e927cdffe38e877ca388631edd64c03054e211fd3efafbcf8a75aec536c5a8899af01e5fc721c82759869675a3e817ef0c2c9d04b68d8f27506f02501b811af806f0079068cf541b525e7631ca2bae0eab4cdacfceac33514d34fbf8b1774f4a09b6cc873e585232e6f1658fa724f30f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfcf794bb0c62fc2b5e7e85a9be99f9d0cd05001c4f14e74eeb19827bbabd9c5de024575700f816b4afb2d00aa999977602855df750291055a96fc738de5d1a110aa5b979b51ebfb3bc16e9ea14f100428a458f63bacf0de92e8da83b070a5e557e691a5db0109aeb9fbb3c6c1a2b9fba2d8a503154f3c287;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc3358a50901296af7f7bc864ce491c850e76d8168d3372b73575c7a4cc541539b99b792771933da068f334433dda42f164c087fedd124c9ecd4fdf4dec736d4e94efbe8a114b17f23417052ac4bfb5558997263161ee1e5df94cc75dfb5da9ef970241e7a5678b71e3a32e6bdffa270b09eb0d581ddd7be6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h79b8fecec2816fe975c12f5af562bc6770d94ca5d155c51f4b0c79fbf07ccca1b1de487003494bb6d5ba7b95c4d8cf61ecad389362842e57789f6c2dac6806f7aa14c7f46409a2cfa56e1a89e7b735af17d2b90f6f6cf5a3d5cb1b42cf627afee2fd24d2f8785a28182c8eee77bdd009c84a6a85d3975701;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e8c6959762817759f88b82af6f98ca86270e2ff0e18fbc527f0d805e7a34d2553616184982a8190ece123e4938506f916e25a45eca67e14c44370b8cbca7c5d1e8551048627cca5c5bcb3e88339e3cca9031aea6f6bc6fd4075b36171c701df2876a3d79030160c549099804ce51b3c3986eaa7b76cfb8c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15db930b97f8ef5e9e6fb9a6b88eaf0354357b66e7be656aa38bba7839d555b1f61b6c869649f91996197fbdc645d085fe43207528f58723e6af6be107b8dc8b8bf48559bfc4605f34b2d20793dd739b7539d7a9d6f04121180661a3bd62c1bcbcfdcfd400ed580f6c08cf21c4fcb1b3d7998b0c226da57fb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h53612d25f055c0dd8e6a2b696755143015b7bad4119e3b3ac3dad96fa24e9341300477f4811a3dbedbc23994eac4aef85ceaa3213e81d6af6444586850161ee6209afa7b2c8c0590255e1c9ead4fe4ad8f556f1547e79ea736fbc6737f93b5e2eb986e9d55bb235312c8f104e769e7366b4881c2bab22384;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13052a5612dbad809b464a39d19565504fa2526daddf29f6cea633a3d4be40a7617393e58f2bb95b8fb61e5f567cc31bbc39e5d67cdecdc8a1d88a52e82d1991708510b23f84a64225f3cea6555529499cf836c264fa203bb7a42204a2dcebb47364c3753e2faeb4cf9aa7415eb6b3b38a7245cc086b45238;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc8fb1e46be14e288cf829273e8c9c5769f54630f9c462bdb25848721df1ead2de77c01f86ba6e17e43bd7ce0140892b3ae31158a217da7ae20c5d9429e779fc42efe6fcd88e007ecac080842a9069fafa4499510e7163a6db1398050a6eafe230cc420de878725e1819948301aaefd03fff376fdb1847c82;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1741e1d20b746d6a760435b266d2edcab9acf96f5599d6cf6a34bef3aed37adcc8dbd4632fb4959f54c8b40194154cd4d50aabe48cb72a83fd71eb4acad943f88978c4e9463f8f452d74f2117e9aeab1b9b3e0a1d7c1a7c08439bcfefc66f4b1da505b82038346fb7aab87f1637d9033000bfd79d361a836f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13c51ab4b9ccb7e71ffd5c728d11cf6604e6765d072e04a04048b867850b2dcc540ef5502420da0781b4c83a9ea738191c7cd2a8c3141044fbfc0ac8dce9f995ef6dc82c965352aa3dd8f9f100f6cfa750a73fa6d6564486ee691ca6c8d1ff82a3654dde418ddd7566acd42545401a3eac8ddd11b4c7fecca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h26783c0601e1789b45ff5b6ef20ca4746b7e18518f669bc4b2f5163210521bcc07afd45d10f25cba618864a693e45380e3269db69fb86e267c8262b4f10eb009bd4a9e89898daa24bfa3871360d930192224296847330f9c6b6c490493f30993830f4fe0f341aa5e5c3220ae293463b80ecffc3042b9e929;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbc3b0b435ac511b87c5f6df0330642c510ad7e7ee84db8ada5a0af1e8c386afd2bcebcbfdcc0f060980800977297d7d9c02fb28268916faf8efb6a8e361849057275d5ca2d409564153a1e559f0c2ed7f34d4100bc5d3f951b664c08db4f120c9a6399411feb5739ab4f7f2898d483a288c746454e4a5946;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h427e3f68c30508806fda6ac900523b494c7b8abbc8be8b71b464ba8e09c745f2f8f8de111639a091ca8c0ec15c8cc91259176c0b886c532764d7bd25a021846936bf07faa0e32c9587ed9bb97aad2eb358656393e609fa11ee91a3c5956a71377a06da5e1c4dbedd1cd1e678491651b1f78e6d491717c054;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h181d46def2f5cc913d226566834c83711b1b3621e9e116e03548d8c8588209df923e502239cab312464c6c2e891963d4007cbe07f30759e7675716e183bf7bd070ae80d10da6005fde125ecbde2bfb00bbeb9b24613db27015944f1e75163d0846f1ff3350ba8437f46d7db8865436675f4f22cab7dbb3bf5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13419a97ed806a9002c34d99480235212ae2bc49360b3862990fc10e920e0e030280d31de2bd9d141d328b1cf3c1bac5a81c924671edf602aaa6d0d157a70954130005b97d0cf79021250ae24af51908dd4b0c999db8e83da636bbd99229e953029a2c6502fb7977ab68a9adfe7c50b4e49410ab431883299;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h408da312988ad250895d4c1e99802bbd1e664d3870ab5de3eefbf0e56ced9547728a5c6118d05bfa89e510500784286d2dcb11c2e3514922c8bc58b052906fce8433e11c10bbefb4dc53909466d09df4286bacea1da3e8565e2640cd79216aec7014c4cddaf491a40890d647a422d955f1274c307595991c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8295016b4c3b46b62bf18f59ea51c46487da4da84aa2ebc9d98e8c7810da259b2de7a807658ed4db3183f45ff0a73aece824d274c8de3620b87465e6be570348c08833288668449b4739b2307fd01481a9ad6e4b99b0fa08177c17af5a457c896a43ace583a8d532c622cfbce88841151f1b7cfa18741e6f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hff818b0371f7d17422449a68fb205bfffed0067ec18284eabf9c51d0c73c948962540a5e8062e12174d43653eba6d761cba5b4d01bfd1a2f96bf887e105e16e802ba9bd6a96ba6ae0746cfea5b36c0213db801a6d28516f56a8a5230aa755e11769defbf04a9c62486667fe5b75201a228a6a7aaf55de144;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h23c64041a1096a1320987d6a980a595401187ef4b15f99354522eea4cc06c88e3e42b335c16c0b487d781027b1ce05250bac107b3fef85797a4212bde8b50efbb48ba69fca2782de695704f5c9ae269d149a68fddff2a78bbddd2f13ce1fa26f9f1e73185cf9ab8cd1271c0629a95b936f6b6db48654e9b9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h86770a3a29d5bfc4788ff99a7aa8fb5ede3865f5ad0a40051793bf316a5ac060a858873ec99dc2f462006f8de48818628379b8b848a2744f0fefa8291bbbdbd9e8477b522c8be71cb2ed88c2dbe40ec42fe7f960df48e736ed1f7b83fd22294b16152a72115f5bac8ba35bdea257c795e0efcbd40879a025;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h462986a2bce88db8bc0a6019f950fbd27544323ea4c1675e264d322799147d62b4791c28e9a53b345701dab9e03e4ae3033ee7986885b811b7580c721c7139e0a3b63149eb043748ab1db50b6bbc7a142c5ec36125980be8737c257a79aee7ec5754bb24ae28f0fc6a121e255f80d9f9cdf92026d28ed74f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h184a0b89564165f98cb758c6f606bc6bfebd7bdbece9e8275e341015eb1ccb7d8ba9509bd8d778f5e68b411048eb6c6ceca60043438756892b8ee7e22de109b000909370a4df028a737d4dd84ca1c0696c38eed82f87eb7a16b158554951351efaef6d30c810661115221b687bc1a8cca82fd93bfe1d059f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d18fb0253ad9a79c710a68fb121f3c5bdc1a31a4e0627a40d68c96013caaf51e8886ebaf6d7be267b0d724a9bbab1696f4635f5d14e0571957927809f91408f31ab5eb58ed873e48fbb965c05f7c84cca7d4dcd28a71e1800c932c9d375c5bef41baad7a7a791a5fb14a5c133449409ff406b8426bc802e6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb4bb9ebe7ca284b650680ab22a8ad52e0b256ae5898b28e0216dbbeb84d3cf30e5fac6e797d255a0b0af45805d583b590787c78e5e7d92fd1f094c9652f25d3a24eea5eb583a28f82b01fc525ed206aef6f861eeec3651a8b5251b5cb7d328e044d9445bc3e52314d517fd4e22438b8609e6e421a2f26821;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h68a99e98e3af609ac3c55d3b82ea47dd0de9d642f4c78190e734d907fea9d068404bacb367f1dffc8f3e4da5521fc0dc4ac0cc6cdcafd05d201e185d275121df04f1a4aef17beb087b964715d1ad4e3054c588e85468b3ec4ae2fd5d41cd40b0fce4aab4028a2feae17022a9b81e390f5f0a28bfc29997a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7caf9150a22a3de627869b00f1e42a7c7ec3a8638aa124bfd6215253b56d9926c1401eb872b8fbaca419195a99c700ab2f169400a7f19bcca52105113cc8b833209dff0f26e0ab4db8bfc43a3f4a6d6457a43ce095a6f28611c63a2c49802b4f94ddab15b4c2de8d3c5142e5e897a93e22e079b10c107598;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc712fba2d4d1e441f9d4ae7441fc86f667e70b9a095b31850e1c3d41e46b9b5ea6a5e882aed585288ed83b7d1afdda618e2aaf34730eda2899706bde56c5ff26ad46632b1105d64d0eda8cec14a847403109ccddfc4ed540617d0b7448ed03405f4f9caabf355aca4447a37793df08200472055cef577f9f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1277634f5cb046a2315b67b096ef4451a60e3e3d6658207ac1370b88e34b4be3d2a3fa80ce5978e8265e3325b585d2ecbfc6efe53754c6e0d599257b6026fa9a5ba19103fcae0fe6da278e75d8bd72ed1d5863e0ea8a9fe60e73f5092b3707a8d137ff87a7dfcc778639e0238413a31adef44f8d29e67a468;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eef88f675ad802592f8e915cb87ed40a36639870cf57054a6f6b42c1c1ed68a26fd202a4cb7a9d361cc24553cdd6e1a376d0710adc2eb7a9cec188eb09c8c3462902f4a24dee2c362eaf65a44528f26210dbd3d4dc8ebb81563dab018e250747ede615d6da44523718649e11b47ce342e4dc2428cd4b2224;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1764f2533f5f239a30028736ef2c945e1e4b2e5d88b5907437de404a65b7368c02cc5ebe0ed1c2d44dc9b9f7c6661d9b2a166b388a7d929bb90807f383ab2fcd4dedb4e0ab6b3a2613acc30d3600957c2b29a11aea6d4b0c8ecc5c7dbb6086de8e4ac39b777e37f91bdea25111e4e224fe5c2820cd4c3d8eb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bc8604ee8dbcb57d124835a0807c9f5cee44d646ac83188308c9952226169150656c89b561d5bedb5a4ebdce524d6ba3392499487fb6bb62aa8ded902e30bd04774e6b2fbd1a08af017dfa37679005de33900fba7402eb2a5a431de60c58414e5da682b7ca44956a43cc6f65c12b8c01a05f09c7f6818d4a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a26f50d4227d2bede1001f067a6ad9018529fd709fb4b983c98d5e52ed1dea57b32a7cb55dd2ee3237d2a565957b0693fe2f670b0c406373a6527089005e07ccad90c3a7414625ff893a598dcf5cde8f317150de03700322488732e1438867188df72e8bf76fd12c87d7b30367102535a3292c23b874cfb8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13140f0a00e516fa9f6c7132fd59388740da9f5267359b3138382a6a09ff677dd7259d7a39eacf3e3127092b3136169988054e20fff3766631987ae0136f8ffdfe5083141f1dfc1644178c44052434a2d10700c2a203a7c87fef8905089a060ba8d00f17d69f21ff8825a6959066a0477bdc130eb12765d1b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h910eabaf92f14230db0af4059898b8f7ed608f80e6fbc444ebdd90eddab34a55544fa2558911d5239b3acbd949dd6a87812845be9afca619663bb293d7a5cdfc5efa2810745c5d8aa2571ff17766a01b5081c9e8591c1d80bc753ae02559b4bd07a28c51f494e73f8ea05d80fe89945f9d0c97f437f66433;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f57e5fa70840cb282b0e038ade4c42978510af610c0ed25ee117dbe5b4513b71b36135d3ce415648a7acd9ec145fbda9ba347ae4d635d1b9ba5c56c9550982f8f79f47dc05fd06382f774f43c9cee5a38935ae315de3d8aa3b4888ef253bffc914be1d2a475827d607734e6bbca17ea7f8f0f078f8b24093;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfdb86992f8ac18434697e21017fece260dfbc738d3b071440dc282859d3fa6cb99b85fbf3a55f05c82becc3d5b426b48b545d42810b9cea54aecc03f40fd1d1e4f9a766819b4bbbf91d9ffa20a6db15fdf684be72e8deff02fcf68a7106d082000528954bc60c0efc3e38864491986dc62b664e314b1972d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dbe8fcd0605228db48fdc9a62a427e60783d1c41929d1ce8a8b6f70dfa02e1a4c2850fb0892a48433618cc5c9154e9e027e3de3acfa15f049267fb79ab609281de73f2f1ff1ed4222763715b73a23b74c12d88c1961bc3e45baf58f45d7e4194d045f0182077f3800348742a8a8995e2b4de01cd606383ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfb8fced4f00b1788d63652ba4d69cbd3431d01d42c4cc26757b3d4ca24685c63ac88219acf5397be187c6ab19fdd90f5b6905d654c04aa7ddaeff8edfbf0e3d65586bca9b1d90c464fc647f16e4161e2f787372e6db4179a7228f9c38a77e4bfbe01f57e49e7e48b6be617119e4c1807fdbc4da85121869e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd4697515df49771daf972c9f20e407f123582e4ed91191fd9d3203e5b630a036a334ac1f2988f599adff7559cb2145051dcbe4e47df21e95b614b3874924821b256364e6097327bfaf974877b737213c6e1dd1dd994426fe412f9eaf2393dd4053416dbe7b710c80c0d513d535b22ffb21668f5232d35a36;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f2ae9b6ce5323aee0501e32957cd787b8311e676d13126ce4762483edb8fe10feeb45a11e7cd6a41db05212928c73bb5e79011b182b0c265a2b9d4fdd9103d1ab3d8274525bf264654cf1d11b133bf4d42be406e1d0f80b83883860fbe092ef2054286815388bee93da7bd30baf7977605018cf9e7eddab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e9b8361fda1c6b2faf22881ceddb246dad021a5354963e1cdbf639e54aaa43b40a1c517d457405f0c14eb58870a6cbcd90896c2e01bc09db7244b0bee718fd59d9581f73df9f059df0b379b8b823848766fe76fd90110fefa66c9a3760c0a08a56874921b7a7d48aaf78a1fb6d8bb2c63ab6a450539554d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b818a82e75c79ce25ed6913c73aaa7ff7a60f6377eb4d1e2c794b83191473ae7c1c697acc8ab3932a7dc834d075a8359773295c8e9e47ebdb133cfd2081a214c64530dd44f7682209a3f91c39bf2dc43b89785ebde40b64f8424e3ed8ab47a944d378b087fb4ff7f05236824d46ec66050b07d0ec7e6c7b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h895bf952bcbc2154517f9bace05f44a03981a042905e2cbc5c1c71028ec1dfe0717c1d4a831c40a792d6b232471fffe6e3297ece8428254f73e518c8fb8b913e82bd0266a67d9e9399a046d15416c0f1253ff700ae743257ed79dc903d65aa11617089d79b25a55e5a1b3f75768295bf8eccf4c4bc1e5d1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6518e2f397371c87d844e8333db749d8581a2fb1ccec3e82bb394099e67353e49c2beb1ea49ed32a26042797bba9c73ae2cf522599e91bb059fbc46050661d768cb963e3bc855aca8ff8650554ef81511e5e6f48ab3d78336641784277c377ab0796e531c65882f43586663605f98c96bc41240f4a53c22c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha7cc3088595e9b41e15ef88507d25d911f51c3088f4fe8390263adc15c0bef3699d098a21517f96c1e4a50365dcfb1d688c36f6b38aef12a3931e7461000e8a12fb634c5c93c44125736cd9eb6f202f66632cba4f2eb9338ea284b022ebd5854c9807d1452391c3c609708605ee50aa787c4b3d8b242745e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a0eedc47c53b92b298e46166a98177ea2aa7c70a3503abde067a6b15843832d9012628f113c3b853ca473fc98a57f68de046227dba7a502e08156d7ca2bf785656605c82b3ad1a95474843aad1f769862d8806d2805a812a628ee4a46ce7b15f3446db7f19be0c7fc5c943011e528b58cc9cbba5216e5aa9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b8d237203b74e9f3e7c2bf74187a5312a54b1e9b680022658f8cd0cd0d0e8bae55aa73f1b8d40f6ef7c8267c4fc39df576aae4eb82ab3ba83e9b580d605ae4e1e8554623dd58d3dee5dcf31b0592143a39862259d27b3b58f4192365c95a3091834c28bc3f1d4e2757c8fd3af3a6a485625b08ca402e6f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc3c6ce5f0d46f2f5d7d00ed195485d3f48a803f7ac8ba175141780280f8a9f1ae93bb6099edb388a21f9992c8a538d4641804e653d0ebea1191b24bd474f958c797db3a8ad3a3bddd6aabec7e54104c5daf0d5cc21c96634d0e64d4bf39e47b307bcd554c81b7792e4196ea12ef61adda29e8392b7c04da7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14af27e9092a71a2714912dd49ffdb60a7a868dcfa6376fa8a2c15dd8dedf2428a08b54b8ea8236d2d852baf7f0408b741d8d9762549bdec58b237985604df4904cb90a3b21e764a950756fcab42169d5a4127b24b4af2bac99f3b3a178937eb108a42b058a509e78591882f96ddd24ef2468b8ae493bcdbf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cc81b0c01416a463bc2746b915d2c39281f5c349866f0e15ef976686ee33c88ae8f3696408285d9f9ce9ad76e6b6a38c57e1827af38494ec93400cb7314c995bac4c93c8358d74703392e222fa6f4ee1ff966c2b92df89e42cf1baf7a24595932e9bff3f9d088f108f0f1959045ce0ece222fd709cc5d1f1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12d6d727c676f99a53da6021b280a791a8ec42277135f82c3ee6158c740800640773a8ee96b60be1a5169f511c9e7383ee3719aa65b99d6a5b5178cfd94ea338e1f83ee67b1a2a84a25eb7bb07539c823d6651766b8ceba80ca77288e11e1571d93a5a13a471fca06366ae7df038c0bcdf3287eac6607ef8d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3d43d36e698cc00d2f1c4c1f10550bf114ba18eacc63fbc3d2279d239cb74081a9f0ce9df0c35eee6cf1a11309c82ddfe40bd76a87d95776b85d35555e60d384fc816f56315ab4b01b1bf00c637e5449109a20888987df46fbbd2d58631e751a9e689801d77ebb8c18e850d8082bcb9759052c9f35269fa2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fe2a97014c278705ee961c7fcc4b504c57e961e9a32c6898946e915977c144c1a9e8a249b558e77a12f68081b56a302ea63dc98d64758679fc01532ed777c7990e8a478e618bf894d0dad56abddc5a1f85341934bb16e6759112b699eff3d48eced4b873d5421327aca70fd1837b8bc854b6c7f5f7086a75;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b44362546da744d551c54970ab42c8bf6a5ef275c999aadb1f2d275389ba8d224ab2ce1c6c43d0836111995185564983f6414951a0ad5ae01facf95a3ded0fa4282eb02eedb43fbcd9cf1f0eba68e940a100508d49d26c17ead9d5eacee0e8432397b6666a2e0763cb2460fb851f6f57106f45c520c5a6da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e447f383b4f9842d9dda6f29699ddfe9fa6dc2cc209e10aee0ae3836aaeaa0dffc94234448e0ffd3a38f48cc4569f23f9caa12196201ddf2942abf88faa0c3219b63452770c40165656a69c9d9c840b817fbd0f4536b351c360043af7937647b3a8ad8063f65d9c1192bf318691bd68638efe4467747fc68;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb39738d0a2b58352255bada24f02e7abcffa81807f55ed8af76531e912887b86a7c15fd23461040c42830f221c10c3e556c2ae39aa7bf665205a55b8356969fd92e875a4d2f3dc8ebe295463f0626a9a1de66b9c890c649b92a99efc4bbcd674d404efd23e3d039891ec2f6130b81e87478927e3d4f06623;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h33bda676bc1f9305514b073f1e278cc7035490dd920c4ba47c246c2c5c3754ba928d21b656e813c76cb7b52ebe96fc7f9b82b9555515c291342ce6e4bd510a1051028b6f26dc83199b68cd3b39cdeea0f0ef418df3728405a19343413df23a74c20c64271d022b4c4cfba62f19c1fdbcf9bbbc113f36f240;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5ca2bc036d9d1b19c7c6589780c34690b7dea5b5fa2c6794d6a5bac38f4e5813a305c0254a7a538c1356a3fe088938c12d46ac27cbade3b9a827479b763f4f4f4c3c4bbe3f4d49e17aeec4b8ac5d0a65541e5f320c3c2287b135ae33681222b3d08a136a4eaad23631a09a60b04703171994ed234677e019;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd18f26d5d6e4623dbcc9748fa7aedd3988103251419ea9cb41d0e621148c79b6ccb400de1cc8123ded055fa184afa76ae0d143ff900b8467cbfff827e42681c41bab8bf28818814066d2ca447bf0f21877c85af9f17f745b1d10d4bd85ad1ff1ac1c657f97a7ab4d30bb9b98737044885a4ff0bc11ebfe66;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19ae779c8cdb2e7bae8c7dea3649cf221534750396bcae498d4f8abd0b5109bc748bfbe3d050b6ac920e60ca4321696bb7cdd53e0caff1fee28ce87c1a678cda280c99c06f6210e31ce3f870d8f1b3a3e5fa01bf1b5816f2dcb5d29fbe01b37c60adae9bd404cd99ed30a4aba70068b5e285503eec3b63d5e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e7a6adba16848068744bd117ddfb537a0b4090e630f45c44e62c446311d81e97e35ce23c6004e386370a5faf6ca694aba8d0f05a4c4f0f33bd9f8bf1ed48a830de84498adfa7e48710abfcdd3d2ab6d81877b972de8f87094970dd13a05286954d8c4725d3dc23b3cc6d9c6f25b0ee0d7d625f6ab569e5bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10377aef5d28b98e5cb33649dd9ede612e8201fd163c282ed56da3988017ed18fd2bf4b5b76b2e4b066aac39c7f881fb2193ec9aa6c026f35edb5defda20f627b16a2366b2ffb79a3761bd76fe1bc9af60a2fa940faa137eb712c62ca7fa959ba337456fd00cfe8c8dcf792a5cb752572af897e04cbdcd199;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2f18af5d5d4a7dcd5aa21347ad9c7269deaf82d1a61fc76066167083f2d6295de64046cfd70496f49548044759327647da3db99b1e5e3d19075b0fc0c419a735782d63b455c98b960b725de2db00ba6fd4462005d644d9c4242cfc5bf266b016fd5f82bb2387b93f9bea3d3943e0d32042efcf66c0bbfae6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dcb53ca47feccc62b5bd6402750f501ba096fd9780fc75a86928b07d4a5c0738479703ad25cab28f7251294393add013450aee3ae1a532c09ecff09fe77cf74b4bf3592873e69ae990fd95056f70718dfde4acaef4f53486df32c6e86edd53fb39b38e7931e5b4c3c3c5d8e882f62fc1c9ad6d0a3cd20250;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h160f9b41d5e0b061d50e1b63de34c77ee5ed8209ee15c4e1404c903cf413917c3b8aebdacac7a5f4f1e153b52e04f7d1ff8bfcbf4ee81829804dcca2001186d2fd76f55f04278720047384c8b3fa338b8589ac380be65b0969f28a29d8057c8a6073a1a0514fa706a2738a9ad5241b14b7895a98e6828bd47;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dbcddda31e3099156f7b159b894ac98fcfc4c3f05f1ae0ae883d7ddaccb2db26d129ad196dd2496c04363c7460657b8467b95a046d7d7619ffe37d6af38024fc9a9634c08af9156df684201f9ad099f4dbca5822560860fbe8f8910ccc3b843e25a9fd6557080fd1eb0d0ca19fa6ae71d98ec2e53bb5b24a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fd0acc6d96f8a23ac5f3dc2cb2b43feb338e53af9da41f481779306906f4a92f2d656d3e3978e0e6b44d4769463cfea789f7816f89f9c1e6f4d89db342ab79a60de4ffe8ef8fa64f29afb8563247fae16f1347c3a9f27345881804d9923ecebd2178e1b39cab46ce19ba776ad0771db39e3e7793760da971;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h150c6d9cca7d6eaff69b6e27373f74c56c0b5a4cbbbe11f98e678dc786563d490aed65f6888954b2cf96a1e510e8e58812b3a6a2c750ce64a4bdd0c7b3e477a7dd28798046e5f47ee87f29c46130ce8fd307c2c085e9b977c01fd2aa22ba75ea0d97aebc661c0205b4aaf9e9d1965d74d3f7e0c1750dc8c78;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h33f6a9fdde4c6d4c62263a6f3f28a692c2b87f91385c8a0ea86e88181dc882dc1a084b9ac617d0bc65f3cdd35aa24c6491a5b993dd73fa4ec533816d9b87903572c7e6a0cbadf0d321a7bcf75797956e285cef2c1d7e78acd59098c63f4ed64876c6f3d05c2d2c07f03cce280f1e1a9185b53fde208442e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h102ad808b5fa71638907fdc5464db4a8299fc0572e47ab699bffcec6b72f7eeb4dbe33e6aee6798b4c567de4b9b285584eb9798b958f149c345e670bd3253517fab827c4a0820005ba3ffb16d747707dfec0d9982c648b88dc73fee8e68e07a9b49a610cceda1ec1f313968af74d326a772300e023f8121c5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h29488da2334dc53b88826fbb62610ed35daf87f44d8f7f9b65bb0c591fcd11c0c3dec428d8be50393780e67de970a54dd926e02b351f2d9d825e4f78fbdd265739923205c405ba2dcbd26ce3d1c5545f27312ec87b43efcf3ce9fc3e940ccf23dcf6fed63532f5c28e34868168cad03b1700d6e32c527683;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16c36a42bb18a90a1be08faca0331f4307b222db34894ef629719078ca3af745e8a763df1fda8e025ac185b16067ca6f4a043f76655b336ccac439139bcefcd34e3650c7abf04842ae9d38a5975e3a5c7419feb693e54f8d9dbefc07ae062e3ab84260eea58ba676fb9a92bd4fc9c0d4710684670d0f59338;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he9594ad335dbf8e51a71af216f2f0d43165ba6d41fc55219bf33770e29d256c5cbd69da82efcbf50cbf4d5a9dede6baa77b18c590f9ffb9171f70a17773e955ace6498d000c8edbb24ee60bb26f7c5ba50648e3ea0448182360d0451d1531a5a3066882a0801b5b2a0adab4c58a15c03f4d741a237ee057a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17092e556c24ada03a5bf8d0bb8d8b788020eba883fad5d185789e3acd352f88fbdd686a31152108a0369d84288753e8c5f196fabfdeca5c7fac29480803ad514aa775dd1b70e4788c9939be55b11f1fca813690b45c66a519b5badce688450a8964ce76068e301802a9a1f9c52efdb7d2166d1c84703d45d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h260c5d15d1d762e28fb7888f8dfedee09a154e5f6ab0c94ccd45d5bd735f36ff729c7eeac02e14237ec05d777997256cdd06aca2934dfbe4e957d8c47ca810753136da38fcc02345b79aaaafd501a0d1266186607f1bc20f5dd9164344b7b54abdf1e7f469643533a772ad7a833edc78ffba77ed95b312bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1adefa01adfb6fa67e11b163d0ec8f637f74b388d6e4bd8285be1bfa629e8b6dc4612d2d31e61bd2e0ea27fdba91259190458c85229035a50fe55d33a91fdfb555d2c6b8530ff0eabbabd9e6506e01f93ef47592db8a324aecf2e7a70c3b552c4844d74f9961b5addb22d26e2bf7d4a92c2e74255c7046211;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha721edd99748559c380bb5a5b56a89425fbcbe4caf5856b47849cbb54fadc0005b0665a656174afb6eee590b6147f96780474a31fbd45d53771b0fcdbd8c1f3ef86008cdaa1fa13f7f891656738d5244960f229c558a067cefec86992344d6c4665a9acce8932f81a95a87d51fd2a2049aac3ee4af3b2bca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6687bd2df0ca32a9bdae3ce2049be33a70e6b53cc2895f8e55961be4f1babfa536223e392f72364c1c7d434a4b220a784297d94ca8198c09785a4ec87d98439e5defec13f0e934e1729fea79582fe3e130c62170762ccaea64f1bcc4e30eb41fa7928a03a98b42ae3c710c5d36f41d06e513a3fb99e8b611;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8946231861d48f4a55a99f9dfc9fb6991e731d5607b0f44077aef94a5a04c7d63b0cbfef41f43cdcfb9df9fe1ee5d46058f6f374e0fc304fd7be702f855e323e02adefa5f4b703a87e1fda8f5fbca3f95feec00577c47ebabbc0cdaebc5f0ee9ef0f2e1f6c2df7d023c54f626978855646a6e64c3452508e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7d67a5253bbd20f07676c9c19b295e1cb9ae568f7f3a70b372a049955f69f2382824c1b1527289f6087f7a96a63385d2fea94e60a10b251fec371e7f48b383cecc1b678f3f0e994842a131d1a157bd0d41787319f67394594831f1628cdbacf6c1d28581db76ac7118f51404d33add15ea6e1ed6ebb5d42c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19c09bfb33c456ca6de655f089fd509b6ee6a31ad159ec6bdd49a8ff8dd054f9563e6e088ac26a369f8f32bd9b89fea177fd335f9fb352c59c3f4d80e029ad07220138361e8a7f044147c789783b7325656ea3ffb19150bac0520849b24a5eb9cc3db5f5f2e682d2a0d5a0c1348ba208e9a613ca5159d2fe7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he95633c7dfa74d4c1cfb3233e987ebb9734af93dcb70eba3e2f8dcddc255aadfd5919a412cf002cbe16e7ffc89677fcc2bac89d01386e91a8901922375cdc4ba7f85a376b98e193d834262ab3ceb99a23a3917294b332ddf7de688d2683c66ffb6f58986b07b4af1d0856c29b37ac5700555afa9cb71301a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4324fcf9a910593fa102f9b8c1f8998652ff381f0809f6f98ce99acad98e65dc219553ad4340f3d7438e71ff6b2580de303268e988be35d9fc40662e74041fc5e14f840efd14f073e1a3235c00e0965d7d07988d05bf81525623a24a0a739be62e565a88b4276fd7f83dcd06dfb874fcb12ac10b38b6a5d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17cb2c165a6ede4efe4ebefdf6763b4f291959db6dc98fbc3dd9e5e29b795f2a33a6de3c3f8e3bf5253fc8b40b90a01709348f83f37161ab79e00d577926d10e04e7e83134f688dc58f0a29fb70869f2baa1e740ed0845813188355a040d977f5889430ed68b931948e228b4f902bf3cfac794572be9f7a4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he40bba03c84f2a29fc856d2331bfaaad4ac9d03295b85dd52d7a7ef6f7540dcf6559903894c5840bb07c096582fc7a9a021360a2b6626698a89e20928cefeff3ce35a89349f9b4d59ca8f1debe3c4d56e68786f380550c38720cb13986e39836bc1d2b1977f92e595f98496ca9a1e765b94f38193588ec5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha187a4e1f0a0565c1325882908ce31401f8e5d53b8b5ae1196145bbe2c1eb1c683598e53e4bde604334513b483595a726d8e11aad606c802e387f44114cb40f0226582da3b3ccd81f9d039c7fa5db457e3aa9dcb580cb182d8fe2ba1cac2fba09805041f92aca796b3acad61ba10137b7eab9fb145629977;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h193ea7053852083becaf3bd1b50d66bed7abe13300f5dc0c7924cdbcdc9eb92371cd57aaa3ab6728df7ca77ab2c263db91d3519aaf9bddd1adceb68a2baed8c0a49e35732cecf56f16cdbfb8a13050b20525f5bfb73701e29b3846382cc54557295fec5fee276491a4b7d2630f83b139919a92a9bf87937e9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e58ec07ed7a2f19c387dbcd8cce158c6e2bd17c1c70f947a268b97a11a5cb4bcc2bd0f56e36ae4e635f31142614d607bc93f0e9ade0c70bb4c296818b0b12a82da23afa2d651cb7cac4c45d48f329d884860df062719280003ae7f42e359530cbded6d1201c748d3fd5e3b6116a33c0a700ca7667d3f52f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h78e17f996d67de3b32c33765f3fc2160eb5d0f79da463156a73c79fbf8e65882999b7487e1351fda0ecb2723cc73e4b60415a9e5d4a8e48a15007fbc184b1bd256fa9ac2427a0bfa62335ea415bc23aedc14372b08d7262b659fc58f70cfe44ac204c34e90d7c3abd87600d118ad3729e213fa8387728850;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h90dbb2431acb36fe22d7c6640e369c2d4c8eed90ae0cf0e61f3fbc838e295f372439e5bb7af7854c1ddcd96329124ec691f96d55d0a24b920046835baf81e19409bf6623a24cf4beaaabdea08261c7345e896ba8086402794499b0367292be3bdd01562aab55f748894be4d86afa52d7abc0ba7308bf59d8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10bd7b730fbbd2068d10fb9c28e789fb0fd220371243ca5bf174f02763522522846743fce4efc9604dfe62735b1189399962814eb59ac59c23bb9e194b52c03ef917926f6f3445ab7da93c33e4a4aff5356c5033c0d2bd8a5435c8413188e1afbac11a02600e978e916c859bc30e37cc82933915881872d82;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h108348ef612f589ee015bef59a90ba565e88cf7ff6d13083426861710055a03e28d5e4bc01812e52498b188d9ddd881bd4fc54b9fea85714f94eacd1889bc548ffed0c4b0f589475e008a661232cf62667a9637b15e4e10d1110761a722e9f1b64632676a7346da9fed9c7f4239a7f297424898be2d687548;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16bab687d6068ec579800b1e8054c77743da04874517c501f95c6a385342ed9de6d848cc73c28765f3e8b70bda740dd5c66fe6230ac00fb25ad1676b3de3c1c40095335f7f47472ea19ba7495bcf8ab683c8cac210ef3b3ff421dfaef3b0e991b9c71252ec0404d94f0d7f2ad54435a16a02e00bfdef982f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h88364b845aa81eb3aa87426fc22db2b58ee3d6b93ebed65366653aa400fb198e51d0baabed708c09e8ba8c4c0b21afd1c1daeb0f4dabdf99dd473529484d194bbcddefa4ef9152334f051717219aba1cc4ca1c1a3821305b37f21efb2ae5ede105215977ad24532894dbc6ba4f92d271b8adbe1d14189440;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h113e838d8f4f1f0e3a39ee6c937b22a326b6981191ff63a42fdc897beed20258edbe397eaabac978f39139d5fc870dae9c077da6ba0c8b97cc9ae80b443dc2d540e86c6349564d4c339a8010837e6e2ea6faf7116a0541312c3bf5fdb0496c394f4dfcca191aee64348cf3c8678c80843810b239a81eff437;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2a557f20fa7980194a5feee84de84f0e07a376fb3f8bf744504d91eeac6a6ec73a83ba211db02ac0298bf7a7fa6a2b2533d94a536b5126a4cbfe89fa26f2eb3f5f636bff13199baffe3db71bf4908ec11535acd4129c065dcf37fa1677c6262c5bc61f2788b0ed1b24d96acdfa101bcd1627292c6eb61c50;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfb43bf61fddc7b340238b6c5b038444952771f872cf12c065d7698c7afb923ffe9abe2f28bcddef147b533ae2b735eee611bbf81af311c0190e640dfe257d9a3f19d53561d1cba5c86d9a16fd83db4106dbf44b4800061a150099bcf6662572cb0fc001dc035397be6efc95734ad2c32317bb57e11a4d749;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e2b9e66658c914ce622948eaeb3758f1c72fe980b1657a8f43b191ddffad3c2b4c5f1230eedd4ab6f274e44709f2bea1de65ed3685c0c2afdd6b1574fe9327b5452dd7bca8f2c13cd3735a291a7f4cf4d2393a25252348fdb1219b55d5a61c57671780ee34738b7ba2d1ce5eaeb153eab77ba75b259aa46;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h175c0745ab8f0c439969cdccf0215afc87d9409e6269b00fe6196de0c155c2d92ae76307e0897b6c0a2cd6fc786623382e1beacc22dd5b72e1fe84a3148fe2a66723c381c6365b260f055152d8d8aef667da9a1e8675e6b0a3c7d52b725dc7e7e975e3782b7ff3a9ca54afc35b1054fce09c58520aedee6ef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14d288bf8bde2585292c16fb7e99f790b7b2de80188fd1821ccb1854bf79344eac2663f3f265162495f996f851b2b13e3e9766f0ac7d00cbef7127c6d3d83e510b67870d3bb8e5f31cea2006bccf9dc7f25ec663ffa23d81cf4cd069f120738cdd6c5d63d6ef0d18235194272c13509825f1a3888758f8792;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3e6f9b111fda1374c143fb8e0a20335ac5d462ea06b18b9f727d52e32ee77077abb3307c7a95b81d5b229e7098ec6fc846df5831da06aacd1bb166ac41496cb15f5fe5696c72cfa507708d3665c689176396cd6fb81887900b72d0d0e8b2a6019526950f49000cd03d4cc8e6263d1df69a0c63bc408255e9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d009b240e0196f187140e0a7f528c2b2b79122cd2555fdaca90b66d6cf8d41d7f2a06e80ff3970d3091c9a788d6ddceb3382b69fc7a742213c9c210d9f28eb898c0e07e786218ddc22e1c58676d68b28f4af9015e7ab38dfc8fa8c186b4fa518aeb778ce82e420b954a12d4884902d43ffb76c91f040bc76;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h462f42c04e6b959c323a032a89f0bba74ebd1aaf635893ba0a197a4b47f744d49d51a999a1b1ff4726f65a9646070233e4554c61570e77f312b3e6d69460c7f0781619a826c5cfd96ba8d0f37e9c2a3cb0fad20928108b1b1845479a81f91ad3c175562d14a38e63b0a4000323fa38abd28c5db85ac9c3e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haeeffd8b066a075d317b8cb1bca2c433f30a513123d3d30f04c965ef584678b0df919acba24072667fcdacc039a4946cc9acdffe4654115bca81b47b7029e92c7cc1f22ea8669715356aa47c64729dd7b60444bc9061a36fff67a83929e6a0b0c0f8527fb896abb4dffe9deaaee904e55adc7de75fc24c19;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc506362dd70fa6b814f419cf0ebcff059d4445505b929e144347fca955ae3a60c775cc31b6752136f043b1665086b12a49c304e3d38f99d53ab6b0a35ce144519ca432988713676784ef07f12490e25372b04fc0050793bbd5a7c39e43aa863bb69689b96bec90e851bcb10094b3a52d450c3ee0ffd6b79;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bd396da33179770cc50667674e0f1a81bdebb9cf9e8cd3bf702bcb05dadf4cd0c50cdfd4cd40fa95faec7f456e890b5078093fb975008dda087348149e4b5f59127999f895f21d4f0ab99e0849d62804c5c7036d10655cefd6547cc7867c2f997bb4676162f48431325c3a6a8c6e322fce408af782a6744b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2a675e3964bc7c5fc5529ad58c80ac3663c80349b187a28dce8339aeb09cc3c24d4f6ca140024228233b8a00ef13728495da4afcdae2b8b3409f7726c0845283c5884cbf9a7f746c22f9f02b5968fe7f5f0d70b6e867b1d259b5ead067aebaa3b757ffe47b052ee9a21749ae0119d407535599860812cfa3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b44dcd1edaf1b82f8441077b116ed6443f50d34d79e2bdd03174d90b252fb7279e8784821e50dab4a3601a815e0ada3213c91368a52f346cf38b46df1faa06d9bf2ec5e16d0556638262e089fb1ec447c5e939ac91ab3f637c7e2115df80510d1558cdd6f0371381178cdf753c9172179cbbf4d75fe2659c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b0929af4675142dc9807c1c0f5aecba118432083c2720df6715d0fc8f473f4b85890ccd2e6363f6512b5a7360bf38e78dd26c8fbab2e5bda6100404c8c69a7eecd02a8d3495f136c3cec0cfbb35234d20530096a5fc5abba1376106ce80c6eac486047f7b09f19afd2d463db35f3a4036378c27bc63ff3bc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h33416706b3e90067919ba99ca53b8660b745857ec44806c25254d721289d30cf7f5d57112f690a37f2515a8f665399973df9f419b50ccdd552491a1da714d8c63f7370ee662e3212aace39cf09d7f2243a3a59a42703ac401144e1e4c7f5f914325695d0429193413f4673a37963c253fff4088d2e37b443;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3877c832e1a4e010ff9498e1fd5ecc4dd6a4d5f6445f835588acc58cc0d0e381c25f66970c50a879e5fc2d3d386c197ce51f75dc5c2191b08a45f845de86319ac1d91211cbb80e66f8bdb3854eb92cb48505e2f20d04b57ec98db3ae9e18c6fe54bac56f4cf7a1495089cbc5091f96bb2a162030a4ce7df3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h634fdc7307e7fcb6ec171964364cb7b4cf6c2bea9fc3a7f19c764200e850566a0cb25e5220b7ed6acd8e6c4526ac400b67aada0875ec62803816ab65dc5ddadd08b429dd31eb90c98abd3193b6476df5df14226bcaf5e7d86513824133ef19fecd7bc3fcbc3fe7b01e2a1776235183597e342bb9d783d2f9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd6cb4c16208f8f9b840b8eb316b3f4b33114f15bb3f4c87014b01e1f30de1b48cb82b641f5e2bddf8de7275a679d861a4eb4a381e415847aabcb9da4f02b3670176f82a07dabc3589c4a67a9f2bc20d2ef050d5be7264902e9fedc73174d1c6b3c08c573cc817cd76134bf94599ef0e50f11848ead1b91e2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7a6f1f743823d93c010eecc2be060a0f005fd843e2fee4fed7c8259334c02c55305e6439b659fde9a9f83e5dc20131a6d884a938395e73eb5daf048c42a2725f1f05db788e6be1c2370080ab59bd2d1a4226a3a3d7ba814a7c31fc4ff788dc9ea3435aa70db0f496cb045c9919358554d1788398d9098ddb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf82c468296d0701fc911621da561614003bdba3862188bcbf8876e736ff0530cfe3e8a1b9f6381c26d8979480498b57d81a0feaa1063bf76c454de73f73ab78ce12465befa24b54f008ef7218d27f69af948baf8e873f80bcf413ee06a51ece9f045f0f817ea111b58810898a6fea0d0e7143f333041627f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha5386e455d674f306e2dc4df8a442505bf6d486f9efe1c53139b790a4258cd7060dd3b1b5de765eeab0f027592581c4e3c23dd79bd4d70c06ebec57019cd8f801b0848330c5c0f0877ded9c51546d7041d1eceeadb1336a684497027ab8211a15faedbd8467fe7c29ffa3e13a1c5c88cb36f89bd9e2ab166;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ab502c66c96d646ec70bdc9860fe1331763a903d966a3c2583c96cf8a7a39cf53aa5aa23e06d149f17e71be0218c8af712b9d015892ae7d2b2be2897f7661e148d919df0f578b366587c41d6a6d7df1ac3e1619ac0eab9813d266d618690c2db980947c07510c8b145e53165f0dd253749187214c3f97a4a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h69580f3803792053218b097349dbdd6e9952ae127590a849a7bf6b26ff3156a742ab3c5340e2ea86845e266a9d2a802caf937efb075aab61d390e113abdf7813a05208217f93a0b83f5c36e63f38069a480151a480bf2e4948cde9c1b596677bd721405a4287dd297ed943e002df93394ec865d2d8ec7a04;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h604585575164e126faace17ce5a8b73c49865efe07e16c29cc5e754baa84ed525390b4a760e957bbdee6eb3a5dcd64275619b7ded2a983bbc0a405a2f42ca4c7814fc6905ff888b5c38c073ba865c1f7d3f8d21f817fca9b59dd3a966de6812acf945efac87888fd14fea138600dd6d05882330e38c94d79;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10164e057a3843c826b7ba41e647324115e989b006f6780c78b8ce2c7cd2f1c337e68605296cdb50d5dfc3c8523be27ad8e58d095ea971be7e0af2a8c600089d667828f4e6e1a71695fdd603ee046e01bb14d07fc7f442a0b3dda1211ca5370c831bc5179ca5dedce9cbb9c904eb071a3888cd9d0e32cbaa7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b23199e4911ad10002f8200a4976f8fd029e143a5be48a8b10bd78cccaf79cd5b002faeb07bf5630fa5c08b1492bd6d45af4d71590356c975e19bb9f5d89fa890789974180e2b2e47eed8c68ed13737c9ff3f5726d2a7d4d5721a4a2b8e053bbda08fd16730c4ddb80c00f718e8bffdbd83c4267d23e2be2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4de98e62178edf83a601db22306bb3060bd95434cd81129f766f3d18c85097085a12a527b6d04d69c85ed0498b3d00504e405b1984eb04d455a889973c9a09af4b36cf979935530ccc77efda864b57701e4250b0c86a3ed170d7c7bb8af640fb4675a21549dfc861c06062e23973addf2aadb48c94373c0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hde07a05c0924ac8ad601f830ce86886ac7d8a1092f76d2bb454dfb6f299402e3a055ff0ceb6d800ffea459ca6e3077cf0fa8e2039d814e2a3bbae734db050dd5d5b15d038ec88e74490450e6b7e98462e2e148d5705fe1d25838ae31fcfe1c97891ff6d36b3b007911501f1e9e1683e14973c1169719e4bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19697d9041c308841ad3183308b13766e6e9c3d5f985c7b58acd6a2ea691b1c8d91fc67089986265473a4af5281781730daee70c884265a833329c112579113eeed7881abe7409e5067f383870c926c27f48398f9110e9b04db2983074c5f2451d0adffae8fb01f019dd9fc961a07bf14f4338c5336d864;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16dd5e80320f0d169dc6fcc3e0641ee71ddc2088ac2f8bbc59a0f84a34f8b04b0ca27c391f284812424151b4e79db88a446b185157c62b4112b529691e7ab6a56bc6594b3525bfd8da33c0cca0a3a4564d898dad1e07f051e684667b76ddcf77eaf8d189a2bfd547a8aff330699926d45aa5ecde7e4b100b2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e18e4b1b120d6d2cc4c9b56c386cfb15e1b0efe2b7ea06022b3242e07e933de96dd8dc05239dd94a0fa0e817aeff276cb4f7fc96b863044b4b919f93c2b6f298c283940e184c9ca4e7e16e56361a4cc55b913b0d50e3bad0babed075742d09d58b59d6ba382ddfb5671715358bb08a8a7cc0fdc6f05b661;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1123c3e05675627cb4f648e7dd8cc71c17aa273d88df65b2c71d58a74b6654880f0ce17ae6e7c7f8a5f6c06ceb6c80707eb549c6952b5418dd42f11d1e55eda74fd959f7795fa93cfbfe27f9c3252f1fb71261629f4ee11c3c5213ce0361e7ed68068791647017bce354473f01cdb64633638b8e8ef5aa054;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b264fbe0b6129fe966894a5be3eaeb77a3cbe3c560a7807027742325209fdb9b65e203c7bd269cd78f2c42a73f0690f8667ba912bf619f5ebc366000ec031b6c469394554799cb0033b5a2edb11f2534ef853bb14a06774e6c2cf866e5e6bd0edbdf006b9a1ec0f975508f0cd0128afe2071cb446a20bae2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9f5f03d0401b963fc66786325e8189b63c67677d36486fee178103b593cd695f0a157a9f9384f47502ec35a786796912e5609da9eb07c8f563addf09eb1d753f48f22ee1e7f87116fba02569c9bc988971015e81f5589d6f03869c054de99b9c0086c9205e4a737ff1d4666bd9316600fef9ae923e25bade;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfb87a08b23b1e43d75cb862cf14c38e3925d237c56db0690285c8f5a05b3cd83a18f68abf479237187aedface19162348daf61e452b951dc74aeaef0443492b8626e0ad0c22ba84ae60519fa04b6a399eb51e1eba3573e591c3e50f28761ffc5ad833aef727210e3aa1bfd675f0510eaf576cbfbc559b2f6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4233878eb6cfaff44db1f60043865db99b6af00ba7c104a1d294a7ae6a8feccd68766dadd6bb706e00bdc26fb777af4da9786319fd6a89f868c227a69a85c9e56ccebe13fe3c3b011a71632ab1d561fd605c677b8e0e7ef641bfa450bac636ab03003a1e8094cd2d16c9f73b7e6fb734167625b6a6ab9664;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fc29efce12a1df198c0d235660e3f5b62f6f353b08fbcb5d4bf6b12cd02422ba4256beba928dff17e52953997d4fb41b5205b9c6792a924898c07016da4390729cc0987c0e39baa64f36bd065aa02dd631d4104269cf1780b867d320c057d03b5c2c20e6165ffbacfb55d5169f8e51d5a75dcd6d5ef107d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e526de9dbf823e09e84cf5e3546ea9edaa1a09f250783ecea4fef6420f502684872b9f9deec43ad959abcffd9992c0de54648a3e1eb7fd85fac6ffc236e4e7166a9ae143a06c7348a3f97f6616a18d3410eec54b102616aa52a1808a87d9d78082983f0a84065468d77b691976a5b6e5ca55d5380cb20392;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hefe884eded34ccc354b5f5a4e1c819699a2b3238b1f55c9fa12f066653edb23771c3540ee882cfca5b68b26e8990406db69240cd68f0d6f67b7c5f74fa4efae5c883128cc2dd8fc3132396d0167e75390880dbbfdcfbfd49d9c3d4e68bc4e2c273170217068ac1a7c2fcba256f7d1a74c043e312605af2e4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h370f888dc532c5ab4044d3020ddcd3b3d2c9e093dc069a2eeba8fb1efa81d4623a5312aac1a99e37779ca79087963cfc217cdccf27b84fb8dc6581dd37927d4ab67253379eae71f3f3987b02d82d8a17f481364500918b235017369c94b6bd05f9809b2de4a32da8b357bad93a4a1208c74cc0ff447310ed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bec6498f40909f85366b574610e92644359b8792e543cca0c71337c32afb84a1911407fbcf4173f5efde2db2b62936092aba06afa0297d485c269b5246f584cd69e50c0218498e046ba6afdf69c5f9ddbf370c01006a5b00df08fd02fc45df6ade083b648611213f835db22aa5199b08c1c3b28c1a4a1d77;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bc9d4c52c86a6338ca3395b1bf40b4927d6fd8ee67ff1182bc2f01c78bff1bcab9a8b99832ad5ca62daa973eb711401ccfa15d26337f4e50eaeea83d92dd729271b22652f2d6c9c724037f4920e38cf710470810e86bed7b3e47b07a7308c2e7ab2ddbeda61ef002da5fe508b0accbd9013c47a9de2b7282;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19aeeabf7315fa9f626e4c00179d9ada6f94440215e3f67439f5c6d08c84728fd1ca9de821a3720083b7a325555ea31154a3ec9b46dfcfc9031356d47f03a8b26886ebd6f0599b5f3f17c8de5fe647103c24eeac5485be2a892b2af6d55efaa8e22cf10278197d744e7436040019561924964432dbdf062aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h195825951dd9b35822a789e69011a283eb65adb8b67d0402e40214078f6f3fac8739b525d6ccbdc88efcdf69c2d7b37c5d7f424ec6145a1125f8d33796df4bb7a5c0e4569cd2f48b9138b6f5e35c25244e174f7d54fcfc16268788c5ed22de312cb20d73923561f54591d9ead68430215fc0d4085670ff89b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10d6744e18f0363cbd8991ada4faba9895638f2dd478c61d22eab9c07ed2104a60bad66d326814cfaa168dafcaf09e603219fa3c84b7b144ed10745ff4fcc053a01066e34c284b813c2b6a2a638dbd27837f90f6596451363b2411dbd4d1b3117fd947bdedfb48f9d386f6ff1bcc847c09aca733a70000fc7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9c371f0f50415dd0156cfdb110525485ab04ffbceb32767290cdc9fbd599566b07387e1af4e4ba1c6a970acde8ad2bccaa99adc7310e9902e5441ae39dfddd76f2b7b0656165990ee66bd94aef5a77e3d48474150f83bf9433cf2d35da7ce37399679de873069e1e09d53f7781ee6c65a86ca7c294e14908;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c0e022ebca3b189d2d0dc52247ebc5f303a84b1ed4cac737569ee96d12adfedd6635c456fe4ad18f914e003cc0c0cda305ad8630380088105e40f364cc56bd804612e107a8c51ed05e76ecaf5f5a2cbe9e8ead97908cb30cae71a4f79acd06e09f7444486191b10bfc471f1c8688e30ce6e334ef1b9d7527;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f6e902f05154f1f026f9202dde9d0cba7253ad32ca19de39a1ce4c04708d2bc770f1e093d1e8b06d3eb27d0daa49b23298e3b8cf6df6b01efe18be77448686d6a0b835960b2033a5528bd7c238ad5113dbe7c74e67bb9c2d191a7855ee2a8551112a90c9820b02ce19d7889621c51d895a33e8363045a869;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f11778515881975bf202630e4e3cd2a81e3ce5d04baeeec972fbff367311e8343d2417d69c0508559f87052786c20b3bf26071222552dafe3973c6c7bd6c58e7252089ece194b966433144d55d30c61a0dc6975526f5135a518f813a18362d59a1fc51e893febd3dcee392f4e9fcb7680bb1c81e78ea0e9c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c777c1443986d9600f279e2fcbeb670b1b63a66053ef3565e8b965adf34d6e26c48f6653fad9b7581c5c9e532abd184ff675fc366d2b9abca58efa53c76fc93fd8a40632df7c05b0b763b92cc9b67bf6d2c8f62426b629a96a65587796d2b7a8bd762ddc463bf215666a639fd8fb0667adfee598af096534;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13874283df385b9e4c4189e259031337b36501c5ae3df554d35d14b3bc5c76d1133c26ecb3f33389c4790d3c5d1104086fe28fd0584deabdf28c9c9e331e4bc852b8f24f385d19ad223b9daa1c7b89e4e9e3d8a09ae0a2fbd57af80c6209ec6253c7342103751596dc066e2ec682ea51560b10d58c07922cb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18827bb90e453a7642b4be47d68ea864b9ffca701ea8a727249e51bc79a61ee12f8af3ec0b1719d1fab20116e2d4ffa209af0e03ba50b4fa09333fd56cb185558b2d44c40beb718c6dc3548b0972d9672f899f39fdff0c2fb558a6cd2d76713114bb909f98d544e3093233a6e849936a2da3029aa50f1d67a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13f04109585980beacb317d67bada1066859a89447440d3386e26bac4e5cbc8ea7be2563a5d56d43d2272dc3227276e72f82cdae5d441caa7be0aa3f7d433b96b3918be2913096951ae5d06a2d2f2a800d70a8457997a58c4ef222b0279e3e52778215e45a7caf123ff53ac525de300b832a1eded13c2833a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17511d6bce92a649a4236a8b13a07970c6913123fdba94222021eb099a2182782d3e4c4ea6c3da5e2686f9406a7b0112e068c65cb7ab74d23334a939f63724bdf75237df7ca9e8036d43da157211c47ef585dc3ea02c7830bfe19d1203aa76e357e8d94fc61b93a2860f7eddc54811f4606869feb5c08eb22;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d2ae1ad7c772cd9ab8ee7bbe4f80c71fc61e30d2bab279ebb9f64c0837487825702bb4e14ced83373313edcc426b957a8c15b8d77aecd47c07e9e63eae593b45d9ed7d21bce7ced64c91067aaef099e303f7d8a181cecaf64d69f6b48ed07787db598c23b56e364306268aad3065a5782dc8eef8d28340b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h88a5d585288782da1f1c0eff80cfee700201e8f9f20a84207db434ebef5558d04d2032797570f167b84aecc80738cc3423ae06e4109690ad0ab03b8c7c968d4021173418e8b3529b77b19667c427cb674aa78c633c08d51b0d0792e75f01e557255ff6e975a4a78e1dc04619c9b9acde95454113666f5cfe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h86370baa7056529c0b911d5c8af75585decfd4c383febcebdbe1467c9b90c60927c24e60629b2aa6b49e476348adfa1b867d673512d9dffb8c891ced049e0128b35b24644431e773cb99e86d07c56554ccd61374d585533e5e2ad42ea776329900c4c8e3490c63980acced4885f1f24daafd1402d6ce93aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h52f3c4dcc2c874edc727a958a9fb69bc368757ee0856eeeca698424978f842f3b88d5523b549d2ff88be1a5051e4a9fcb4412ec6068d87a7ac7f9b742dcb3cbe052b867957eba0a8d1f3dfa7bbfa65f4d90c90d77f2690d1f105049074c9f163db2587a0757d17e1ae600335442bafffd1752a8e82a2708c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b451b1f35ee2a1a6f6a615906e5ac35e8d98177fbb87c704492c48f712c82ac78f687d87466c2bcc2524048741aaf110224617ef88077c8c7ab6674cf4e1989a04e4b6859ca725773efd9fff786187ad7641a428a8ae3c8576b69b64afa72fba5b198fe5364daf35b3489b5da51c38d4f40be5dc8c51789d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5d181eb9479bc2df424786a04d1b0188f9f6962e03793d8f04428ea4aa24b95cca2e3261d533775491ce778f2592dbcadf0cc977849fc83eb1ff9a5472d12b1d5f9533214917f0ca32ef1227977d5d8aafc10e8e72070cab9a8cdd0d9a258ec2e5a8386f5c5c28d4e684c860f1a23ca2b86db8c69a016070;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15577cc51abef6ed1b487ecadd2f8f21f8285cc513b588728ba8b5f49074b85874b55cb683fc39abc3017341147a4617a3bfc06e1ba8d71cd9a4fdc0049496781c150a475dbc33fc67cefa8bd0dbb76bd72faeaaf8c3112f33b925e23189246b4098711e04129f8428c40f8ee1d19666f0bf1463e8702ac1b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4d6d32798f00ef34d6574dbafe2fc103ef55ecc136afc201a83bdd185372a53ffaebe6ba93461c10c7b5e186433c7d2da393344ed46632034d6e1281635b2ea54a0292897fff3805418afcb5fa5f625c633f5e067808a64f8af6e65ae12502659bc0cbd42d74694fb0cf8b202d84e0a1602c7bfa7e9124b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb18a81bf14225e7e67168865eda226de789634c2ec5dcd162511c17d4defb223cd80d2e151b5f286beb6b8c866bd72ff7f661b84ff4723243fcd29b60bfa13ae33f54b2b60aa056a14a15d7108f7a9613d8d8062eb9e64f8baffe9eda139085e7e3c2ef80f9a0770e864694656f5ba05be48d5ab7494de16;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h49b3db94ce0311ff1949df79ac1c1a24c5f44342c0544807a5b209d8e60de6ebc4dd80e633976a4f69ed775d62f76122352f9c2cdceebdd867f36457b10048021d42cf24e4f35c94cc337ed0706b51b273e2ad9bda0e9e964b1cf9b24834dab00867fc8cb937784be57416c587701c39e73e25f952d9201a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f23243b6ee357502903aef7ec33d6584e6d9f0bd0dc455c1a592a02385ea347dc8d9ad2d8bcdb978e43e2d92f53c6457fa092b72b4495d9b84adc9e3892800b876bbf30270683c238dad5cf217883cd875bce617b196883788943341cb129eeece5a7211669345cac21d450b10b0eaf3544b4e37b32998c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h43c2afd251d367946038d295f63915f46bdf75f5e4d85d4f496d6f5e5dea86bef42d371ce5644aa62471fc6bc3377e120cc9a04b430eb8b0dc48eccacfddbbefd5e84c04f7bd5c0e3af32e31587f19cb6cc458417da8b9906a35bff3e779897b3ba7ab871a7da30eff9bc7a9c1176108c5bec71389f1f788;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h180298b003d049d3f60445db4671952a8aecb2376f98b2824a583bd3c0bc8a76d0cdfb7b64c81a744dc98e16fa3de655848fbc8d5a894f9155875782361557c714956afcb14cf90d26404347a6ab1a4043188d651ae98117d8e05dc612451b7f0788ce59863b948417ba431d0c7d57e0bcd6369359595b81e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17c9d50d4d4bb34402677d3f0ef3f286e2d221fd55045379b608f495756b8816d08cc62be6735dfb0e832c2c052b6a7d6b51532beacf09e11878dccc0e6365747c330710f748b00a7212647d967daf0c1817604bb11312c3152d823ed5126aed4897eba31e4cf81ca1f8686ac8faf9a2267e7e3d84c6321ed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17a3ab9bb42d65ec070223b710ad831292ee3f16989b978ad34efd04e6f039a43116a2f27ce4a947e92c0852b8789a874aa2e04e49505e924aaeafe812a9ccd964bde5d55ea5ab4f9207f07f004531b48445a1efc7a86a2e4cd5d6cbe0052c429a5110f146120f1de519c4d675ff940752fc5684aa94cbc86;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h260dca7e47077eb286761e999be3f9c11aa89391b876c06649008948d801345c71120f567527ab6d100c51dac65c4886bd2067ffa9e303278f176619ad5bade40347bbc3c5fb5ee82d8c8824f34b393687aa68a0f440e60c543fc88ed6e610d6adbdbb2bd490d0db7e6460290df44ff0ccdffb3a329d0508;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ca1a2bc984f61df795762d55d3b50a425a83efab7a43eeda2c6c73079f0304f7118d441de515818eec40f9b8f268303fdbd73e4cbd1544e51b13c44fc7fa0b32a31847b4c5909e6e0cb1e44c2d9aebe205c5286d7d6230ca36c6a2db7a3e67de55c8f3f868409de54af2f08b236abe062f35712e108e2214;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e59aa1bf97adde94c4f4ade55a2f416bf457fa674ca5768d6ce5c74bc7f704e2d36c81c8bffe7271d725e6753fa75ac684ea8299a71def4953fd4116be2af51c48bdb643dd2d7c70fc7549f4aff4ea5e493153bd19fd60375c5efda8111e449c497984abbf61f5a76cfbceeda633b38b5987b027eeeb1b64;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hba7283c750819485e131e89617320a80bbd92f4476aa85ca6b61ce539f1edcbed75eccd2e425ab7e011e8d3c0534deabe73f5d9bab8e094fe849e19bac6aa444b841ca6e749ab520f3ae2766069b24a3a5f5dd3727763bfe7d62aea3100f2a583b5091268c99d8a5d565f2ce98d4dc9108fe0e9fde7c0909;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h70f2a9afa7a7c85f0210d0840dd900e5944df5691078cdc2bd39a5f001e8807c1026fa01b003beff601ae9c780f1faa24e4ae44ad7381133baa29e2c2c9b23b891592e8338eabfbab037879b61023cd37dd7fa0c8d815d6b4502659ffdd4b0b6e05fa17f9e05489db105fbd7ca3823e6581589a1092a00c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14ce95886f06f806412346c9f9e3e81985f9dca28166fd53478176ce7df8775254889127f59da64c70e52e95532664fee60ff5e439feaf89df3e4077c46b1df9b695212db1be420c7c8fb310d1d20a24c6452bc8180dedc58a476a6aee7edb1b6e923e0914d82ebe3ae613da8e5b8ea968037269ed2e9456e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1120bb465ab90a6317fe4671aa5bb27bc7f391bc2f4fad728a23767541150a8d485aa6362cad2c4793c3dddc4d502f16a9db04432b789bb52ee392692e93f785c5f2742b41ac73b767b87b268a0ff6a816f02d0646eceb2ce2d59c51e0d0957256b464aeb731661db8ff20ba624354b0e8f20cc85a7620a3f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11f2380ea5946fbce4464a6b4a9b46893922b96a64e4c64fc5209048b166b24fe50001d1ef4a52ad55b57fc28cc2515449fb83de68e248ef6f726c1603efe511f80fff6a0b64a86e14b07d24eb8ae12e0fc5f8e0c5d26701e7fc47637fd80915f1e1680ff31b2e8cee79bb226afaf9bb2f98f7c7fe3e918d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcb58f1c62cf4906037f65e43283484ecbfbd17bf3d3ca12d577b1e2df97566066bb7e7b69680cab4c477b8539052b4671e14c388b24a48554a0669e3ef90dbe83468a44da356b602ba99642eb4030e81d4c9a85b73dbdc7d2acaf50cbd128ab17aa3b410edf7808c6c925c71dc050720c988890782c6c2ea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d75d8e8f74399d12dbcf29268e553a7bc07f05b584f5b493d4e991c533ca7251b93c57a5e58a09d0874ec214fab0008ec7d9b0c7ae2a4d9f0362bcee44a2e71e6b0e6a2299709bfb09d1f8e846a850d6489f8398059748df4bbcbef265857c78590af1dc1134815aa11ebe0e8a6d95c82cfd69089c8f27b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h34b057205331307c15c36f4187692e40fc6de9ea613e33b2a08f1adb6906309d23a230a7297f3285243405f77e79696724d3dddd8fbf5cd90b1888e735ebecbc799d0082b8e6d42b0c65f31dd4e45b27a4824b100a58fe012d17ecb4be10dd8f06fa0388fbbd6064c1e715b9c61d45d5bc2e0356a66261f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16bce016410fa809c291d95812799fc80b22a916741dd3ae47187518b7c25223bbb27efa3aec6516a376a6ab0ba2f2c7f97bd05e566fb6faf71af2acdaaa83c04e100c1d8a6de2073eb68ac9e5f7949d35fa71b5f6f46965a584ecbf287532387432b4f7fe9dc26304c3c299287dd592e92aa85420034b196;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f4b2042222176cf5859ae6989d576f731c56c7f96c2ff783fac83bd0c2e70585808087bd0abbfc45b39d855eda1f0c1ef7a7526d812dedd8630e26ca7c452cf819cfb2a1be80d12da2dcd7f24cb130141cb8f03395e4aac7ef9748f230e9e72ee6d08e49355f8e6147e504e802a67dea0925b27e6d7d5b78;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd34260bd8811e4edd3a9703ee6df746152c9c9519c34d5bc84998932d31356f74a6e0d0a302288905beed17c1272d4366c14b11bd7b84d9b6597cb3d645cc6d103b0b2191a0d2a38f6b3a11def8f77b3eb80922b8f8187872b0fbb22450a23be6392ff730311333029131935931ec30e8bc062ef5e27bb8f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f67e0c417b0d11bdd39277d62d9cf23b673e9563a20ec5f547baaf2ed4784f00f31d9a408b03f7eee3df65bcf60356ea5db4f02f9b2a7ecf8fc60fc25045555922fd97f88929c6581b776de2c0dac59f611b8832c6f3075dba82fce4142ddbab2b9187fdce4f6e5fc64395f0e9de84bf013361f0ce2f40e7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18a1f9f38437d4422b256b13c077bb6aa4657dba02cde69d80b938d73b785a972056eda2623f3df0d8eec649fd61fe118a36228be4b5d028db270bb451339566c9d2d4591b311108324eac2c953b0bfeb76c1fa2d7d9a2ff33f13536b3f67fd245eea6a683539b82f758513c64e17f099fa91b1d95af16843;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c5c5ba62c30b48b890005a8b1e1fdde5b1d5778cb22d0398b38b917bd505c403fa4990c45cc465eeed8b6b03888d307152bfea017457e0430c05dc468813fa5f02459022e8d5be0f721661978d4a47936811db03854fde020af1c1861f42b195fdb1e53b7c8118aab973910621b02c853e4a8a3463994d3b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c936a034adcc7d336732bddc687f65a682bad91213c85b8110c106769a5a6b55346ab8d60e773f2027c2ac904c86bd8092243953d6ea0b2a9d9695abbb238722fe2c4a4bfbc170cb85d324dc09fda9d372687669e968963dc53fd5aed3df33314315d3a5d93a16d43ec0b8da8d8de934adbdae11b62a0e7f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a914601addbf086f1ca4f355977dba5d7f440bb1ae7326defc868541e408dec3c59b95a87e44f4510439159d31f0e8380537b7ed630d891a542677dada0afcd07158b9d46245a33ae3d5aeb20d32a1bad972ca3ef5557e2efe15d2199a46aa2a0733f6d265b3e585ec7a23c03231b82c83e02194c8a9d268;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3e30400bc61729a9757be629fd00518163bfed86b8610e6a93dd1dc168b6793d404f0225c20e68d09208c632cf4822c2fb6f00ff950f94b0438ec39caf5bf83ea1843e6f48ce02d59a58466994f8a407f120aab1030611394cf9f873f5e31369def8dc68ae1e185be05fca9416c952cdbaf83c0f5b5e55e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h57411a1efe1e7c5fff799f09e9f9760f89199105131ba44c50c4c9802cf0322b66b2c2c3327d40dd191f207d779ac2d6f22eeb1e8fa2c3cbeacd9d89cb130d5fc15e234b048c0a96c675a49f48f6bc0c59d8d4542cc50afa086e697e19b02d5151af74916b10be581ca405514a95683ff3b3b40ecd065a67;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfe9facc3553b999e6b839acdec867584fea2ad0868299e07d3f23c9874ad69ed1144738cb893a2f5f7ff705e69d6db42ad034ec20bad4656d3908e0daeae277a5fed921e4350e79b37c6f304c53dbd027068bc22aae27879413012fad14ba8392a457e5a6e5d63002b8718c44e5a0849f5a7aec9a1254d05;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5277335d3d65803d1991b49f795785ecf950f27b3f19ba8d8bf658ecf2113ed3d5e055e0bac9c089b2062799f604ff0ab752afe2d351ec470d2931acb848d8871ed4f1c9f90f84bccec934e6ec324132473c7d2b53a169640b9dd74d1b0a3ff943a52747bd1ec69a962534c6c556c97cd039d7dd45d99788;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h556f9ef267309f8acbbb333f7419725d0faca606b05e0502bc4e0ef318d340544e43cad75f866f12078fb48190d01abbe8fb45a6168bc0767a63d52d20ca770557f0ca188173914122817f54b99f4e43933578f52911dd4b2bb40e3d81b955116c49779f6343c3149c71a4c894a3722c94073a841c53b994;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12e93aed600c38d4436d07c384d88e55dc0e4d6b4fbdcbc57cd468bcef9ac91dc8f2c68f117c5b44b64d8bc38899a437a46307bfda4c0e99d1897279c9ff5d6a11182a674290861ebbb186dbdbc41f4b05d5ff7364c34a34a95ab37eb71205376a2114fddcb9dffa6c41ecd82b7f1244dbf908be3206ace3a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc8b8118a37b10963608f7b5571c8199b1ccd5cfbc92749bee6662968cec3ba263981feab90ac8925eeecf2ade822da691d23b542d42885ec22364d1bfba9930ea9af358d34f6729d44a56b7d17b393ec09cc9c3ef6b8385559d93e1997de2bc2a2673450295a417e5622b46321ba9a23d84893a445bb8717;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h189e495f8ff0f1998f8f83567c95c4b34508e7eea2e7c871f8e9c8b09cbc3318476fccb3db5c0ad3a104c2147c62cd68fc5d9847b0531b6fc8d19fc66b12033630f6af6cb01feb2df4f08728aaa677e4f101033788f39155451ecbeb8ab627df75618993fbc05d696a1e208ec32ef79aee2381c6c4e4d28d9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h99736a6be3c23fea6944162d73241a2376b5435a6f0688b04568f9b383682d33a36f8f6928b45752a95138270512515a621fb0cd7e53cb6d762cd18fdea6e7d80d53a330f98d3a10851f6e0e63540386bcf92cd352ccf4bd78d5e3b924b0c2121d845edec5a1775aa52a38478f56c519e8a09669cf56fd81;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h100f5b647bac32a38d2ee05fd6c9d7bd20d8440462818c432161f9ecc06b0bce75f169387f132e632edb465221a428521617e2a6d40d29891389ad8d6ebf6e433ef0c80c341814c3a5a7fe99b7b3db0ecc7314fdaad6af4981bbd4f4c6407f512b24f707099f0672f4352c95197280894f1cf2bc3857cafb4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fd274370a5e9b261f445e3a9740a8c32873ac2297fa36b531d2fed739bf1f76078deca1c690f5265bd5d74bfea086ed3b671b6f949f13225f8927445e80ccede3d18e045a18b385b8cf0c830f3c18c880fbc9a493f09792472cae5455ca8d30fee8aeccc6e7fd70668eb8db630aee49bdbaa3b32fdfc0740;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18a1e37cd15babd4d229d3766cfda6033e8ba7a03f7f1ef5004dce81ca662a1f139b78d2a77369a34702ac7e65c037e5dc1e8fa1a82d73442c37ace618fc6d7960239dbedd7a3ab1a3ffb964c57b234f09af5bc5052e59731d3568d277635ea9e44ef3d87d780ef184d95464abe3e6c2eed3195a3b84d7b16;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f07271cd913fb0b0914a28428b19325470834d1417fd0c063ea9b0219c0d43063ad3e3f6555b33955e34d2e5d50d1b5a83535af983e8d23ffdcb4ccd06df328249fbe1b1650fab6922bb495f90989f5d1c596b11a946499fa90082e24bac83ecc352ad250e90ced6c51a532cb4f640be4424defef69615a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc8fd066c843208e35e92f2053fe784769e54d2495d58689bb4d13a78998c6678289c4d33dae76774e32d20b8f2f7ce1f5afccfb8eb90b96d114fa757cc5ba13a7462ecd5a728f27196018430b45bdd8c4a1bcabd68c5bb357f3d66cd043fbf3766504c59d30a64deaecb343809f08bf58bec84fea011a819;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14ac02460de4f996d260e4163f9deafe4614275186cd509c5ff563de2b1339b32b727c67ed3d24fa59a0c7bcebccd8f9b7a59539839d9349f25615f0e6901a136f9ee6a63fd94fe603764d83e0ce986ae48df75254120ece6da3793dfbc42d327b766babb9175268d181fdc3c3ec71ab338f8abb520ca70d3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h184e4b28da69c817d3cb5422d745653fbe542c20dd3116255aec77489ee69f2751f5ba84602355aeb3c1a42785d43af80226e91d3015c2e90bf08a58da501bace6ac78d53d99755ecb97f613f69eea8d6a716091677a6630d750867f1db89522cbcaa004b92398d855adc5e030cb3f9adb2410bc3c6488ed3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc61c9575aade843c0d4aacc035a29d94eb5f8f96f8390696c435ce0c6554e97ac558644b8d628d04f894215126425d2cb70cd7793fd44145111a615a67195a689f83a7f8826281d4637c26bd05de0043a03565c42d9ad4b6fb9b8ac5e38f5d9ded8887d7215854e13a44af8f853cb3e03e8d0645f36d887a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdbff8c05108960fb618adeed5b6c0f20df71f6f166cd012b4ba02442409ccdc8cfe394686d37ef0f095e0b39ac63f40524f82114bda0906770049ce5ac38e886e165f58fe86d51fb4c641a1d7a2d80bc28d16c9c0935f0cf8c7d1a98255c1e7225d9ebc306e25a160a6d9547024b8b631ba24423fbd077e4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he44778715445866435caeb3d40d6d5c99e637b481a7aab3cb36ef3e44a876b70fa328ca684fe11cbe3bd1534f9baaf3f554e0f77daac3f435a67f9e8c81c7ece25675cf31d0499e977569c35a054347523f00c9405c11333c86ac8f8df70b5cc20ee0ea1f60c6f1a73cd7bdea540ed5a56b5bb10b9eae923;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd7ff38094b27e5e7d0ddaa80921eb7dd48f11f1692bfa5f27fa6aae5337e678299fbe45be2b1c7201b3dc40baef6c44fba66783080ba204a4a178125e8a155001e3e812633c6a2533cd81a47336264f3000343fe2e8f72ce30eeb23d5fce16246af328ae4286b420d5372ae92455c99ad386e7c3806a9483;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h28d6bf09f0a77b4d0cb5b1052ec60fae40643773d6cf3ee822dd9ac8df6300f7d8878e2339caabdce42bb3ec728f0819c19b343367f21531db1b82bebd37a9c2f86f7a048badab3867204b9a27435c74aba66560e195f536cf88538f5d8263ae8fff07fc6df57c8f0ff6c944714d50fd218147d315fedeeb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h195359811c9d77b8a5cd0ac6af65b90cb0b65e3194ad674a8d54a6ea816d3d4e929dd4616a894e83e6db4b50a3a1e316a8b97762d3e7a4db49b8741c0f13db738ae746d05f281e712cdda066bf62f003c3d7935dd267ca3acab489c35620a0b3acf12d2034daf5b338bf944c605bef8882af52004230e8b14;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dbdcf5a0e16b89de5f0ae286d883863917917bdc97e0cb818a30300e9a68ad3cfb83522663559bcbd0436cf7eaac6fd6521250340f5867289773daadd494dd083a517fa1ea78692a726eba79ef7513d90021b4cb9336969cedef22ba25c9352d61e622f902b798eff2182f0bb3e8e1c5c0bdc918bb35ecbb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4a23e968a13ab06af05272c0d18e44d1128b030079ee45b3fda1c5902bddfced67ed36470e75d9173533f1384a0126efb4fe6a2a4677d36962e20ec8a2b2fe307d9fd48a02f9536a90523e908fb307e45359e321e3b70684ace7320243dbf0b7f77f5c0aa4cfbd5d8b0613dc338c890e215946c6f10f5b7f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbbb95d6a10889d0fa5c931c7c4b92b1a6b8efeec3bae53e2066086d2e1b46c7617afb9f85a644bd3d6c04c2af99099147137f225af8e4259ea465e9979663989db39d13b5977d0fc073b7b0fd026f8a4e2efee42c1a57d6ff35e36091e89377effd56565c1209e6e4673e43798b08d55e90bfb3f2bc59995;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he1057e8255d9f56aa0f910311f44085aa8026824cdfa3adc7363b69eca0e2cd81c63c3b880e8901bc4cb7348e3160463bbfd85a6ecf9c60627aecfad0f05ced110dec75e55be153de05aaffffd31a29d7bd730b2f2358cb54dbe5235fe37beb6bc3b0f83d52da2492a15c423f49d417fad9bf62111fd1d4a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1819f73c162b46ab3fccd8e1ec9841277246f3b5cb4ecc6e60e9fdb193fa8d9df355ea751bc349daef568f7e745e7b7c8a6f81ca1dd76b8d6fa8bce2a35818ce82d9f6614c6615f7649520a309b097b7f55d571b08f3be8404ca1516e0d3c5c25802aac18455adb301168a1376361a3d68054e5a1139e5ebc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1076b0d42cdd2d56d511737005f3f321b43bf309fb00657342e49c9123c868e02c27fd1ddeaaf4f7c8b5b6816d929dfe0af200013705fb604a9bba05cc5072ff6e58c05629c376099272a5a5d9ddadf74df7ac515ad33b06e7d24f019e38a9e1cce53699959525e88d57d539aa0984add48d04f7d6ce30cb9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13747bf02d71f92d6c956838825d2bbd14df56383ed35bb2501994ecc060c45f75471c779d2be0135b6de77f723f0e79fdc997d8d4c13dc7363c8e613a97efca15dbc4adc8f9abe54abc9f77d279bc937a0b8bbcdf6e8cd1456d74990784b46be430d50443e48e010083c8ae66dd50d091424d0ac84f87768;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16a931e457c6f6d112e7e1d913c8372275784a59766d33d645ed308a60e0f4f6cca51b5019fe6e2c4e60416d7906ea8c68953a92b071ca4da47be4e66736b7abbc6a55062f4acbbbf749e90e2db34a86eda370c4fff0b7f085b6344f7f411e3cab9c3c86420eb822c69ed3f25276decda0bdf6d2405128542;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h139f7c805043c9d2c32f161246be489dd92d65dcfbe2b1aa944e256dd45c3be468022b46786b14f8df954bee564863eb1ac7a90ba01a4f929e774bf9c8a2f45f20e1c95b57f8ed6b872779290ed47c7f7ac899c123e494a9d07d1208df2b663f1f0fbf9525a1a308b23a13fdc48a0045111f6475dba69108f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5e27ef0d82f33effd8fe3fbd9b62f500a8e73c7f77b505bad03de620f564c56df2c90e3a2812daffd12aa565ad8c0df23107fc84ba6570d96294587058d64f5c43010fc8d6d4be2c6f1b6774dad1fded95cc3bff22e6aea40959f5ca6c06d6fbec1b2c06879dbfa5b04ad154bdbc5da6ca23fb21ca114b22;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1099699f90f2fdad5316dba0df615cc5e63516e5ce719ce6ce01c36f53bb51799ace445790c21cf41fb2b3096c3df7c129e00481282bfc4af3b0622201bb8f6341d9b321888208940bdaeddad5685d3a1facfdfd0ca37a9eb7697fc7a2995f014feebea0254e5ad1f32e4412248ea8eccdb848345565082c5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h103db2c1193424b53f777613860cf5370850c424c8f05be06e10df574ff3bcc8f7bf2508c16678a6500ca6f0dba34d0ba8436c553395d51b79903e79ea338b882f55bb3ed7a03957d63fb61cbe982fbcc7e686dde5f31df34e323061f48bc6b2c890702ba8603521be8610c5c9dc4ad32047e8ff908c5a74a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h940e467f30d00ee5d58aa513d738ac08a8ad2553f049ec9fba863d7d012c10600a6b1edbc43c60ba5ac4d19bce7cf3fa4fc58f33d064849e10599772b4ccd6c7054f0f7436c48fd3733b2e883a9ba66daef904222a45e6798d4958b06653471c3d87ac70cbb513c0663cc1e41ba5c91c84b014bb1b8bda05;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h142cb179f173f9373b3b943cb1f4c1302da40bcacbd8eb631684535aad5447df551bdb73084880873903c966fe4d9492f76e9d5d0c7ce95caef9cb43be530193bb191c8634d100a0001fd52ff8d0917e9a68058961a074bff365041025b82a4cf773cccdab69de6cc0270d9ecca6b404ea20c24edc1eb62b5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h60cd05b829d6c0d7eff76785a12d18a14e75928f1a75a3955961355d023edca52b9bb992ee45a931d5a3c8dda88bb90fb1d3a75fa38e759f136f8f5591d92e0135f463562d4a1c17f0bd263960cd0153c5fbb9a8989306489abbd0ac99a98d8aa5c36769224c50a9d75c84ac626cb30475a3954505f4ae82;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1541666df4f22ea89f626bbec9328d916d3caa738bd65f9348f4c275de53e029f6dfd66c3cf850106a8430056c351e6ead3f2e2b6a1238d60259d3b09761528b161dcbb402476ad13637dafd895543cc542d95a04b9087fd4a285eba42f9033cfacc024957514e391add67fa319c2e8a1cf98b9b0ab236e7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h71be714cc87607bfc3345ecf596179685ff7f2dfdc8a4496decfdc6a62ca9694844520bf0bc05b6db7acbe5a62f5ef0ecb6df53ddca06522a6e04bae8cce2ab3c1377be5b58af2576cf652ff2d93d97cfc359c757867268dc1a314e5cb4d6f8978a9a935fb7162079d9cc0bde358c865c473eaaa14ea9f2c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h64eadb7a7a3607e7f9085912ce6212f6204d0dd784d9a6aa1d4fecaca664c2d37c6a0bd0b6c6a9abf863a2d94bad228767bc071be8d6ddbbe500c8676d5aa8a8b2d29e9237d95bf96804f1494edf974dc37a1812483052a13131aab3b9bea0f346ea6f1db158eaa1c6182d71c63cf8522ec6f3d1815532fc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15deb4c5d54c630589ea8c60c957e8a652d9cc563b9e52edf1364b1cc8c22a0435f230c6913dda663f2f2aa3376f1237040f5e6b6fa0140a107c304b3496c2d37a1aa1d5c6b79bd2426d2c6094f9a7b100b4e0279ae34b0dadfcf28c2c5f30f09b210badc60397f87496988bab2118e10173967ed5c8bae8b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4abe38232a6d8af6ae69649468fbb337f3fbb371230644aaca26930d127ae1c8f542b8fb59b3105a0836801f9243f1af129511b33a9ad6b9c5dd407a75b44213f70a8010f026e38fff676b00945b4ebfdbf0c8c0deb40aac41622f2ddbc7d7fc2e9571caae260fd83c0a4c0e473a569cf5e65efdc1c4f892;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h400441a1c80cfaff593f86a8de8b377d6f77aab547905703f98b2633e257f5dcd8900a6cfc8ddc35218010ce8ad7aa28558b99d9150c579023cb3bedc72fc33abd315ad513f63e8f1294e36fa0caa9df06fc7b645f2ad0f5ebee5abb7c6f94cf8356150a19854936eea3103c22cb735e9a2b730de020e7de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c69fc046a601d3e6898e6267615702c0d16fa24a16c0d2f6afde0b1416cec850da5bf60463f4590a0e6dbbcac8dda649aac58ecd7129bfad448d1be67f35e487054425f788d61fed44996565b700350113d2a8201dd5cfa918ddbd7fd32b71cf62c11ba29d0e9de5a5276e590e7c2855dc102e7d8873b7c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h35e894f1a651ad8c5bac2eb159b25beb44c7d8402e42350e7d56aa14f55419de3e1c8b6e08dec747db297bfec269ca94c0e9eba79b113d8baaca7e0e4e2aa5bed01796ee3b8e50833405588644167a092256daaa22b921674c6383f4cff666bd62a3292597b0e6ac41edd2fac92219358d8f3376a12e9308;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h186cdfae37f47891b37878af3b6d0245464a20dd7c9cda1d2fb53ae8ab34a879bdc0740dbaeb194dcaabcf8555459e91370dfd93623085954165e3b14dfd8fcbb7868c956fe2eb7ff1412ecb15178d79df9a75be7003ef8e44be04cd12d1d1214136398a39c279462623f6088517e786ca2daa30a5a7082;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5772174236c749796454669520acbf1a25e95ae99ab07e2e48c932bd59df9ee3f2e6b3871b1a31136c8b2d4f389bc5a39d11f21d5474f700050d276dafbe167d31a25c5e56742ccd62ea8092f7d0cdd3a62fd2744e9a87a470174a571556481cd62b468e877ac4847708c06763c137eaeb74efe565a22871;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb6cd3a1f2e43b4ce340170cb4b53bf3aa256468e2712eeea8860f7cb614dfd7bdccb9b2d1ab06055555387369376e7fff73bc0efaa3a860d8ab6cef65c3be8908bd9fbf391c88831cb83da7d0387bc4adc0610a20d6eac435e3f38651b50f87ce92493295316b984d0575ed6be59b4a1840f76355823b2cc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc7177f09eaeaeedbe030ed9b1c60f89f241f9e76be51baf765198d517465e9213974b402534a877bf3806cce972d33d3e66cadd949915b55b4026020c3812d3cfcfaa78b05d536dc7a04581e3cdd9d3cbe612bf8eb6e526693f19fb0e5886fb76058db2cb99dfa9978e0cd2c6d15334c66b03fc3c4e3e97;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3eca9a7341b1a549e1b89d98f23d2a283aa938a21606662c710e2f563dffdc10493f63f297e360148f6cf73bf6778e9295a0f4d847056d0810ce807bb80f67cb4bb36de18ed1f2c8de4b4c6dd7c2eeea92c951dddcfcdc663e35cf27bc9b90558bbeb413beb814f47ad5c57192a0ea3bcb3ae890384ba1d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19ac76de586e5855ae5217bcbc5c6c29cfc0187fd2cde158e700ef732a5859acc9628fce99534e9093f515ff78665d21e9f6bacc9a7f4cef94b3d0d6ce05d1ef1f1c4370dcddd846c1ef027e939260c25a58362e8e423a6004f3b97e5e58b9e13470b0281b5f2ad15e4f1105dd6ecc61ba80c5ad4e67ee6dd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h182e79bdbaacd32e0facc363f883df8556f5d1d6d549b0e2f32f64257d3d4100c17de889df5383210482b358e4054ce7bf8f1301e4c45728899e987dbd2e5f2e1b79ca360f68374b8f1f3ff556246a4f5c17864fb767e178f405f9456316dd1117d8d1fd97b0c77cd0229877d3dedd8d4c443929fe7b29dd6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13eaeefc889ffaa08be004eff1c281cfb15e833552517de12b992b5c1d6a024d80c31c1f4f64ffc830172743c2925812b848a714a3534eb8e56f5a9881707dce9f1982f25a1d46afc38003f5c6dc3a7b4ce32e54ce1be85fe2ba24cdbdc3f2d215a447d82c727dc9f1647544b75389db72de6387eca3788f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hebeb273e6815cb2a3a03128f6706664d360f65f5ea609bf269d7d4c4253a919653c28c8a2da80fd8d59ceff4e7e8734a5a401eb0eb36b0a4d55decb5a815afc0e3463ce6d2bde6c64cdef9adba72bec0f2a397a857ca23335ed4c0b05fcd84466e9142caa0412d4d9c26f6e4de903355fbbd1066b183f6a4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e0c84481e44e478fc8a5d264b143ceac28c24d5331c72c61a4d491e248b4f3445d4b6074d3d95e802190d91f5a399bb2fa17e34ee020846182e7ec5d26fcdb26f57e5199fec0ee83d51c93fc455cbfdaf2c6c33b07e31a0132336ca762b7f35ad60632bd1e97c4911539494eccffd0ea7b981ed090153b0b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15a01d5bd9b90e0f2e3c3479f3c53a307b16cd58fe5000f3c5f07773d1507242b192d504b5b1586d88a833159000a6a36f70fd98ecb262a38e5631e355f61c94e09cc05cea95e6fd73428388adedc3d175fa9c272adb3dc2b7d7ab146e3bc1888a178f3ead1399d81e9d125e3d505f973e0fc9793c83a110;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1845356e599dc9f45208a5fb9a73c320a5dd29ce806adb2dc7da8656a48980489d2e743bc800dc4ca60d757002c4252da150651e0a908b9048f909078444ccd80b807a211188271a96a9de1e54661586bb40ce6d70a87f6f1591dd0c85208fdf1ccd4800647757c7131ac97007330258f86a75536f932d400;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bb082ddcd4a766651ec23391fe64c422f91121994b721aff12e8f579c32f3a73738aa0a2d126b0f0d144ebcb830d267310a1592cbd8dee41ba3f4b7ab0da8e6a78cea65bb09d9ce2d907dac6b76435f2a19a98cbe46a0d0158f8562b95c9233d67bb0effa865d42f259d0921e3cbfc5fdf7fdf46ecb3ddfc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd9176771def5ecfde1e92e42d7dbaa227ad4f97e8a849dc7b07de1c900e368c2fd70345229f187a85b18e0eee239175cb01ef655d418580ad03a7914e32e13b6bf198386779207bf28d558f4a253d26a1b9195e6136889acc16bd20c136c5e69671d983d3ddd8d73dc0cf388feb448f5356e96605bfbb84d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hed72f09879ef756640ff0fbc3ed54d280ecce497b5cff9d5180bfbd3a63ca97feaf28986dbb44f2a2fcea386455dc31499bb913cfc037a5b72995bd8fe701f9e7e49bed2603eaf653261b7c6c6b001701595bdbff532028cc51ce36a79ee5a7bc9e38ce2eb67fc47899b2b0a874406a59faf862537119374;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h194967131723f5d67402b97130a5dccf02441a24fe5971f4b6251935a19263adf4eb19b55630b17de5ae57de3b70b91acfdb6881017be7ad0325be04f0e548e92ced96f54a93ba148de76633f443da649f4b353a606546defdba6fe4340af098b2f7143e98352647df2374bcc54d76a5e680d948331b0861f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he0c1141970f8b9acb85c5da53287ff1ff2ec4fe0416f5d4421e43d0e97c16789dbbd73733a0f8f3e4bb21c49c5aea4ffb227c39793de36acfd95932aa9f3813e125fd219aa108bd1a91e843005f9e3c1855048cdd189f36ac36d3dc3ad7f0a37cd0afba86174e6b6490343b54fc3562b921e5a83627762ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11590e95cc4bf2ba4df0d45d42052fcdaf667d29c7ad9d34bdf1b6ed428b76931f46d007a1c7bd6fb347781ed106e06a3b4d21f3fbf2a0a911ed9a15ed377a58e3051d36ddea6ed99e4936a381a54be09f8dc81c860589f324946f4f9c70953e7c72277b1d79200d03cb92b6c46187e0f532701343ed9fa76;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h66dff8181ea76b1415fbff7effff4b7d966eee08dff5181ca69e8b749116e72d1b6b4298f0e32edbf02456fd6130c1e2e5c615599ba3977ad420c36aec34c0754feae65409e6e9fb45b67e974b1ab6d6eb7b64053c08246c52a6ff3830612ea703e228bdcfaa9603a241bc5e256b352ecf11995b327b3dfc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16343fdb9c90538789eeb968463d352878d78e929dc52b5691aa2091a2a1f3c759711a4aca1da315abb3df9af607baccba9e74b401a78871be19aa25c91fefdeb5a9bfe786829cf458395c89e3bddbc0914a5992572bd0c33a1f5ab5bf75bc94e8123ec5c46dd311de6fe1cf9a39d16ccfa2c36598cddc75;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h770acac1bebed892e1a6bcb339f4ad62239338214c306277f6c52b65ee243d40d1a185895a344b01be2ad8dfaa7519abdbeb00388cebc97fcc3d38a07d2dce34bf85c5c0daf5b3d9aaab16019980972132bd197d590d801f9f6f8fa2b21faac19bc5c8683ded0c77ec11e3b3c5e9c1a8572dbc167d2ac220;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbde48a19f7a01fe463ba38568bd6194b509b7c1590c2831a163be43485f3fb7609138304378a446b90126fe90e4bea7693ebc7efb52829d64e949276ebb118221cf95a315caa12c3744c492cdf0854737322b2e2d945bda71b5e965fef9a4a861f7e87a48898f9a88552049fe16f9e0971f235bf3e81b3fc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb87ab17091671d20b72dc8e1b2ba42256127b142d040459955f1f82e83a6b50ef3ca332c0cb7132bd10158e4b11ad0802017d6175844c5402d9efc91d7c436682d50c98c5bfd249543298b09f143875d7baab0b26a90f753c3377ee0f859b592a6bb4050cde38d0d31fc22fced8abfafe648648f67fc7ba9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12248d5dfbc3ebcc4c5083fc37e4b46900dce53dd39cada456516f19207979ff3642f87ef078bce8462d0c69d2f9b08dd54e45236caa5b1a7c59d32f61516b2a224b2079af2ff9455307446406dceb377e84580bf72cb7decd66415ee7cb3dfab66310762553d5902b036a1bb111b898e2f4b1730ec965588;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b0653e9fdf4a2c9f1d306088821cd94567e9da1e596b58a699e1510c843373e85ac26a7eaee5bd57f8350a71ff5cc1ef21106136fe97b2b93fcfe26d2946a6e2162e0716fc452206f2d7cb33942ad22112a1577bebfddf7e0a91e4ff084a6d83e312c3a30497ed5fcbc588b456efb2113454cf607cd79633;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1131393d72a7ee36ab670536b16c3c46548fc2a040672eafce6d7dae85a95f1cff96edcf34c76acded0135bc178db1110cd193419700434db5f0d1b12aebcb2a27284965320b57b2d50e4b3422d1a61a59356218ce65e3c172034440ed7a693e62338c29bf0bc9f6090dbd50d1d964520c2fe228ed4ed261;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bdf3415ccc828cbafce5b9c9601fa70f7bcd21d9c2ceff5b0388adbe385245ca59eba821f75222141089ddf00c8e0ae1e95506150a76224de05908fd352fe19ab69b5a04d060d2747c25f16942aa76af7b65d2306b9d2a0ccad371fdc58b3eb73667b6643d4d4ce035d185b1cfab311c9fea4630d9b2ccd1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13d088a33a3f4b7c09e167e091c9a46e439ebbd68e5f75af972f532360f0febff9e5d1233f432b6752f411e839eeb10e2bc53b8166423e3c64f0c0ab275bce668f0dbe1489d14fcb08b7fec4c797d44e607d21e4da25bcb2a838490180b42b96f2edb808459fae3c8ab4b81171e2712700f7be61d13b7e2f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17a43481cef267fb061ed08e4ea514536f14741439ab704a3dd435afe29b34c3a2d0d5886520bdbd42055097982d432443f087f9e49f667db217c5fc51d9ed83320ac4e923d8b3fc3e1164836256d58c74d8bd47f084bec3ee54a616865831d56bef4ff66dcc86ee78716d79ba48d0fadb09311dc6c2e8f89;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h64c23eb9a982222f36f411aa598b78d1850b5598a08fece84721190f6fa72c3a6ca44e7fb08e4872216402b2ccf9b6b5ba50c64bd3a9441dfaaad2eef7c55d59dcd0c6dad3a8d84fb90f2f412b22e3fcb2b1a96fc1c705a07939677165e2d47a150ee0272bf9b758008562c36fadc42dd9809d004e946085;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h106bef3908fc54231b30e009acd6b65b265bbc2b6e4978681bb261b55e99e485e3fab2fe89790954ce4cb922da0ecac57985cd07afdcebd80b905303b8b3602600c6fd65befa0cabde311c10e9f27fbec3f5bae050834af598fe6a7d2461227edbf772f0d597744f6c55f052550ffcc8d8fd71f56e8594f3d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b206c11ccfeeb31b0696acd1f821a0b28b63011729f7661c3caa374e034f3d1caccdc401efa7f60dc424eccb027f292af2bf3fd0406bc29f5aabe3ac0c6d0374a1b65d01571e3c11f94981b63b24c9417c2d7fd747cddf8e24cfee63e4af221681d4fc81f489be46be97f26fda9d80ad7f9baa689b8e3823;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17cdec2e03ae1d1a95c8b6717b89928012f7065a5848463e7a0de0059de0ee199a4651b87dcd73a1aa9667f036fa94b14bf2ec83e275f384cb3671ff06c8aa5600b0fd9a5ad8716344b9c6bae60bb1ebf4476d3faa39810cdf097b153c7104ae72ae5661156a200b6616f3fb30156faf654694b0e7a87ea1e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdc71736ac6e0133cf7d49e411aec28e466727bf8b6ac681234083b8d7712d0ab77d7defc85f5462f34d1d3c1ecc5b4a0d21856c2e9e8380b265843ddb607b09ef8d7afcdf5d61e6fb41f417af73a4875fdb6ca207392fbdfead76c308f0f811411ea9507c709bc15c6a3d7ff7d31aa39a9928aeb2debe97d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1228ee9895c8d4a7a4a2581f82bacf486da94ea522fe2d332fee72a28275833a7af3f3b6548a409cb971a77c0fca20ebf67f9b2ab14058b1aaa0dcbfe2afd95e101342e7c86c2c28391fc8c2bd5de0c7d02845678e519231fd50685ed861b43259eb069b69e49e70722335cf2a084bafdf1f76b86bd9f870c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ab7e07568ae53d4f8e1f304936bfc2ac113f99600e74ad2386a95dfe60459f56ab04bfe831667fe18c7bea34aa458650e7f86f4065434e973f241bd91813c13728c8fd647a7c3a6fa0aa606b10c7f68f42675f2ed3b55fcd0b7c4aa8b047777f8a8692620db80eafc3e39961aa476fdb7cd0df19e1d73f5e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h919df6f3e7382ead9e9d0ad43d923ee6927f2bef771a5a7767fc7af0cfc197d4c68f2ec22873c2d75fcdb479eb2d9bf6b6b221b054bdb3f6e108973dc5ab26fe09c1223bd81d7e5b1debc03c8558d1f5d95b147197bb56d73dab60984fc74875161f32f5f5241c3538f786cbebb5c2d48a911a6c05fa81c9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15db96826b33db65977a2d12f4fabc2e20719974901c6febaabf2ca33e87d635231f197980d83cf10c43555d2e9f24f03b0f71859d4f67e094cb469e66001da6e43976f05278cc11ce0664687cf3c07c41c577e55bde1a81cc3d0ec6a1d241fb40a8658a5271226b82afd771f18be5c88e8595fba5e767d3b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfb500bf3f193830911f6326f59c494310fd1140fa3ebced48b4c8cd5eb49d780d41d9e700d61ce4f7e6cbb550a634a536d16a7b001c5fbd6dc8c195f51fe6b8d448c6cd1c2ea4bd3664acd530008054d7894dbc49a3a471a8bc847fb9dc6612268138ddba689b530f73b40533e7ffef1c8deeabe5eb1fb89;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2e0624439e847ffcb2af4e9752ad9459901382ecda890aedf26c5db2bdeb594e629576ffaa24ac0511a67d2f3c83753a9302afd1a9b1bcd3da9c9c3f02f7f830175c8fe14cbf3fa419e137728975a8ae54ee1cc6e2687d9aafb1d9b94204f5a658a027ece0fd2599dfd0c907fb72c87e2375cb3ab2d1b1fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h111d7a38f51b3e309fd6f9b40e52f2e66bd13f47d131cbcdfdf94139265ac202e9b0139cd1fb094fd6bc6f0fd43ccc9b8eabeea8c6f6e41c2d4d62fadb6f7e07d9152611ecb5fe5bc8700fa0c250cdf37ac32ba377b6882fef6f8bb1fef142d45754410807e00e763195d6ea363bb494fe0a410688352dd4b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha431d40274a65d2e4c36eea63afd90aa32df4492c7c4ace18a539d04f87b24c4d78c5079eb5b3e498ab76cf0c4ebebfbf02bab8530b9727541e4c55069a1d05396e8e48e9e301d3c9a96083e43ee18c3fddf8b3d63b33e908c1446bd3919297ee588b6eb25772719d6d226358a4a596b851b20ccf31e9c09;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2cc0e9125e9c10c50d1a977a37ac74fe43267e5bb44838a790a714e59e0e0acc86c6655fffeb9d7e08fbcf784225c400f749060c4924b95f7368336b6342fe136ab4327b7f135c9eef240c2b712565ce1c4e569012ee3cccccfff0c0c366bdfd316a7628abcfd72a6003b1c8ef06d2f567421245fa72ed9b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbdd245eb9eb39801b16777a2b35461dbd2de0cef9c90869213e4f9be55b015fa8adc3ac76a2b8f91ee66b65d85703817b4328d2b3dffa7783bedf609f86a8e94b2578067b10260aee6c82d86f2e71c80f95470b39ec1436f94103256a2a8a1628edcd6d4b93022aead1fe0973eef9aaa5aadbb53eb47c075;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15b85e8083513bd367659cd814bdc38a0ab9aaa23ccfe563077a0ffe723568d4da32f9a3ace07d87a13d0ebaceda0cf375e955622d2f37537c07c914c0fd11dc0cc4694d80543b5643b0a6f4bae84987755c599debfa485421916f6f81b59d904caa56aec39aa81f4b1f6b3e115df9148f931309213c3af56;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4d700ef648fb360ed3d48a4a280b4a9cd5b43082edbc776bca6b45b0ce2016d913645c9d5e19e1d0c6d29df718995aaec8041fef39e3ac040bf48f68f7884e7f8b343c2455569a5bda16d4d01f1785114097b419c6edd952de2c60f9c977accb42534676ecc8e44ad34841c52a0597dac4216f5db021e59c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h133e336608a30ce6389eb016bc06ca4f501ed47673a75d85a36ba648f5193d8d8a08707982b5e70ec2ba81cd32b416e7d831fd524acf1c0b48a35d96ea885b0766f9a52668de183fda92b4f60a208ecaf2f20c25de4a591f7607a6d46de07e822ce6f552a7844d26c8a0d538289668cd5cac9884ef0137fe2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7d5e37cac615690ac5a191b417801dd5ab1577bd7af39de7d6bee47c0d4a94b248e497c117e667d97b5d76d6fd2452bc03b2e485d90174328c6ad19a4ab602b5d27d8f32cfc82adeffdd50bc1d2d9e48904ee91f18caca2e0789e0326acb449b928378fc88243b2df14598168b1b6c73881f9987e03d0460;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9c742656ab28adfa153d4739245cfb2c0caa80e43a5d8afa03d7eab994e01b733b22840afc566b86bac54da1d016f693f0db50c7d8c7084209dd30f2f2538486312bdc851e79221648ef4cfb8d1221a925ecffa0f5460481eb8cc72f9862dabda520d34338e022993259f14ba693ed6d994bf54ef2b5a96e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h122cef7b028cabe7e71348c7fcf2a9b44ada7b116b2d22261e01758f0e35bdbac6eb5e43408f6509745c54d402df1a2ae5b6c294a36c2d9e431e91e8656c823795d70ac3db1fe933d67100588ff708e15226d6327203feceec5628a9f0617bca39c309648dcb1e915e2fbbd20a9896c3dbb7c128df437c371;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h63a9b9d4234c3075bf917a0967beef31228f58c54cbbddf6469b1e1b84f9f01ad9708dc5ee704295c5c8947a6905c5305a63f7e3097f7cb16a0523c79689209d5bb91a0c8d5692bdcaeb90f62828e7b89ec55476c18ea6679d7bb1a4a8321ae817a8140e8c3c6e13262a697ff630632a253d219193ebbfa1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ab461166c6d6ede72c7f2a2b7704ff4d2453e9c997c18e08445318936b734340dba1f901898110d5556fe6e6261162908e9313c38be3ea5bd6932d9848290ac75ee3ee5e2a2af3a0ca84cef4a5bfe7f4df01c83a1037f319350a5251f74277bcea75ceb0467d8bfa4bc2169b6d01e733f66a9647f2ca0a65;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4d9b873c491d3738a7530e3c83dffef52662124759e66341b6239e4ab84b2430a27dc7b43a85fc2dd310a1e0fa1be0bd84bc5ec221fe64643f77f6ca461c7c6fd518099f0c6e985510d97df9d39c191ab7db3ab1e9d24041c6d0d8c3a1b7d48200edf89e9f555ecd078db9b75e36a69c82f73c16594f0a6a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cb1b6ed5f765a754e31f5ebecae7624b01815e414b6629cffbf4bcf444ada6cdf7009e2040ce98d9abf657cb319437618f3217dd4bb4169b710ed71054daff530428f4cb720bc7a7ad1f7665e60427d73cee1672c0348ad980fcf515d931449489bc7c3b82cd068fd13d6948bf55d7ddcbbb85b248cde221;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c72104a9ba053af58f972cc35d39b324f2b471a47e0f497810fbec68e28b13387752d019a2819bad39661b6fc21f49bca03ea604a030a19a1bf7e39ad13d42111c193e61825ad4abe687dec4c22767a325c7aadf8eee34796d1d88c7ec934aa02ac2444abcf5a300acc1a485f089d325061c5582aa2f74c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10d645599bb88e4b93a0c140e27b3e2fb21914a7ee8e1e0fe7395441f673059dd4478f62fee3d5c6ce50135e765b4a05291aee5eebd2eeb6a767082147e8eb0b4167a622b8e8007a6bfca31e8da2237327dcf788cfacabe35c535a3477f0aeecb12151e88b2893c4ed363f243cab898a800bb430a2d8e0221;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he99eaedd1cf06404c211e8f1deed2532d4a1dd96d5493da7329d8e45cf15284448f147454bc070f16592c6146310fa6040e636edd02841d67c17f4df5b835ed62a25b2bef5570a9cd0e8ed01148e6cdd47d2e335033b3d3609ad660ad401feec950c38d7f88a0c6e67b1f4440394daafaff19fcbd7256716;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf3a7f0dd0e09a9c3acce7bce69be9cba5d0a75d163161cad260520076da6de4d8ee739a2a4258df84bb9bbb1771773e4513c8ea277541a6b29aeaf65e7c58f31c5b70d1cb9cce36b106e355830e02f0eb6464919d01f92d22edcf5aa6f8cc550ed163e1602bc529d8b64e03bae9339282f6562ca16e4898f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h164c34dbc424a338abce26817a040737194a4053a2275955e8cb81716c375a38b8241bb55556453aa2e4f4d53b7a9f2cfef13469cd689a539e5c53e2a80b0b3c6d04a109abd612c12512f148414119029664035d401ebd4548dc0ac1f982a715cb65cb980759d96a8fe6b06b743437c076ac954c8ce61d7e8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbb4d655118c675a89e710158c6cb9947d13f4e114ddc83a8bbaea1a138320db357af065e098ae6537a28d5eec1e7ee4d5c3ff2e1e8d646d221a4174bfa10264380f1893d62ea2bcbf5920ce4889241986ded021b85357e7d719f8624c90630ee2a8e0dc62950726ad2786f5fb2d91adf6d7c1ec32ef2990a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18519944caa781cb11169382f7e5b9c3c2630b6d9e34e31391732ef9a3e2e794a585235145327beff932640d957dd2a4abe46f3ea768d96c81120c7a3f2b9927458a3aeb0935cb3a5b5a29c5a7588eb494855379d21e66bd056e34a1e6380b271c6993199d198d880c41de5e6fa08ea1e3413043caeb08edc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12d4df579b71be8970263932194ab6cdf502acc2097ed5331d4d1615ab86c58db30da6bfe7c68e9d9730e53bbdd8653d9287a6273d63c6af580e3783a5ab936ce4d5d52beac08d6ce2323dff18e7220e2426fe07da225102ee50e63c353d7ed9b9b1eb283990cd999dfa44ad8a4dad74f32c39013e037c950;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5a5a4d7b8934bedc17366b4287c8fb46b9102a4a9b27bb13f8445ca6ba396040e5ca586f20d6c90d7c3e3f8715ec15a81d1edb3875ac7804302df312da2fdd5d6d4752374b8a1f6986f4b350d77cd0d7f20dd3cfff55ae249d53930503f5fbaeb76f592acc8d287765048708c2b8ba4b230588e091068297;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146a9a5dbc426a68ac46ab56e98662232dbb5becee9202d273a6dee4134a673b98aa2398ea2e626b01e9af7513f348f55480a3f68a1f9f98d79c9ee51164f2d9f60d6499edbca15bad300dc8bcd9762ef3200f65586428058f7fcdd11328d6599fcc518c19e062871fad9ba221d94047b71e50f6ec6736078;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13ed4c19521a8440615b39091ea5ef0b6320f67be2d8c2ecd63b615ffcec5437673272d1e619213b7c85c6f0c4b9750ec5353021ed6a13fb6f5ecc4e9d4bbbc3e290972cb16c15179fe1157c517b8d38d093f82118717ae8f677bbe3d5fd660cde6fdfa8f63ec0d4fe67dccf9ee9fdd8842c91a87d1ecd16b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ea03617e961230c7be2a30bb2c5bb4516c26fa741bf5df881f950b375a87c7a0209b4476a395d927a7c278784cc8d4683ecf2efe591755cf72ce4976f6641e1abdaf8eda94427261dcffadbc03f1b2261b2f7e03afdb5ad6c1dd3adec132acbced5435d3cbd3a9e6c29c3ba937c5918ac934b8f0c825dcf9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14bb787b9d0a8da0bf5c8b3813d24d95a78dee79def894a92846bd27f002eb11b00ab3a836035d05e71cd7167db932f5d99d508053b25e323c1b1448dbc0880e6a56b2b188bb48ed55b36fd43f3f02c71370d8c4fd240cdd95047771289a3f68291b25ba9e775c493ef9162fb3034c303d4f70f60b29711c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h24320fe43790426cf4bbc932cc65e94d4440fd82a646b29818ca3e0bb354990a2dfebda8823fc1161c102077261fdc2d62d46291d8c8eb1fb143d8b8e4a87711be905941f31679837ce0ffc8d511e3ea0d0d1776bdf26d4338fc247c31d5f54a0f2830ad6dcac11ed4f1ba80252c240de56d7c6abad91292;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f937c690bae7c309d805be703fe6f991ec6145fdd85a915ce64495f2024561e81a3e4e926da32e06cd1bf6fbcc137b11acd7c27171f578c16709d5347be691f2ddafbaf9bbd7404a9de001186820e7e25b012d52e45a8fa008270196f8ad59e6aac87a94761f6b6f1af02daa8a098b12df96572a396f9749;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbfae1a6ad4bab5dc32264a45066dbd0b5178fc66e38ec5831d3fce1f06503a3296f3245d62b99f3cfed65f7d2114d2c40d6de241dec16db1d89882d74916d58dfe65eeecb0037583b80d9f9cf8e53cc6a3c2ef35abf4ab90d45e1843401df7fe4da92fe014cefe0b5ddc7b0c77b6e9a0cea2c4e923907c6f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h288422b02d4c65ee6d06d4019a13925e12482f8ab45517a50cffdabfca859e6ee353e866a66c49428b082fbe1992ca263bde6a0379ce762264f18e6b6bd4b757a7164d5d6509fa0c2244fdd53bac5f6ed8efb76617d4b7e2e312e422aa40eda146eaa0fcf6617df6af8a2050110ea6ad8a03bfa279cf9387;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc264d80ddeb1c902e44a90624bf8e1b7877f5b0b0fff50c686c52816fd5a0cf4add07e1b732decb6d12000a4fce2d343240bdc9685e70c1f00ccadc310218b80f3826cd2877c1ddeeb1f740a7adb128d5326bec98a8d3446924a4deff1abc7d44bee53599cf9e8e03b287bcc7254525a1da898c131b524f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h165aa516e6e0c92d919f2456d66bc2d30185bf25894b8cd77db63382d509df5bfc7e0fbd8f9032935a44b9a16222aadc295eaf217770723e5ea5ffd559187b10fb9331beb84d89c5d190669a66fd828039aa08519d3f0b9c419ef684f3c2091cc1ef81f2b5b5bd16140cd4e934197ee7ae7151e4a5e5327fa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f2bdef812ff7197a8fbe385757263cbb877fdd7651c2e6d1e520eaf3357f75ddaa6bc47cd7230bc1f00c788b469d671c13461a1e21a305c5e5291fb955eed27b1c94d8dab1560dc587bfe842323208c49c6974a7214f7dea109a970ac66e8da481c4e74a5288a27c1297955fcb8d13af2902a21afac9ca62;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h401a8563ff1a2b5aeff6f117504ceb02ea75d120e7a2596192aec45318fe7a75a9988b2fd9f5dc1d4f6fc740adf3546bd276bdba4c61bd64ec25e5221863c21644a19c22197c711e9af5f9f31425d68513472352917b690e0471e63458f6268bd35c87d9dd94a24e9cd33995611e9df7d97f06fdc44f9500;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18e8c64d958edf28064d6ea23771f6d3e64daf32a51a9ba9d7a7e5d413fa3868753b71dc63b75f1e764eac8919e41ad2a8d709460fdf75029c9dffe8389801a1118aca0af8a41be077df3530485cc9b9c0b4691cca4c2f22b3943e9e495947b6b20109b6a194ab01d5041e5d84c11c1add7d5f62a11033e8d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h587b97d072fce364b19879874cc2f9141bb7ecba516a40ff2544fcbb7c86276b4b49cbeb7f490c29ebe2ea2d3c48584c023b90ebcdf0f42fb2dd57f85997badf87fc7ae01025046a94475d46d6f8b2767e1838f8ce237913298ab85dc3bb88701537b862dac41080726ed51096b84438c617aeb697190aa4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc8dd2374bbf18a20a66828f68154d3e97bbc4ba3f1b85563303365e87e394a51b13eda4177394ef9d830a9884ee2db23d80182892629449bd6a65be3835c35a767554d950fc895b05516b8e509971cf43b644b0f0774ce6ee5bd66b39ebcfaafaefd3ee1edc51e0432984287fa44073e23ab2c7abbab64ec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14dba18364417bd9ca5c0a3e8213f479645cdcc343521ef17037471e312d24b81ec9af79e72f518c1a9b08d8698da0795626c57713efba090f11d248ef4ce9dfcd77c538b4129f708d990ebb6ecb628dbaa2f3fbcd8a25e6d1fbcd43690171d294423dac36f0636a9dead8ca63a6fa969141ede803a19e75f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hadf037fe118ef93f7095d7a0eb20c100a64a84a82d6d078a8ea8dc2ab5326b4ee4cf19cd58ea9daff0a330fdd762b5a5c91439717b8b2a49cbf9ae9ca7f7a7465ea10c0096bd3ff0c2224cc6494694b767d3cc92d0319a81b8258e5531fb09a9038337d15f885eb734f5faae640a579e89747fbbefa475c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c703c8abdcfa53af1be39cd3961e1637277345eed5a4d5c3d7f59cd0f926c3bea7a469e7f66439d12deaabe12e7af0e3024796e7fe50f853f11bc68e82d147a4e319b65fe3e1f0234d32b3f78df22adb6410c8461252bdaf972be865e1cfffc4c45b14bc1517a597e580af8a3df2cee225d99ce9b756d9c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h53e6699b94202d82c226a586638cd6228f90a3615183c798fbc465c4f5120dd087dcf2db71432882f9107a7180106e04fdd064fcb95cea2240c20f27b2d76fd8413d6b99ce70cd96925af4d67f5e73f49570794e9b05bd3f8227ca9d9c1ac91ac5664cc014fca4949f3fafc46febc96b582e6336ad3fdca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hae7eeb9f9a3c53a3e9c51dd1d55090f6b6dcd123184fe66beee59f8d9c9002bab7c6140c1342ea112eddc66df996507b7c183cfdc00db051be278685009be5d21af1b58d990d16933485c10dbe194fd9911eb6c4c629c315aed04c14d83314fc4b7c6c805d640a45fa6943f24b980acf01a741106b98fbe4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bfef83424b982091d0b83964b279e902692b40249a552267f739d9ce3459d8540af7a507e47802f8f7cc36437e43f5480577606fc1a38bbb36155a4eae935a287fc9799ba25926829cf8cde6ffd7740769f342c0759058b2508d0d204d24984dfeb110bf0adae267955cad9b7384f5163599920a9aaa782;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1da6bb4431fa9bb9c49db52de545a3cd5e88082cc1f9965b2dffc0d487e3abd004e29a82d8be1f0d6d300f4a3d7e33ae84588b0f64a922f4dfe7830eeb8143b6978f8ff5669c5b008caa7dacdbc91479802a021c3bfa0a80ed59290cbb496a0a6cb3a5741944a455d59915dcafe51631129ea067cad8fa1e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1668b0ebb08cc9ce06a651c0fb3b64fdb4275b982b8e759057974e2f1591afe358ca29892b39621a0d6803ca41fd652eae75a02653719294491f99285e5b0f6b2f500f7e6ee8f70c1353e24f00de81a23123c89d5ebcdfe98055b9413605578635a7a841a328ef49dd4a4574adf37229e546fce5f38edfb35;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h910d20ab8cff65aa7ce98ded5c4bcba7d85a46a732cb716352e40f4ed31ac5810e751d5a6f19d680e82f0a7cb302525e6a0f102236662f96c274e2518be2f80f060ee3f95085252ce08bccde70df64fa92fda0dbb70df4a6037288c9403c0e00ce84ec54e6a3bd862c59696cda770e4389c5b386450b60b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11cce9745f15aebe9c981b43fc848c67897c740705e655f79a2bab7370a1a1d571cb35d06a18fdb18a054a7f6af1535f29a51a801a94b1b283b86ff52fc8801fd0fa80cb181bf7ad30dd15c33497296660f4291622f882ca4ff1c84d138bfe9ee10f988082a47e57b602f0b06245634e2b78a5ff1bf290a6b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bada92c748d7ddce451b4689ac781482b96ef8c7c309703b50a7f5353a360c9745495250cdaa7fed8a34148f7d1a818ea08f77512eb01b2976e7158e203134e159fd6e3566100b3eb29a54640e28289e6a488bbd387f53ea3b93f78308629a15dbe1e9d31601aab734d075b0276f97e7c31b0d0828e29e51;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1682707d3de11193d258d67164ca3fa58019849b261dead2e0046dba5b18449c104914816bee8ece7302e4399abdb1c71c766276de6783681bb6932b6269fcf497e5e23b579e05c40278bf9bf211427a5d4175043cdcfbbcc185e559b419d5f9f001b7cd2db76ed306b00095e82ef63d379d60d9c4001808a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h138be421a3da4d27fb640769131da378347135b9ad081570bcfeb3cf25f7b96e520950e1799019b8e53f4afb13d1e8f20f9eaa4eab522ab92ba90f2e8b8b11ad6ef092e76a2da4c761355c8309b1ccf0d4f6389a022ebb99dc2cbe86b27b8de9fefb8de69be8393c0e8b1b7e5536d1b77aaf18aaa4c91c750;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hed864aa615aebf1563b363d91708ddd00a9b4d53be333e3396ef33b585b840f79883148a15420d77c7b8200c09588a971b9e8a85cb581f90246fc8e879cb4bed71490abe3739382dec8d99068ec361bf772775f506c52baadf0fde0ab6c93a23b8f8a2baf6b3dce1dbe537e6b001004cc2245c151508ae49;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a2de216b12f64fc73c82f0eac5e17e1ba73621ba1ac89274bf315e719b2dca96a57e1b210aa8604cf8e36369b13f96f82242df54d123651742afa42435fc7917bf082667d5ca076c6e2f148701800cd1f040e8003027b16353485d2760876268835d94ad2efca365706c257ed4e5cda32c574fd61214c9eb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b4de58f4d42d8d8fb7620219f6b838e270cba258dedbb0e6a665729ba95f2f4b3e0818192c7c69c2bd759eb281e8e80a0401083ff6d1c794a53e2cba2c98ea94dfde74cf1ba00c01119feb016941d10a3b2fd664e6b45a7a576291ad5a3da7f44fa60821fbaee1c248b562d5599146ad8a1aa7977438f04e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h191720f9cdd75ea97323e5f02a34f4a0cfcfbbc4740b956e638f94379a3a4aa5c3494bad07cb909782482139aa14131920cb07a5fa2b9593fb1fa4c1543cf71f957d83d961880abd9e9d80db23c55ced4a6c4e307be159539ce9348c4f2eb6f81a4adb6d1e61f337099989cb866feeba5b9cc60eb7961741;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h115894a896eb813e0d9de62b5e741f5691f8b34f48a82e0576d949b08786011c7292c3999a78197905c3cee9c07079c2e55182c6c6ffe293352e7203b04457009bb9f4ad7914f7e5a023ff8b12fe02d34b5e47e8c3439077e943281f60ee9ca607b890ebbd75e78e849b10083a5066673014bcd1fce7cdfaf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f8e249cb9edb90d766cc8ce1ca47558f313408ea66bee9b3142fa66cc10590bf349816fc71d2317a3cce4c4f16b12f346a372328adad72cd0e819f17ff3e06e480d77031e176d2db9c39ea776dbadc27459fa3818e669c654d31738521192f0a73cfb961af6c1714ca277412eabb0b9f30dea486da308a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9ae652316beb94c1ca5b4652eaefd3632d1275f11371f575a02d3b9ea634f33b758842665b0daa78e484b2a1c5cc9bde0dd13122c3792f682b3574259d18d4152c1e619fb726735c6e794d984c2311cd0aeaed9b0b7a634068d9f59aff0f1cb1fd395b0de5b28db9d458cf9e908c1b194503fd78d15210d8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2696d2442577e5b41c42b9831a82e75ab2f886ada835aa59802309ea9d2234ff7ce7bedb98348bcb1760892b725eb5d3618cb7e74679be9b09ac549ed05388c7da80da74898e8b2f2163a9fdb4bc8d345f0959d35978f02228c3f4741fb486a63588428e7fc4d1d176de3c1d2c1014952473412c31a42629;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b94eb5312bf2405e316d4086c099798445aab1eb0978ecb28fa81649270b39f5a87bd2bdaf25ca5eacd5456f2b3d54a1f192b62f2b8b5a78b114d151a297dd2d934a264a0688e8b20b6d82b61c76c41cd0d0517611445c6b92847376eadd909285e14bc1b5b14e782cb4fd888f20b1ac5a2efd9a9c8e7ec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c8bf1ea895e7b38771d32702bbc66856b3f40a9fb4fb85b50b6d628206e7daab0bc894de233a2165808f12c980c731f4a5d702b0a0e2c977de2bca1202914ee7606a0c562acc4b9680a0963464b6a191f6dfd2b8bfb3786193a2bdee8f00873d0b08ed53ce61cf56c099dab9c318e09ca3915e9c007632f2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfa0f4548b9af270b092428ead39e1fb8d4dc961d1bef89b556b9209ae4774c846c160909b8f45c436ba7ecb36ef1405a8267fd737d93ea7de2446a9689caee94c760ce656fdec53d4288840ac2ddee35ed9c144a66bf4ef6c2237e9c3f1f21ac77b7ef8d3f200545368303cf157398d6ea6e2d252f59a449;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc9fcc40e6c27e04e4b8a0e580f42c9f52640f8e15491db271e4779e78fd73e2989e23bb428252e96731e44e0c8cdc49b8dc8c3605ae2235b3a4a9284db4d9a2172e889c20f56dfcc64233cafaddc473d340d3c4df68eafb9c14cdb2483f9ea1661c27549762088741ef30f02195e1aaaeaf93229abed5d42;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d5130622b3c18b88fd97313244f92d2a997efb6d5745bbabaf341fd683c9b4da5bd932c87617cb274cc6f95987788cbb237891509d85cd80176777e03b6dda5e97d1315deb1bad9d69ec31c6e1c7be96ec14392b34d540c22d79df4bbd28e40bd7d291256a4c68afdc628892df7cdd5eafd90b2dfc312e5d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1493cb1ef424ff48de684d6d1ae7abfd3ec01b6f5a797a2ac01efabdcf65761e84ed545d7e92684c464b39ce8241643919c1dc44de50b9b1bc4b1315cdb1efef15b24d6099dda7e8b0a9881f75ccc0d657f8ce5a303ff705d12bc566b02cd89d60002e193979b62d6c2125921de578276127a49b55402b44e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16bad703d49bbe2d3c164446e0b24d73a4407ed641e8c53508f43c17eabcebc5ed04a2f375cedd4f30fa8bdb0b1eddf0f2d361c7deb9d3ce88bb362bf0139cdd03f545400f26809ebcfc12a33ec3531a18b03a4d395a4701edf9269e9b709f764b6336bafb7580b1f156a36cc78c25385c2cef2b8bd4e5513;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h449e83fbb42d05940f9b73c88a3e673725b7cb7c28e5da77083f8aacbc57f754fa1cdbbed08de591c2132b3245757dff40a315a352133d79fa943ea08e45d58fbba599dad912b48ac10774369e995cc1c7269e2693329f6791c610de0ef67d79cb6f76435d60cde51e2d103e745655e73086e6df04f0bd7b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he3a2a8b190370db1cb724eeb116e933a32e20a1b99bf541e149648e816f7e9c312ae2c5347e7d3951f2e74e111165625fcc44a7ebe29d37153bc4f0516504c94cbcdf31c38f61f2c6264508a7158c2ce3b13ac0c744dd1b0fc00dac7fa47eca231f63eaf93b120fccb1c9a70aaceedf150ff0eccbfe7abe8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eb7d1fa13cdaa64bf56242281992b794543fb2c1f1c295b02094a709524a9c2ca0bbefb8480dbaa0c34a554da82c1f894f51e9f61f86d05f5a8160e2c3a1f3f0ed02c0f03f9d60219af2292a16cf63c1ae4256148926bbcb8e242b8125a7f6ef56d03e9bdc1a5b6166aef5407352bb04ebefc9c31d4c00fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h92027b937a86edc8a54f220fd1d70a2a02ccea9583a78e3897b674b53d9ac10d09c5197bb504c85c11497ae4a73a6e360a7b55d368ed83ba81b85d122ada7d47466b07732fc457bff437996205cf2910d4439dfaf9227750211e204f290e4a70921cc58d7c9316f2f8c9aa32f47e5f0e5b04fef1b543c3bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b715f275064015af11470c3eafb8ad142d3a86d701b296182811ac0c03ce14fe57b90f7150081c9dc98af18d9816842fcde42053c856a1ac6b65f8fab87cba175ea715198ca65a5d867857afcfe75a53448664b17da28fdfa8536dd7d143ae7a92a87bf28159c905425356fefdcde3f34679d157884bf7e6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6c5e45208194593c1688e9ac8ba598abaa89bc860de6db2b1974563dff08602a66dafe98eb9daefcfce0fd78f0bb77dfa1a51f75ebf99a16f97ca25303795976abf0c2787b2eb055825c7abf7b7dd31c75a718775150a1fb37fda0435e7831ecee5112cb46491dbe4734ef5f15401f56e59fc88842fc2bd3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19a428f0a0d5b39a26f014dfb922380126bad9d23a9017ca1ff095f046a0d017d0b73df5d805ff3abe6486d1ee5fc6142677dcf1671bbd04eabe0b794d11a56a212c6d25f524f5ca22d19cb598f368eec01f45207418c6ff9b87668f027d008dfb4244ddf1ff291a5aff456ccd3898044c1f710aa4ebe3944;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ff9ff307ad9f96f25ee54eac921d315146c1d5f73728cc0ae1dc19a9fba87e48b8e47c32e2cbd9bd8e79d501a47af966b20a3fc3b45659e42148bd85767622c9d928a1c2bbb1264429965e638fc941427d64433eaf6e5c94bcb5e4ac91f9feec6c88e361dd3b2a6af7237ce825e612d5849bb1106d234c4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1550adf8c28e213c22d33c5c2eed662da06c31cebf280ffd1b6473a6f28dd14711dbcbc0481d7845b32bb44cacef38a78957fa00ded1ce61a21e9badb962130f5cdfb017126f2081cfddb0a9104612804db38187f86834b9e3ccd99f226ad4d7effd1d2cefde932424206c9f4450cfef44a680175b240d83f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hea4c5e9ebc088245a4eec1d990d500ec10e6540b0218af1d12e3f87e5633588e308a086bde625799e46c6b63de825384166f4a73d75cd9647bc053646b4d29d07551c4f9719a35ddf2f7a6c69c4d06f89da05164dd391303d0ef2f6bc120ee8e3eed3adcac766f5f0a0aa262ecc731465f706c5f505f3242;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h61a945fbc1d7eb0af64c4a48750d9f71758dc54978e5825c5807e0667cac032cc8a235159584cecf16adcec6e38961f46f018996453db7228d44ba34eded15c9ae1f7453442a91555b8568e5720602cef2323ed28afedd0a32bb97da78cb74da3091f3e3c5daf6be04ad726145f618eaace38cf29d4f3d60;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15b088ab7890fdbf2f1f46ade019303157cdc25a4de280425efebf19abe7c6eecc33c5bcf5d31abda1601105869051b168c6e2b2ef19206fcf52a9666b7aa07804e646326f2ea39da441e8a7a6d0b5a78a4791b672b592500f5fc6795d532a5ed8a794bb43621c2bf429dfcecfb4b28e61fb49cf8263b2111;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcbfe1c59c1521427678b604e8294ab213506900e409967c04d371ff697c7554b3c2333a7dec6f1f548996f9cae4071a33f6f5235896b91603303d2981d2c6ce7281c8d3ad33c5ac1378020abb5d3c7e0f5a06e5f920e6d23a2e6a4968918e274e7398c0bbc24ab18d56d11647f4a3c8573e7f5d8017c9efb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h43479a8220ec2c7fb4e4504f30f6fa7dabc668711a4b46a37c0558441c027984f140591ea17afaefb7860993cbdf8111bb9884174224b5a2e8a6e37152bf95240f698b86e13414ffc2d84d6a2fd1dd4577958288efe38491133aa00b45e8ea97406813d9580bb08d3cb6fd9af74fa6f737aafff35564b014;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b47bf9ebfd5de3b6b3f8cff47b42ac2f6d52c5c8c80f339e2e38fb57bd655a6cc81fe5184a64697ee506fc003f3f4496f7d7fcc58519ca5636947fb00af4ba163b42feb382f77aa014d57bac19fc8a9e2d93403f70ce99b1e704f3a8b9554c3d78a1eb3ec2968a68be1b3b9adacb1752f4669d36b871e1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cf2a3d4efbdfa63bb8a7defa83e0d09b9b61a5c4a3d6aff79a16eea22ef8c2918be914e242aea32fe7c64c6b078cca3c7e2829cb530aad379405d6bd17b196b339a9cbd13acb19f66bdfd259621ac10bd829d0d1eb594576513c3fd2a84abaa5d3c9e69b251e5e5a592f6b3ff801c477dfb090c449ef6638;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h149f9e0b240bf229638ef83f326b62637c545f88ae7e0e7b206238cec31e6842353cc4b6f70f1f92f3d1e936bac33f1a9d57d4ad0bd5e2ebe9ede79978e4403f07f29115ef726453f777ab7f3e8b111b948cf012be406509efe053108c92b4581259564ddfcd42528fe7a43fa5cb1f154032f9f48f72ed36d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1580351ebdd9509692ac9425198f1e74a8134afcdbc8b9484e88d084708ed3838911103f41a680e6cc16460afb6423559b242235056026caa195b89b893a7e5dee17aa4cd815d318849866ef7f1d08ac752d010e697f06da80a45a8c53449858b23355ab946d1a4de492b8041c53e92237b8dd9feb5f98941;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h90a5eca73e8a2a46c876321385d9aca9070901832723d8627a976ab56cc5ad4216be7a543b77ac83e4ebcbb98d25357b83bda02a1632758d3642ae3ac3b83433555bcc8bf29419f326dbde4d1dee12e330242a9e68710cafde9a67d4b866154afad58a07b983b22064987458334be0c7abfe7e49f2fa163e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h187c7ab9cd158b6716231f6d937e647ee3029d5a889b26cb6885d126d8d90f15e7a5aa77fb0375ec018e9a514d089ca7ac5f21b3c8ef9c3004b38aa8ee5e3dc955a86ae9403d8ee77c1772896f94203d67f0c83e4ea787d8de218df632115319fca7cd35d428f05b81a144ab18ac033d80cbbe0099022a823;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19359d7b7444c680f03e95eca32913b33154b08308a384bffac090760fdbf2746b43e4e066c29aa5e1386c25e6b5bf24051e7c6489fc153ad9b6029d9890fd1d56d829d91ad4df2de11985976753b948f52b7156d2705e4365eab688e17ad480113cb99230fa3fdf55a6437f1420e7be74ab68f658ff9b0d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd5c08b4e76f078cfb063005b69498176bfcac0b6293708e22f62eb654908b0d18b50f41e9dec45ef9605e4fd336415cbb05d45606aeb157fd567dd92fb7bd613e5aca119c60dd40feb989803d8400ec28a1169a4577cd76eeb50a3707982456fa93fd8fd0c011523381bfa8037168ed77470cac941e138a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3d89d1bc4a6961e60a1a3c3fef565939c861c75b9977a7ca30b42eec94613214922c4872bb385a4314dbeaae98c9453a5fa7205ce528dff29ede55d5e0b13f4ad33686f679a5285af15d8cc44afa9ad3261efb43fe293273cfa91f6e32ec122cd25844d22c55d53ace69bcb3363a2a272420acbce8c02dd4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h197a65daec24231d0e23f67586c459f0be921e9dfb6b44c53d6bd52f74dfe290528c656851bef4c5bb6af10b57b519f5fafc55959f79955a91c5fda9a096987cec87a4c088616279535c1fd4f2ef26f3ff89ec77de49737fceec883504ec3589df509418baaa8cbbb9285be2d550d169d7c14ab455f86a353;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12b80f4078682718961d3bc09fee195cccbf77a7edb05567efa7374d9a78abc98288cf020b5d8aad9159e00bc5dd478f9f621346825eaabfef2d2efe686ab2436f42ef52e0546b76bc4dfcead54112cae0056955b33533783c30ed8b8058c90448e5bd936f25c27b0c824a839e5913b16ec6f1cee32de9f75;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hee75174deb8c3694c1b4c55aa87af96489e041d7d21f6867571c58e2553fcb09197ef9ea048e1bfad72e41805083f51c2a2b679f14bc1c201b002cda3737a21ba0d42802700ce3a431034a28a7e141bd71fe265b5922b2e9306ce80188eabf81a7a241f2d1a46ae4db70a4eaf567a7539d1489e02111cda9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a30955e05598806682f307a804cfc6a2c8066cc70f1f95bf57a36318af06aeee75f87a82655ffe59c33ace0e25c9b3777786746716073e32be8439d928e9265cc34fb9fe0b6f348e73cfe02a36f27d4e94b4507fac77fd6a4f27e3126c1d9b1c535a7c81c11a5f0d416bc20b36f5ddb824c9e0b748d95402;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14f6120121d00fc71e71b886ea1668d7eaf1828c38f34e234872eb225d33ecd1ce5614da44aad238b86be180f7af613cc11749a182678d31697a6234fe354a80f16a90f296e4cb4330b4f5da309e5d6bc486ef54173761be822c8ba605d90b66830b7e30367b5350edee2fb5acf455fa235b99c4c328aeb99;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10d205e1401554413775b288e4b446addd6d8c3d770e2844dbebd613979a2d841d958bf12b4d25aebc41fc7869afe2922131afc210ca881b1b96da7c08e6bb8b0355f65b890e5e9aaeb4029b1d98d2adb9cb479aff2cfdae0a90bcdbe74673cf9dc6809cab4aa5776b4037855f7c8703b40ec049b96df0045;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h439062f7e6a01097116074287c1b35cac1adec79948be5ede68c4506a7d259d902b45bc5dd7337d6c262b8b84dae119d42251253f0489802eff843a1d167063727caa107ff4d4ac346d9bd477cfbca57c96d9cc324ef064b4b065905668715088a4670900f416baf60ea09ef86d87cc92a3005223856062e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h35ebb19205e7732dd1a9fd2f21508081eeb6a1168692647e452e454da08df7a0de538fe67d9564a2e40e8f9060040828e09307aa80a4b056cbd852792ef575e130464b20a4115717a2e49a8d00a66bedc75e4169e158c309b4bc9f6fab9e72fcc4168d342215f824d1016f46cae7e343b71733d43cb0f8c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc3aad787844578ea7e55faaf785bac46ff8c9b8a23a47cd3f0a9559b13825bd554bdda8d43ed0bf11d19170c86be8f94c9c5767b2f0146639bf6716dea0c9a2a3d995f9669ef8cc99175d1e352f7996318163a2715ad6dc8d78479c03b0d066bf4ddd00469a544a1d597e6c108cbfeaf4bf649af4ac19fc4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he187c61ca53c51c1a287994c8b0885f10c41d7ce68d4f370d202f4f02ece3d435c1779b030a9a3e24a444b034138e612ae824f04f4b19255e03f03dab0d62ef929b7a03e6324a09a74f9a276360fae3efdd151bb4faf6d3c9c66ef9e2da19a27626821675fafacdba7ba3ca99fb5ead72c4929dceaf82df4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17f3e98a94d585cd52fc54d9a2cbcb2143262e9c7b476db7af28a246dd7366036aed2fa9fed880ed9165af53e2a63d31ba7a5bcee7ed1aecd346306db9bd43f7d9813d263e5d32bb4402f3e797a8dc8f454612eb91d461632a61800d50aece9b01daac2a7373034f54dab75dde928e49a5c6059e0801ea02e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf78b317f0e712f967bf6b6774b0aadf40cd52f5028b051016541362c5c92dc931785bd9f4a7b3d26ccf556fc6ebed71eb3c51d676c86547415f5d57a6746e2d888754dbecfa13d5549c11e87f56fca2f7d4d0d4240861427135042251b7cc88876edf4bf367f11692972912cb5687e5ce7f4b2131f4dd03c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h100f9de512b4408a35758a21d333bef02f95b3e430168661d4607ca9461d6f49412fe1112e0cbda748b65b45fe7ed1243ea9c5096b5ed594d726de5518b911c1eb0e88bd6e09652fbc3fa8af64e54575c6f90b2550cfc457cd529845c6bcb2e3bf39d30f1e5e4e892277490fc5ccc5687ff567db8814c4247;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f792ff880558af30ffe67a3edf22954cecf94099a10c791819fc1c20440c828b09550f3a4956c71ff5504c6db4c3922bec76c6c84fd00c7016262b54133e7e91e53310919896f3d4ba3123b17728bf92ea63d3aabd84660b7c28f98a9d3d09ed5c8ff89e531cb1091349397eee7ec2805e10509bfa8963cf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11698e650857d142c2ca718b0a679e9cba6650975119b4acff1b98ffda7f3f50c4c067fa888fd98c208a5a35af1f153dc534bb581517e440e6cdd7d42e185e12f4b7d3a855a280b292875acada86e87cd00aaeaaf1182a59b9dfa98c2ba255335ab592e393b758b31a42041a1e6553cbfc785595ed61ae821;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18c80c8f12e7216b80c7c83eac51b4297145afbfd0b3f69f255df9a57c77d9b5a7110c5bfcd7c24788fac7a6edd67b25652960b5794fe768df4f197882d78a65dfcc707dc816bae425aad120a1097d0ad09cfc6a4be0530893fa18806a6750ec4e0bc26b19cd4457e77b787c80f1212c6cb87b7c81921ce5f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha3db1a16efd22f8cab08b154f607abeca805c29dcd46ad565fa110c1d605134f044f52a90fad2786710f36b3c3d0aa1113cce01bbfa1521b19b021bb858e3ab076a9167f0bfb654f97afbc3e0c6c35ed481e329eb1282997b7015d7c9fb107851ab63fadebb678df5bd2b04d6ba0c8daf99f026e8a1ccd7d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2a3e2c7b3d1caa7ae949b9ba96fdf012078eaf3aea944a82b4403657e3cd5f5dee73568d775ae68ed261e76412f3429448d795a62c1b80b9f7facdf6f8603aa10f7400bc6a4f45daf685e85253bb6ea70096ca0f20bb27c5e3bae33d79b5ba96962f3426562a9dc850f1791bfe38f271b8e514f8e07289de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hda1c90accd9bfefedb64a5401f401cdb41b8bfaecdcb9e93cf51f0f37c0477439169504b5915ffa67f9eee354e58f17e246b83b1b1e6f4a0b5dd6f2d5438d61c135c47c7781d9c30edd5818a9fdfcfbac24de53b902b88218c3553e5b436b612bc29496b9087f8c90713bbd93bec913a2abe64ffd8f6e00f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h140f253cadb6cae013d1f6adbc0dda90579351d01aaf5106729d35b90087a5f9066bcbac06a38bb391e00850d9be9554bbfcfc25f95ed5184ad21a0d4e626ffa20141cf5da4758d4c8986ea9b99482e6eb90f1273ee4f28d34ea0348dd3a5af477991a6cd494b9ee049992261ea162bc9cbdd0e9ba5cbee80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h156841aac4614669407efece37b893fd3a2e296a3d88eff9b0cedda33229da6497b582c418804b8247d25af8b0026aa40afb848d2393f377d841962d080bb3edef13680f5f27fa77381ec5750c89585ebdd3ef53aa9c741fd0fa53fc840e7d9134ff13307186fbf871bfc28ad3d4ae2f6587390a40291b0f0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha4564b15841ea4475f21aa130a0325d032f397e0a60000da89e5ff28e74716b1b9d313adb116f14745aa150d58a6aa2a35a5ecdb9490172393dd9f6722239a87f9c520b3ac231c1d7607046518048cd47eb21dce94820cb20858a86c3e32d302f214bc51283c2a3cf7c0c9379fa06274bd78c97ea94df4a4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h44bed0a07484f8a6ffb1f7b4aed73b8234ba394966b1daebdcfc223268b0c84f8b363433d5e3a33f4a1963d267f060f6dc7afe7bd649b8370470de1d48c9902a1bafb7547cf6556cddc529502aa4bcf23f50d6d4cf7a268cc89ae7c741612d2b696f949e4f07732d90bce91509994fb540a9b5fa718e6cb5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1958bb4149e1603652dd681c0347c92ed88e77bafc54689a257e3c4896e01f0c1f2500c6fc3dc48f04bd8ac78c50ec80ef7d666e350f770a0593c7ce33a7f1efd80ae6c270567a7606ae9e4853251cce3f7c31240e2c4c9f5892222af0ad969a66304dcb5746af8030a3512288011e856e7a69ef40bf033f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h39a6eb042c1e0404a94d4b8cea9b8b5ea268057c15fa8d513d3d861d30947d0aa3b3735263d5b663300aaca59b241469181b99da7982fdbc7c553f012138ecd69e79eea1091b2233d145a10886600cc75bdc64a947ec04cf6f51667224009d05199ed28fcc17283fddd9ecefab57e29add8f3caa3dc63a9b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h83da36391a16c78a5f841e8bdaef0ca3f5c48caa34590e00909f3ecb9874da8ae075c61dea096d744fea8d676a1e35d28875dbd849be94f95c3931cd53bfea30970b3b7c367cd5c267746c1e7ce610d98b7f58769cb7aa8675c98e85ee7d83e1dc6ea4684300c115bc908bc2eda4cd2961d88d70d29f92d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc2287909f6e8c1deac85f282d23cbf49b21b7b0006b0cd83f16425cdca850459f9b0d5c956f3be754aad43d8a5693abf541d8fc0341d1a637625a2267016e1344efdb680809c76145f8d7085f8321a9014bea59340b6127973fdd3bafc1929d688f6978ab642f108942b5872251b0aa89e5d113fe396c4aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a3d93a69f73914cc152ecac51797ffa3595484f2b0fd97cb7f25fbca70c02060381b16c644491fa07019fcf048b021d98170819898a89e85e02a0308e007dd5fddbeb36f7ad0c621221325ad445f9567c5f778adae39373c3e9851034d798e5716205ba52e13d9eaebc8fbd85f9e4b4d4652c6bf12f4f7d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcad5673231d466d76fd92b6aafd6dcf1bb6cd26bbfec4f443b297aaf61149bcde9ae554ff294b579f240e76457a654cd8a1c27e80e9eff403e7c31c751c62ba7b8c4a183e34ac105f812863a4c0767474d9642e39ac905bb45914a17373d5b3acc797bf5a5989cca7e014ce82b815a60bca7d78b8f9dcfd7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf92fb9d30429e2e412dc20e1cbddefb63db158d697fb043ba7299ecae722b0c5b9a6ef02db8e51c89de562577d514c4b6defeabd9cecb6dd5840e829c7d8662f9a9adbc457f4c9bef836626ad3f44100d6d948b035b3c17a51083051456e327434eed6e36d7dd3d5365cd4377a666c4b65e1f2f67aba00d4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cc432512415a1b01d83ead339f9d3503e0895363fcf547dba5904b618899d217b90fd9f36500e65abed6e99d26aa92cf78019f3fe5a6c4b2dc641806b18811d4b9ed74d9b6cec024b78b7d62e7026d3f76592d0b001d24a2bf89d7e02ccd1600c3de3e4e21abf1018ffd1a0c71cdcce27c1d9aff141a49b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7887cbf5d0f951d1b3900b0cb5c9caf8019324085e2e7ee70265daaabe4b933bffe295c9a0042a7b2fc19e554ad69306743ef8ec45363c3b97c41750b2c76d026d1e4d23bc3788109d176a6f4e808caae51d8c92b1834c9a4bc9db0a1c5c659b967a1449650cd37e75ac8d3b02a9878bfc44761a26b212df;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ddd13012ad9d6fedc0cd4cdd4e075d3d4f50b0d780025ad41e0442c4f36d84422a6059e5f69e599331784c7235776800642618e12863823f702e58096644ab924b935c38f116469579a2728c2d157209ec1e277a242ba6095a43e00addc14b26b5e4f4e7b119d0304c6fd643e5b0c912b4c7aaf2d97a6d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19af98d4b96b5bc3450996723d94c0e6b1fe3f26182ee8585a814e0cfc2c23d1d65563e68170c59061ac37caf2e46426f1284ea0836de4930f57a9485849c0928b44d45dd7e5af4dcdf78c86e25390b2f79462d94dbdbc913944dc04a5c5c991215b2dde11acb87fe92222649b7c7c25596385881bb534a7c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1241169ebd823d55bafebf69af0e05565aa638b944dbf0b0fd2e7ada264d181a7694417a9dcacf9c421e3335e0abebed361f4d844d36dfa5d932e9c8ee716b3567563d56cf10027bbf662e65a212254bc7f35410718754ec32b0cc937fe878a8849bec00f04f6d18d2a9159f27c206217076506c637e111f4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9b07d4a424b6e68d45d51cc629da5a15ba69fe35d890c0303cfde4df7017d87a79bbc33420ce00eb475845008e3701a65c72ff17503830a7a44200440f2ee532928d08e5e024e1ba2f78f2f3c4556b758f35948cfbd2759f6a0e5f064c96df020a2e325634f170c7f1984ab83f74918768547a3e606cad7f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7e609d1ed887fd9062367c2fceafedec996117d1ff97a2900e7405b747672320da9714031ef53b50ac57bb9928d4aaa27d7f06c209614bdf74f5ed66aec516c95ece4b704bff799c9056bfd26cf04cfb3c93d3e3165df0339009a73078f7904bbdb44aee977f7736f315aec1245922c7af4dce9d4d3ff6ea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f3a91133054c89bcb7e408cd48e1457c61ad449377959173d4b9f3209c088d058e386d457fd8b0d910e64e6cf9c776081e730cb05cc6bdeb213499f53b7eff01af7f6d2ec2c11f374caae836274a96d559a55e6682bb23588b4c1b03f627e535e2ecf8516f4c4c1edb93872a6f42c5144a73cbc339716c07;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e6b7fa8de6bd14dda04879f5dfbc0c230baa4e22d1c02b71e651cc9a451e47f954c03d0362b9f857b24b92336045f96809f28d6f064e02bf2a51d9e81dc14444ffeb98f8ad17c75cdfaefd2758db6919c2c1431c0a13d858eb5b5abf0c10db86715416f5a34c139bbfd3d9d11862eec70bb0e86271bd225b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fd161a2680e7b828b8e37ead9c5f46defade93fdf81018a297af2e2fa0e0a818454d0c6732cfec3d6eee7d5da46a22324d09d5c2df52a7e5f2a17446e06ffb0cfa68fe62ea585d2a4438e3f61438b270a6529baad8c9d1e0e779ced9b719592a923f4d7c8599808777a467fcfeeb5f35964d9f66c031d9b1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12e8d69f6d77fd3860c743f915c3b1a978c8632dea2f9037fee7c9f6a8e0a4c5596868915228944e2e674392e3782ef3b6c98f1ebe79062eee294e2a4efd39bb3a3827e52765d625a4e4c723048e4dac3077d9c8cc3940c920cb19f42f47aae0ae8b9c5b62fde8cb9096f30bc2e4a721620f212fc4d66a942;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h174bede7b322186f3e34b8bd9b16bcb3f1c017a72fad0d4ea54ed95de5e7b931add71d9571cb97890668a7a5d657c8cb9ce84da1c8829743661c0b9e65a73c547d780c138f2d4c92aa5e5e394e2248240f70b8dd340d4055ed1abd3527e3c5ef0ccbeb0dfe86085b9f545e9f6d7f1a2d9e9904288bc89d658;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16fe0c02f8c6762a9306a4cfccc3959af80d98c9024e1b46442ca240bd5afc21df73dd8e4c133ea0e36582530124650ebe39578742ec0d4118f5942959b8830d72883e06bf1009be3bdfa3d1561e693d3b3bb7084d8f149a931f7c7906258b8c5b2c34a759933be5572af2cfbd0934cc9a90025387e8936d9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9db50a22e34121ec5ec2c5dba4ee228a258b644ab8c3201b95f06b987c6c46f99bd5184253062adc437d9392c45050d3053e5cadb731aa580d30e1176541af4256f4dd5f38d491b9e5fcb5489a762ca092f94f721a0d4b29623f6ad1f65c5019df9060474c5d1ac94a9df89c5c7a049849186153afcd5528;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hed1db544950023beb038446c1a53bacb9d56760e2bffb27f785c232e152ae11d0e5e9659d0476e1e24b287fc9a789a9cf483a58880d43335280f6365acc3693f6a0818ef9e57d6dab625201d9f41ab5ef951809ec99b086ebaac2f1ac9973b2890662d5faf401e9d8d016b886ed5a148adc1cfa7e4080c9e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1190a8ce3b28f07ce4ce4f26776642f9f8abb7f427feddcdbfb8a8740fa2605dc75fe5c3cacf4a0902eba72a301956dbc7e5f835ebdacb5ef65166f2aba82ede93df6b0f71d2bb43c2857956e5a48f687fd494abcc2634b837a72d008f6f29f972a94a65baf5609e07cd96f3cc2c207a2b347eaa7c02f2024;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8ea9447f3f54198e3b6788e6877dc6596a0db1a07bdc74dea15d7efd579a2c8bf3b5e2cd638b99d1696ba57be5967f88106ee883e2e909c858bdc3ca590081c5c1b8aff5021ff42b89337da5b663cdd2da3b8f64b8c42137eb4329fbe6558145788353361d3a028c9bd1b1f72b91d9a8ce3795804e6bb0b8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he87d0248e6b45909d3e80a61fe2bb892d5205ebd6334619c4bcd1d9d48c9aa7a4ea66d5e3daa054c428756dfb95f1068f0fc98ee17c2f7495e1884131a3b5e08189f83474aa614ed44bc966b683f50f63f4da6be065e8bf2db3fa051ce32128a98ff7936fd55fed461f631d22ed82c3778b0433029b9d438;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17cc9429c1d5f6b5d1442eb085cd44e7dd2b086826d6cc0d39ca568fd28667cd380442ce48366e36a273a870164139843465ba17445c1425f603257976eb50e50fc0b7a53737f25b3f937de8ac5a5c2aba4fa0deb9c4a8ec467ff3c324ec99b56bf3b84c78b91f82cefe73d373caef23af312de89cbecc800;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb8a9a1ee0d137792836a925458f26aee99c7fde3578197c0856865d767efe921393e7e18d034375a119d99a24015a42b2f50a9ac7ee6d9a81bad24532b34e211e9887f9364f3b54ed371da3efd934f44760c08229e66a5b58cfb1746110a61516aeed10873c852088939de9845fe050def0436bc49e507da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h591e14c33c1f0ccb98569863f7090f9e173c83458211dce00e7b75955c847c833e1cee37a97e920dbe582cb19877f88792bb3d06b358b6245fa5d2ddeb0ff51d2ba6ef9d31970707edd7e75396ad60d923489a655f9af43ac9a41dfc3b6037725287267a65a97c917ea3e52124ab04e9becdbd76de7969ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c31ea9cd1cb5d355b00559430b65cb85fc57c7ec396960fd08ca240a7bb6fe51e522bc22cb6d7076dfffab667b2afa5c84e7e517637342a8712659e6ef584c462844816bfff9adcf508fd5957f40e7d5b5b8e4f63227af127125bb836a2971ebae32241ff474bec126e6dc6cac7f15aeef0d3cb364fc5ac9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1174793fb435666daa498f4cb1da9eb4056964ccbd20c986ba06a6528f340ab641ecd95e1fdad151325d9d7af10fc7e39af4ee7475fa00672570936440770c0e2fbe78b147ef40b4b506666e58de016646d663fb16981029ae10970aa3444fd0b1d93e64e9fc4137a67a771b6b8dbc0f7a4a17a966152dac5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b281a80da5ad15247ec977fbc74e8792e835bae2e757fafa6e9b0e78430c0672885e4c089e1135e0711dd186f0b4f62c19c3925b571d020a18807ee7bf3afa452b7ff136963aaf862eba5dd15fb1200a2dca26cd56ae743e0dd1249e267e6e34b9c5746e732213c182817769e9b32ad012235701c9831f08;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15adceda3ce63bcae15c214ee2b158f50a80d4af64544e1591c7d45582ff9ae954d3a219fff713a1550dffbab3b3c470e5f24c5cbdde88c3fca9905b8f2f62677e167f1a1c53e47d8b179ed0ca66e3b2437703e908b778b88a7d975b7dc1af4c5ea1eeaa92c6ba08dd2090f1b38120fdc47b9fa3ee5ac3225;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd20ff80aa6ac1ae4132cdcd64b5434addbaa8bd4f4350f2f5075cf02a254cd66d707da8cbb0af145ae2dcf9751acb9c6cd3317e88830e57b4ecfe5ae26cafa460fe933e8b96bf82d7b2fbcb096544d86db01d3679279115ddcd2eabc160fa4d44cabe0e3105f09791d2e205f994ed5e3d9566c3bcbee7691;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9f8b15498b46bc9f7f768bb323662aa1e409dcec7bbfbd13f69ce6e860a5c8a9d46d3ac2bafc5f5bf78cd688da19588cce332dbe040631d961d58ee2768d240deb079010800bd5d47e01e1b8ac6cb18bd1802626c025bcaeb27b2f58fb88be189e7a4d7da046cfb863309bc6775f999b142974145d3bbaf1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12d2d30f7131ef56a60d3f580272238f06ff4210d970f0e9532319dbc33399052174c743fea47caf723deaa18bb0c7315ca47ae778cfffcd02b3c33bf903a33d8ff7fa8db9568947afa5bf9a762800fbfbb6e4657597dc4521776445f5211cef1aeb16dc9369016af7a41f9c0d07c5e5d12cd31fa9c3219da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb502e76d4f14e54adaaa1151c1fc87141d716e2ecb6185a4befb0675d4a679dd722e6ba606e196c34c394d65565fa6ecd951f0ff7f8f8d7461774adb1423d6b7cbf62687593176f5b53952366c369b3169f2b8d79fd21deea0b378216794ef743a8b7d134bab97e7b787445482e64a21c5136255abfc9f10;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d0983de91c520a311046c7e489e7b13298316e492e0ee345ba3f9626b893056181cb310378a0cddb0bc0a7c2be28234fd2bb72b2227d7badea5963d70b25b51a9f0fa383382590ade97def537f2e3088710daa9e91a2ac1f8410b79fcfe2098e17549389eed63950ca1ba94c9e5825ba4ecd90d7363560e8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bff7d2ebc2e67fdc08449ca831c7da32de583bfc26558819f424c0f22218c750f39ad29bddfac3099362e3b8a9525170f530dc20bb8a5cefb66778ad08c9e53ddea5785f691ba734f70f10f40756096ba502443414f99223a36fd7cdb3e937ecd97fd10407a6397f910a4b7fcb5b9df89b01f66a5abbd2c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h913c2e5cd3db201434cd70fd2064a0e858bcfe39af7cc3c8b29c6818faa31b972ecb6ef01b4c6f8b96b9bfb9aeec6145e3e044553436e9e50250f1c16c0eaac51e70981355fc1ea38645fce2c98cba3353b33ec89f672dac65135af724673ca1b61b7e90129ec7a3f6a4944e5516e282a87126ea2d2c62b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10f185c6b409d617aee02c1da5b95dcc164c0a7c0bc7647735e3ee1693787ceeb0477124f93640eacd53b8f132d3c5852d41b627da308750ef384e3ac3883708774454470ed2013ddde99882a40017296a98e59cc8b7954a12acea7e101196498a980d323c0c6f4f91be2d4b2256f41e2fd3f90c1d658851c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12b9988c1c0fe99eb973bce3a7d9f6c8774bf82927ba0f0c3afa78b8c3dca8d7d55477f15c973865251a90207ca82370c555096de6faf56e76a0e171b1cff55c5ff59b5c949480d1027655500a5277397ac8e8a3abafeca99094779348237fa2d35720a68bea8a5bfe54b15583f525c63b9171d092fd3b878;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fdd7f127507bc16c43f9deb5945a7c02defb69e778526e41dc062373142ef846850db10f2237c51be6aa55d1a00e589e3e55b30be9cfa5b1a07c2e0e1ed1c6e7ab258639225a51a5882fd4e5d3adb2fbad5275aa497af66e14947f25ff5cb4624b47d75d860b7262bb31ead6cbf93f749bcaec2a4f2237b8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h121ebb650579f0d703b98d50763ddb1c808bb0e6c931c87dd84dd4fae8c6bc069eb45916fdcecdb5fe68ff70f0fea791ed77777d1dcad04139095abce36dc56819fe109a9414bd680e485600b1133583196e23018776e758327a094c67dfbd04e90cd16dd5eebde17490c7bebb476727672dafce5964e9b05;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ea01f498235853442085f21c2d825a0ba7cb3963dbe7b7af9106efac87e433ceaaac14beff6733d7c4ae691735c6f29509728c6e1fa5c928292d575d2101a4000ffc93f4d9db7d6271d135e2d81775eab94ca49b68c6956a8d0d82f10ad0086145607bf6b993e230b1fa0bcceaa7be25712b44250ff9e45e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h175938bf590524356dfdf62f02135d3fb51bf068e2eba9be20bce52d5f16fab2f642a3d00458e1467c67c325f1d08964d09793d2f57f29f853e5a0be0c78194302ae1ebf0fdfe5eaf672531330c2c2a07ac4e94239cb49469647d8efbe061fbd4e9eb7aa4d45860d89c059f99e7d94530fb2162777f1c6740;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15bfde4257268a1f85158fad82ffaddb0c6aceb45fbdd7f23e4bca768273b800dbf2bbb632fa036b678d7e516082c6218eaf07944d6fa7238043e7f5186c98d632e2babef1ccca544c243c88f6404f672016cb837522de59aea8d4f719a138f840db18ff275cdfbd50cfa8acf59db3efb6fefa2fe4a5ad0c7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc7c060a425ef67626cc48d27dd75ad432d0046c4348c63ef319db11a5baa9e785baabc85d33faef5edce3fb6849c79247be06b8c3e49d0ffe4b6ab88d6d7be0b1cecebb7a9f02e613dfd5987452e8db995ec5429a2e2e5ee0cf07e8b897ecc680af10c0414b7c01bc9b1652ee069ed0d99b9c4bf5bf9a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d0b4cb8b664763be166df6ecaaa1c9d38e747816a565b0ce96e1d0e7893553cc0eeab1984ba6327afb9beb4395fa1931d5c92516ad07f3b9e0b864c6e1330edc63503bf13541256371994c252e27ecac774b06f3b3c3ff80622dec99556098cbde6b7ea1917d2b2dd0cd978eaa586be113a6fcd980fdef4c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cda60d15bf250719abce6671cfac39ebe1603db39846a57eddb9f739a498d243e052c8e5122640fae42475a85e4a854a51c95226aea182ae07fef7b297edef513810a002db2280e9004099c554805c2c3b42d48a31abef831985fe404d4dcb60d84e2da7323258360f8f608ba4cfb9c25a27822e21ddc741;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17aadfff2e4d553b3d8b6fdfce3a7f77550f7adc999787ee65df8b24c1ac886f64f79f823a4d7ccd4bbb984760e77856ffddb11ed8afffa4a09698ea65783a77b28bf4afc802c6aa9740d3c97d8bd9e0215d0838b6b7b644dfb07a320ea1726483e02746be41b0a0ed5a1cc0fad4f089762731d2445c2298d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1348bc73dbd6d28b27d9bdba45e77eaf8d0df1c6089b6df86e82629169b83134a3f39735f6a1317ec043a9cd9ab43dcbb8529896d633e45583f2a2087974b2dd14f33e5d954de07758d681f075ad2c2e3cde649e97c57e1ae0e83eca6e9ce7811eef345ee47e07d5119a93f7bfb3f7c032bfba2f458363055;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1960be690151bcd91c17f13aeab38e482b2d5afafd92c5df65f6bd44261bf58306abf0635b457abbeb37ac009ae59724d5e0b1e0aeb9bcc53b47ec3e4dc5a13a0f95b0039df9ed395f2ed9252af0dfb7760ee821e98849b9b681f366ea522834772bd25a30a94836b3b5b83818dee2f884fbad5111a2d02d9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h449e1d5f672d59662588362ff5cfaeffda48e674f6278d0cf208e6cb447e5bc2c41f7f7caf984b87e0ddda674bcd99af907890afdbc5d419e192312ccf9a6606759d6a92078443a487ae5aa4e808007dfce74892ff136939065692259663fe25b728b92cb7a5d825104e8764013309527e0b710076a7ef58;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h123543a25ca4ae5c776dbff74394c382e3ce3867b21b20ed123422aaa110ff9e33de17f8f10cae1bf9474cdfaaf9167e50330083761dc639e33a035f1008915844f0c0d2b1810fb65d7ffc2b8ee03d61cbe29e3cbb3ab4851464f0e9e49876d744d1a91fd7131b21c768336bd44c5ec7456f04e78cc618377;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h105e7dc69903a06caaadfd04b6608887583c7098e2a836b33ec0c85de15411205b3ddfee7cce3fd4d0d613f093f17585ea11d0111d3364cd25f36b1a64021e127d4656c65aac60137791175ebaf486cb1a848031e92b2e307034bafed08379ff9a332130f92768f2e340c31a4dc1aa7674b0828f4e60ce43e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h81b18df09f09bd66a36e86a6ece1bbd434dd6952fc75e11203dfa8c0274f60b118fda2ac2c1e57717beb334ef8c4d60d1f7b9a4ab1fb13a8291c15e7cdadc66ff81df61bcae90a1c0409c4309cf54ff9937a8380500d5b9339f944efe676f2446861ff8c280ce24e6dcf3f9825257241af69aa25f0014a23;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13b2cfc08002dc6bc2b3e8067e78476d31e3f20bf6eede421c9bac0794e034cb73a1284a88c35d9c3cf21188febb031b866820c6a6475209cc04ab1300112f91c1f10afb74027088cbd3267d4397a019a80ccae4d0f04d802cfb5d3ee38eb653e5f302c05e4023a377d5e10895acdb2ca1a4a1e527fda6ff4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7a25870df5be60e950debf7d291147dd7de06da2cbac1753acfdd7b38e89e94085ff1971120139d4d7a05f22c8b13e9f89c87821278652e126bfb3c2f8da42df7860b91682553a30fa88eba5cd738c858206feca5fed5c02d042f9609ca70152739046a2fbe274b95642359962d7675b092de36be15d1e74;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e2e01addc54ebdde04e31c587fd54ae0d60abf44deec96d73dece0a6ce1261a817807efeb4e4053d5862f0aef12c670886bda75762e5eff5a32af5955aa5048488f80f4c73816dc31ae61ad3e4de4b3e659293c9e8950f3372e7644e6a71e23d823ab4ecd2f7773daeff464abbee49bc73485bd83c63c522;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f4d99e22fb94f4c5b78068fe75c42a1ad2cee600fe1a3c19fe26473a00742d32bd285374b0bca7a1bdc53fc9ff11822d85f10622d1b1e1c356585ee22dc77598eae38a345f54eddcde242c589da2eefe5e7ea26a024af1c4962927646027f9f41360092efb24bc6c4bf80cac5cd0e97b90554f8c761c019c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e442d5acc95accfe26f45ba2644a2cf78316f09cc137dc2e5b6c62e57af6e2a2c5b97bd8877afa28df79ebb0280e3ed0f3eafc73cde861287afe4c946c4187596f8f66bfae0e903fdaf102560ffdcde0076f16bdfbe5a12e66b184e821a0a582322419c95db768356b8268e93620c62ddd5da7150db52057;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h193e398e2cbd9bc4fb4330b623ee86efd89ccc6fdc4ce2af18be47e3489bf5c59eab5947443db537624900bb189ec7dd56c42500ea6d9c387bb57bbec9a1034b60e93cb4bf0ceebf4adc65cccfa69b8067d991a29e343419c3d21400396d8dd3e93425b4a67f02bbfc60eae6f650cfa35fa4a97b8c15c7d45;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h787a011cb048ba9f03bdec396839192ea8983abf5fff2e2f32c247583422c2bd63d7c032eee256c87783efef6da5e45dbebba58b97ab20bceba7827e2d7ef2be8f0a8071160331406b4be3c7573c3c9e13a033ae3a3bbe82b38906b0a1062d833bf6cc404e149a5e8b5b9fe6f9c32ae1ececdbf9cd056ccd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1822f1f9d44c6e7b571ac65df94d297fa83008b0b316878612d519f26f4655d2d5a24050f69b58c47ad3bbad9a6525d74deae8d7fb25f9b2fa5dad8748cecaac58b4d6b59a9e0edfa446bb2b673b8c4e3e633c5efe5e61967bd1a8b36e1fc9eba454b5b54a308e432cc37a394542b742aaa3f11b795849580;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6bd10d5a874f424b57f7aaea794f6b05c9e259abfa5514e61fdac02ad9f79e9b52b98c1ef43faff189c53ef1b0bfebdf5ac71de457f51ccbd04dea830f9c18faf9e2fae58f2b953a14c3870f009122208bf186857cae6bffacafcc9ad806a6c47e688f46514201dbedb921dacc6666c9ec60e27f8e3177d0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h138e9d679273eb7cce22b3a85c7a3c9fcee49fdd2498c6191d852a95f7ffc32520febccce8a99f847b55e86d3fda5b76ad033e567f4d47fd8ffc4ad90d9e3129c39a5bb7f6c1d238cfcf888c8389608204e336e4a99d60da50cf4c8e278ab67b8adff62f54ba2be109e117adea692ba4beff2ef424a8e4951;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19e549a8dfef5ac454fd3645532f5b48d7d962cc3dea16fd5f07dc8da82ea63a44ba06156064333100f7a32d30b64d7aa0e283a53e0fc4e0040922b7285bf0f7d3575974b61d3d99c41e649944436a46da184e6f30dd26ed31c1d304354648717aee4db14236b155dabafb74d8ea29b7abb64e32fc0186cc3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8a938faebd438e6fae405e5093e85111445a1a2ed9ea1ea255aeebc3ffed73c5a41b66f66e30e4a9d60200794939708a75b84b795998100576e9c029ee3d50c186e5d72d672b13edf8519622763ea50e29c1da3fbd235ce641a89ee4be782c2f49af801791e1e655b6ea3ef778f3cdb45506eb3c7d1feaeb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e4ed2b70e19459a4e2bfbfe12be275269b7f7167756f9fd922122543a2b44e41771afbd22e53ce5b68bccf506e501feec90b8fe2c068283803bec56b6e15ede0bcb1c2555367d0bd6d2935b92740797938ced44762b96edf0dadf57adc912e82513f77f59955119935dc5448748e268d91ca27056add95b5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19abbed40211f7097e8e073fe0581230b9eaaee0a4c2d3ee519e2a0604e796264098dc25774688db3af2d35d4c838275915058c3fe6e68d99723219829ceb613ce38f32968c53c87ac453817cd30eca93d94eac97fb3d822ae0c589ec30f7edcd907e81b83e585afb1c1a275fe070979ece8157757bed4d85;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1226f9fd3c132a0044791a141ee376d0a7e67d02cb780cb4cb711226e5761b76c346943d424ee7d3a03094e07d5a76fbfa0ec122c7fd73991457a4f3d065a902e3d905698e24f08c8a543a14dcbc7ea69df32f142a53924a26e2485068ecfcbccd70fa145f434ec7dbe364536b47b322753f58d6e6c42a3b2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h147f0737a522c68341bd9acd19393e8ac93a7251c261832a449596bd36ceccaeb9be34a24a0a9b58ec5fe1a8e47eb6d66c46c04e6bb7059a806fcdcf5ae15dc8e9d7bbaeef481ed7a03372dffd16fbcd64c28737469cd7b11e484d5e9b3e3926dd4bd6c0102311bd754dd7c3979936329752f3afef3e723c6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1db362d359f02332ed8a3e8a40b1a3a7eba9215c8d0cb09200e97a7a9351ec801bb38c11bd15c359ca7c407aec62f8d2700e5f089d919f03f0f0f28f066b2bfc33a2978d45e14e8ee991453664622364e7ded4b61121ea00248429e1aa923b53d07ec8cbe895757a1f582b087725d5858bce08424ef0c0acc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h85f89fccdc6aa0b559b1bc5947d0ad37ef2a8ddc82e3a6fd8c8a7ceef8b9e1e03f5ff9165c8a3d3bdf06038111ed2c8750954c11394aeb910ef008ac90d8b5a577f7da9d3fd06a35b93140072ecabadbfa66062b1002803c9071eef361a99c0b4e141e33e6a84ca55917752e6a1b808941ef5af0ef539ef8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10bf369b6ae3f709bc5875af6fe421c98fd0ec15632ae822e8282cea9c815d1a31f19d9e189943a4818689306014d92406c2579812892533518997528f7e9e95031db1e84dc2a40723428be8146141be5ca8f051a9635b58699fe10404ed25836221266f857073f77b66a4d66d38633b1233f571e124787ff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h446f757e7ede607c1a63cb9f13e9c65e13790cfc482415c81552f5f476f1fc5d4d24d03124bf1354bc3380f46fed1ecdd9bed500982814afec9f4a410ec25a833206a0c76a4b60f0c0b185487ee2c36fe461291f03015e59f1b20e6069298ad21f93259273f2efd068ed035b32dc4c05926a0a9af1455d02;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdc021565eb1c3bbf67815bf2601e38b95de2348b3cc981bbe3ff2d8fe783f681c040c9995f56547921e34744421d092a4be24cd4f8da08c13ee6424eeac498ff3d7168236d2c212cbc2aa21e0bd82e4a105c233a692b5be4499d30b167581c5eed17542316f5e70422269c8219f12c480ad3a40d824ef72d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1027aa16c9205325b379b8a3e1314465e0dfe1d01ba4cb56f0aa4cad10d8b9a205ac1246c80e13be98e739cf11d133a8c0fab70a4f3c7194f332f5da189fc1e1569da26742ae02b8ceaad4554495c874f5410fa3a30d36f2743f71a802dfd6cdc533df4778d1fe2d12d92ba33ea1c6f796fb70b47198564a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c5c810599299a6863b1004bc176fc9d46e839ad59de31824c4ae13af5e28fb5200b34db30b760b6eec6c539735ec01ff76d789ec8f905ee0a8f1877b5bd464fb43d7f90b2b6db3b45cc437569abf0d4ea9624fd0ca45701d97500a7a9c036baf52007b5819a942472a06563d990e09b28a469c5f4ec39a71;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hccd1364f2449a6beb3e04088f5d2e084cf3abef2f002269d2df1bd7a5e6b0e93e68d142c4a5c23c2329443d990e9b81bd30322109dcee6153c688181c97bf575a6172de0e61beebafcc5eec7ab83d07d9a7569fac247f91702794b70138907227f29425578a57c2e2cf95ce46cc879b7c55e070e2359f680;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13eda77ae24e8743ea434243bbf4ee7bdccc646daef3b7d70f987ab4601007c6d368da9ca22d152b95da592155e08b6ebf2f6b815632e2dbd07090d652fccb22915b571b3ecdadbc336373642cc562be6911bddb94865a8c0a220d1ee10b11ca3c661e8d3e322f226c1311ee6d63e93fb21f1a770a61db2db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1285b7d7b6230a72402620633b598b2a8ee8e3f8ef9382233443e2e8cdd9fecb2e92fe828b39939bbacd2b7c941230a53e9e3c43c87997cf012a6921b54a4a795e07ec00f334660683f5957d0f01b2eb2cae52aef7a46f2990d433c86877780b8d54b4d99312e5e565ad7b97f6649b9597980bad515e2663b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15c3267a7d6955e7c0743fcc5e94013ac2702d63e81b5e7bb06764cca0e1bbefeafaefa2e3c6a796e63414a19c1f0d2ac287397f0c12fbdac0f4f2653903468132a67b5554319c62e2a3c8bfd37868bd736479124a9af39285062e71280e031324ab036057bcbce9c5da41f084de7c497132d091a9e62654f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h114ec1d0ba50b69135ca07a271a7a0ccc2772d274c843467f21a7d52fb2c09ace6883afef34be5b962f2a5b54cf5327db65ffe47c176611458ec23cc752725f840d4064e3bfa258bf0a759ba481c875ee4f9bfb484204465f99accc49415b2f24cf41356e78b5c535c728247f23caa56d0a38081ad050edc9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2e4a45f9f2cd3b794503af12bf7909d1a0ec1cf4beebfc8b61c7498c5c89e38f62e1d3321cfc1a80812b39919b97c5be3778b30995a09654eb1c18262157046da6fa10e1a97eef4660d033a0365acee15b6bddb13c0fd0c5d9d83701ff9aea27d04832931b1e7beb41da0be2a30ec6a433e594881a1fef75;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h59be9548f0d5d0a9fb12a73e5c40d335cc3b4e0d356869719afa850de1afc0ecbc3990ee6cc177393aa53f42834d93453dde7725e87a323c66ce768620828296f40ecf2499fde604afe44a8705371d82670c87461dc91d35dfa04ce6285c485b9c84010ae6aeb4f06b671ada8302f4c3f9083e3c25a66c19;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha4d45c26106302a8af513360359db48edf7261c37e2ff8fd2416b71e72b7184536467a4c37c4b04a5a850150214baeb90a18ee1128742bee1ca389451203e8eeab3de4bf8f226101b89df1fa92ab9040bcd95b0a3f1f563a23852b7a7d6a0e45dcbb995da6dc6fd8f76080f174c2070deedbdd36d09714d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17edbc1dc643a2482e1495bc227a6b51f0e2418e557ed1b8db4c17985f3b45603050919cf3df0a62ac2e217a9e27da4d49c8dad01199fbd9dd6f095a3de31dfdb62132e57bee0cae5589ade5dd9d7d6b9d8eec7fc78e2e8b583a18f529017f41ee446e2107e779d2a903f384e167fd4e8125cb7936aae8069;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1952a2ca069dac7446ea4ae9ce6757e87356b3d160b75b4ccb5e8922846efe768acb7972f3b7f191fb16a1e6000ab0fc08112974f4b614caf2f3aee0cab15ee4aeb57a6448eb0a3548ff9d50388c633e21c5c67ea5d87102649974958bbe12f7f93cb4cc7c83f90467c5d81c1bb45b791c3bd3a3fe6419985;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbd522df3f039a7094adaa8a8d5b478d4a4ac48a6b89bf5fcacab3c78608e37c96837196e54990e21522d1558242a785894f9dfb4c63e4b1bddd82c1e0e79289c2fc1e171eb1d02e70a26649a8ec9eba9b6048124158db55c6f604d36168a11917eeb78efa51ebcfa5d99fbb5e0570f907c1482adb9a24a14;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5c3218800e0c4e0a095d497b0c18816c980924d4316a8254bc48f792051b92034fa3db5bf27dce726900ba877dd9b7a19578ff4792dd1ef35c910b13f8511eccb9485f42be3762250d91751e7c6f45494540dcc309a2c7ed8455b8185253aa7d6db6d45020e99de1b08c224d89c76c5938ec02b905547568;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f6e52f1ac9f17dcab75a9792fe179501cd91c22642c37ada0d967193353e78accf49d1e92f26b483067a6ff3d8c65f70a4abb0ad9e41a0c844bc447e74583ff29ca13e3e11da66edfe4f1074e5190f95599ff8697e83d92608acbb197ba2ec01417429251d05d322fa8764211728da05f9aef79959c95be;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e3b25c9b98513f55ed4400da7c21ab93a3fd9486259d7790e35b300c25254cbbbfeec532833638eb9ab427d4e70acc49861997cd12c9555b9239b633e953b53da46f7389ac82917a427d0d0bb7895c53b8d554f9382d0de4840986e7669c451d2d67cd6615681b7f4d82706238308c35836f3fa45adc2131;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h23b714ab14a10c5c9e3b545f11e74c01f24625166f6811402b1e06f11441fa340833b63fc7270f0ab90560d4531eb6adae781301530d8e45d22f64a11c7a14704fa96cabd4d4405e6d56c2758dec356005cbf3e682e41d69927a0b327ad7e5cfade2bbec306d2db5637489036d972b631b6b95873f3d865d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d159465e5f75505c710677e49e57d0da1491370f97b65f7b7e17e4530a7486ec4e6e8e199ab5c4d0194d1fa32278ceb9acdf6a4bb0751ea5b1c626e026c54c671e34a744c8f0255cb93ebb1340bdb137e03b331ce19bc080376036b5051cc02aa486b1e4e187cbf583be542753a0a1d96949d4d621cf449;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a42506590d0f034266c82c10073427643b4e3249e16ba66237df42d518bd6604a7912200f8eeb168c89af621855dce0d5fe44700204653012c26c448ae61f8ed67a787e82c8e8e0536b21356a65e3ea29562839ae94e1ce5d4aafce3329134edefc3a1cf81e0437a0e196a45500988496ff6d09a71646ebc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a1b53eb1764c39a92f6d0b9fa98ad86e8200a897d8530f0d1c6e9f35893d085cd53076f50a7c62b56b35944df5542f0cd96335a4c1c95f176926667be0e9c83c36a2b5020d7c5c80415382cd00e08633ed8cbdbb8aa94d0e9b3b721de4775a3f7414a9fc7f4bcc8ffc3665c43fcdc6503fd1d73583b3adf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fa1eab36536ef504190ee5e9ace451ffa3beb64929bfda2ee436329823d76062f85ec07817cae483b3a3c9929789b3de660a3b5f4e4660c71496a6b3af8f08f9b1fd8d8ce5dcb59ab0144bf1badf9b4927e432a0987cf24193ac241fb335bf8f63fd64400d362ee1c6161ad20d937167a0ac675ea228ff32;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc0a173825f720355b8c0ddebe44be4f84cb2eca05f8947437122c6ed91c6ab9b6470e4eca98c6d60e2a891ccc5fcccab67a9382c1991bdd3ce39f244ee2e077c5fd951df84ee58eb6fcc12c0db6665d725562491f564a6787f910a909316cc988bfc4801783d0500e5f40db7fb54eb609f1a3b6ff62d2f99;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc91f9e98172b4ff6627480dba2d4ca61ed9846f169259a1105f83c95dd0e99f2cc4d2ae717d076e50dcf51747417799f2c46d164334b6a917cb256b495bd7e7dd4f01412739795d5c49e4870e952050b943b73a03d60e0fa0a8cada47442c42408a331eed491ac20eca7b9a93ccb19a7699d480e36e65ebb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7637d64796db4867fb8eacb0e41a1b52d9632913630e8d41b46b073d89805005d2859d029a74ceff80799b9aef2978ef3e01cbb129f58f4404893b75cb69b8691efcc8325055e4dc6f93e51a88e8da361864ee814ddbda2dc8bc470d1f3664bb9d8ded7d64c3896cf9a9ec7e9de6b5cf5005d120a209dcab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h168e957d5750205b2d7541be6e266044068539a92a9e4b7c6da34611bd762a8329f12da32f7c63a1819bd30368124226898ee4112c5755761cddfd78ace70a646a8d7d20b9737b0a1e818a34bd1fbac91a4c457f5a89decbc5ef45621ad15a878ee970833c159977f0b8ea89f5ba727030a3a30ca700cd701;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h114ff3ec829d6ab7cce2c66a4c98a249015f7addba3e26ec68e3a52a7fa051bd96a494763463c9add2b2f146f806d305b23286283c97bfd9c0fcde3a874a00e0735e6d2b6784d353f44d38676d4256803cda7590bf577f7b7dfc031532e74345f3b2a10ec0573153a5424d5f396f0b019ff2efae437e57ecf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e2cd1fcfed5d03b8754452ec89c9884a83f87683a323e7171f8ecb102120a355c95308bcb3db805c13578009d2c7c09a9e6a219d2305354f732268acd54e9128e54a74c186496209e868da34d0235dfd04b863dab8765639446e26dcc195d9d64a050a105002465688d824f83cf27304772e85078bbd6ae2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19b3fa2cf2fb7730f72d26f04c0653f634eba3d488e2400b7ae6c3ea9b4b164d5d01259d3cc4de7aed661dbf6283da8edfccd00b49fb6d36905f190bf1c2593f241fddc3eb15849d376403f33473ccb07a9b30be80d0c6ab3f132fe463f9e8a263599c69f28b18122e6cc90e011a0f59ee3d67bbd4bf084a1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17b773f905259bf729fef2f7dbe1626e61d86e1f848e839bda9611ba6adc2a69428705891cd4e8143cda7b6cd50f71608376af312a294ab7f9de405a5608049ff25e32593c5e96ac2d0b1f2091b59ff0a35d7d2876f2678d34dcf7e2d780c8696754a507cba7fe3b15af04b244cf15be541dbd8a8bca4f2f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h899a792165c4b82182db92565acaf29a3171f47eadd49bee2a44307d1be968d833e2b5b6289a3458e003454a92fa9d63540765ff329f13061d3ae958696d96f926fd71f0ddba55401bcc3054d7a9e53a91777127283d9514307912a64bc200cfebba585ebbcd49079745b17485acf4c92a4712e3792b2bc5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cc33b640bcffc314e41139c287b3c76a1df39808e83328aa1ae1a2aa63b2c5032acb394e0caa9249c374f99b1a5ac6da76c933f57a4d4f2ce7f99ad13b1aa8441ccad285eebf1ce1bfa5d6d853dfeb1c64c2c0392b193e91a1589931c8b0427c62eca670a9e4d57bb20539f08727cf4a1361e0d5d61051ec;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f74dfb750d4fe2e520b26467fb6eb32f83ad0395397ab22dab1d057f6c20403c3b6d4ed9ca4e0a93512e2a5d3db290e941c5161da12e92ec5205191c3603fc47fd474a201854ff19453069007dc5cb7c4ac00d268726851aa07a66b2567cac99598d50aaa744f83e9dbb9992fdff8d5c7832516df7efa04a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1224231c18dbfd86f065055cb03d91d5548664ef1bc7ff3d66a5e1a4fae75e67963466921d8c34935d5d14d4b64cca47e888708e3f031fc29ca7d8b05728be747a3a737b5a72d7064f7cfe697b9d285cf097d2369db807dde36d1cfc130aac0abbdbe20baf1890e3606b21f5c51a0ff98d773191e1009ce67;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h113f2f41f69f36d890de9e18d730536c683ac0e7e624d1e25cc4be1bf62328efe8f77d5c3f656f90fa91e74c96cdb8690b481f945b418544212b1e09158b5d66b00ffdc257ec36c1f8049a7f6aee85c31ea094db439a2e35b2c333af5f67b298ebbb1ad66525c891a336b16f3ece242050930f90bcd3968a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc8b4627905512af8874a0e5c180a31d8cddb83f3aed1d7068d4079ddafaab3690229d5032a154bf4296dbfd7dfefb4648e6badf13a70612dd85877cd7f914e66b6dd12b6959591033d294565d2d6187207ae7a9df81a9248616b4fa5dce6aa88600fcbb9d867a14f5cd0f5daeb136e1096c6e0e8f4dea077;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10f364c459553ea0ba06064b4a03034c8920b852068ec545709371220cfb5787f24a29f73d832298f8006283e93bbddd54714d8ee593e52e69102b8217a64edfa9228338360d0cf1905bc0d9cd09d415711b45ff5adae0ca486c5bc3b1ae3faf839661ceb2ff65be7bf42b2f6b08d7ae977ed167854f2c145;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16f7b396461d739fb575aa5918829b943d5b05a7fd44fe02530aace152f39ac07bb58a155bfc94aaf8f9e884b0917cea24f6da1717d53c2417f1483f68d30b51c8155d8d6fffe52e7b478919fbdcdcd6bbb3746c669f17e6cfd6bf8f1494d74eb533e3b70ee6a1a14eaa26327858f2517bcbb91d2cae019b2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hac63e7b0c8d1f90cdb5d1a6e289d347bc0e8faede5f53139b996dab67a6277b9a4805a046ada41ba05cbd202c037e2719bf6177fc26dd7899afedbd7f01f44534a2c95b3cdbd097d1d2f727150cca1ed1a6819e214d2f34b2bcac878e7080e37e58723217e4ca265dcf5467445bac1b2b7fe3dad5303ba4b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b41943b7ad49863ee534eb39e29dc44614a969044af0f55c3e7102ca78de44e682f8562984dbd3f2fd6bca272a3deba9b535ac0f8ca5bdb1fc0d4a7297b07e62b244931b39e47e26b266a1385db7eba8aa7fb971d9bfaa79235f2e6c746e0acc230ff2f62048826a9e805f78ab934826d72fc0aa1d7828dd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h669666d774379d4dcdaab8263e15a435ce3cac54d2373baae9f92c0d1c03dfc0983f4a007609f12583ee2d9bcc4894fd7b353bc54c94adcad4f1843158e23eebebd07a78d51355ce050e7075b2daae90e8a917d7b1827444e710db1586b8f4f60016e2d0add7df69349224fd06f3b88799fbd3e6f1674add;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17aa0bf1ceadeea9569e1aed45e8c002bb38a2bdeb73d675954e68dd3732c42ac9d908ea9621d3f517718b59bea75297e7184a406ef7a7a1317b1c77f9fe4eac77a2b6bd1e64a12e30de937dc5ce56031281aedcef9674c95de00ec75bc7392c905988980fafbeffc69811b920ec1d8bfa4891d4d565a9189;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c473d04b23d0bcbf201ffba7fae3cc3c392227ace2f59c2daccdc24ac04de0f66d366e152065cbd6ee239f378c5b31ee05f6a2d82e521255d2b3c9b9a50abe6da082a3061c1724318d3f2932b28c90d6b4fce1501dfb5fb41f0eded13053347b03a2fa478bfadf0a703ee227864a3b518e26e16e9e173bfc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7a55f8d0f88acff2c15e452c125beb1d0b70dc0f9e2977be348effcb7fa02c643b0a497dbe70f03c6a9ebf960bbdcab0eac9e5a0389b892645e958e852fcfab49c0373cea8f48310b1ca30586b1190a33a8d070912efd92e7825571b7b7e2ed507920cd417323612958140187986426eab189af55bdb7b70;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16e9539192255820dbd051553b54f1a170ed7b4f3ec170c8e6f1394774c5133f7958a103e0389036283097890b6dd51713518e2ef0b136132a232a03585ed8f143bbd6bb7ddda840dbe3fc7d56afdacd2f56b9f2bff5502ab3ff5e40eb1ce4a05719a5d9024191a829c592986b52459ae5a87334e2a3ca5d5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h125bd933c84ff8478d3acd5cf8e06c0be8055a8cef3c6785e3d6fc1dda928aab880f1ac4bfbf1b8ce56aa361457dcbe12e477717eadeda5fc56d31a527115e06b48d391f4147210df0b2ef0dfc57c27d5cb604ba25b3cd241ca687f154e55e7269452993ca0b6c4c88728d326aa560ed9a9acd22594c7185d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h193774b25c334df2d64274755ff8ed66b3d21c7d3aca36541f9da14d1cdcf0cefc54147ac58ef279a339e834a8def0062e9920c823fcfd34fff1b41660a28c35872f184ae9df106eec65037b42d3f71d506ee6daf0d8747469782307555ad7609bc4d3aaa099d1baf87df18d9a5976a1e0344f1cc135605a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h78314be101de30d6e19d516ab92ac8fb3c770ba3c2003f00106c3628d946fb247436fb3ffe8ea2dfbb9ab6929e1d2b9342a147a51cb9bdf15d741dd3ead686bc9dd853f87a59c0537e6eb79a228bcae177b91083b78cd5d9b068f4c9efdc7e8de28e77bf431a3355ea7c299921e9a3cdb140d2b65ec3fde6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a4aa3b9fef0eb60940b8e11007977d005c150a9dfcfbf9ea60bd61ca090fb8a5284fc29662aecaefad0518a025922b01f5c3c23d00abc9dcbb0e7cbfa155466be67ab6ee4a16e51a6a5c9e84d44750a03e9c34b4662be7f3e43eb60f81d454b40d16856ef7242bde10dcdadaefde9fb691ebcf3b0da696b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15fb1f23da132e69acac02b86fb672fad64ccb3d2db504cec17d96da8cf5fdcc013c0c96ba7a5e235736aed3cf5e7d3072b8a425e7aa71d22f5a193dfbdc76998dccb4bbaa06ca007369fb845c4b20ac42d50e270dbb5c133abbc477c69562cf6ee7bc1157451a109de2ea145adb9d75e0fe34c059aecd584;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h26edfc3c97ac88946c033d3197923b4597cadb8ffa799ff2c0130c4f09946fd0811eaccdadb05cee2f8f150242d5465e71a004d62424b9b65536b24895811e4edcd3b766738d49f0699185a38e9ed7fe3a03f4df4050009679489351aacd74caf17e6d22ee29fff043a435be9ce06e0de29e7e69b211cf0b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h190f9f0e185582a1c3b4479e50d706bd40e238c317332f6cb450f5bbb4c8ce563ad917315034568a037860988d8476ae8fd83f02aa76c4490621e3ae6c6a9e520e32a68574d7a57b937b81f680d85468cbc3f6aa048e000336c269981960c52ef241ab98092a39a8dd2731d3a15a0f2f4c33b05886df522a6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h976615b80efa81cfc4dd9e076b0322be8a7c9ffdc4f839a33b063dca4c20707c8abf64d24291bcb696955a27a0f48f3345fba45830a912e40e712a1b92f5715bc6e89f51e4c95ebdac13aa8b3d64edc10426e7e95310755544ecba8065ee7e6d5edb224828b84b1cdd7888152d7de902df66d8a8e68390da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h99d7055c426977ed4d64a7881fb20a59f31ef9b5be35403f6b3182d6b977edf86d719896fe1c0e6a6a76c1114bd650402109dbdcce243b63d6f6c62bc82164b1f11e8a555cfff05d3200c20ae9f3789eff9da920456c9f504592eb556e8174339532ee3abfcef885ca86cd5f81547e2386ee1d68a2af28d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h580cf44f739199709f1fb7d0f5df56c9d2b2061f29af94119ddbb43159cdddf56377dec699839db381de7b76d072f6fd8c9c1f6c828b35efdea9581bb048147eba1e799cdb98b90d4767d6063bbf8522139359b7638d1a9f51bd8500705558ea0bac3f04e6cfb4a64c3ec2ad5518ed2ddfca09887a0b0bc3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h482555f215ed38ecfd6e9bdae24020ce430f1ef0eea5301d078cf4c6a3e2c60cc545688fa876bcb31b4f24126702020221ad2ae59d6ab50bb0a9e8f215afaa8c5fe588619c36162e89d2d8121948142291867460c5ed570e62a520a37adf24b8d036da1cf54e38df3b10c1efe9624fcd7566795485a5d399;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h411c502880792a5b075f0f848b678e0dc9b536447353dc7d63df76daa69caf5fddb688f574375cef5c327bd3d4b3bfdfce9c4424838f70bfd52147c6dca0eb504295fc5fcdc48573e3971028e368b93c4fc0d95a9d4217ac7b9d8574f1405d960b2207499e99ff1a0e0311c84a263f0b2d9edfb69f7b3e0d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he1ada8699ddfe230940834c88042bce3b63a8582ed8388856727b0febe0d12df7ec9e726c8d4574b18037bd2ba1c5d36f3ba2c768b06d5801acc86504e7b87c0b177a7c7c9f200b65d213162d6505adf048442c612e9cdc626b7fb236655614fb5a09f70a98e0f7a7db485ae571b057f02e4af573e4f36dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h168e0dec2c18af6fdda2fb162110c0f9e485049a480fdf31add3e7eb95b35c5f7a8d9dae8e6e39780491ef8782bc6f5089f4a29e5ea296c075b906dbe876b6046ee275fc62ddbaa0c14741405ee1f03da538c7e570067c9e572bd2dd860cf4b4db0e467a54f3bdc0542a6cf00772b00df113ad267b8fc016d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1da7fbd5d30bf638cb67b7834177f4f506a1450f6d0a89cf3a62340ff0d1301e870883541d38f2557067d4656b4f2563b4619775a0c03944deb7ba7e0e70a2d39e96dae4645b335bc97c74ad040295918b7757a6132aac9412d655f94404399ff07f646a0fc4847f9b0a6e8223b98b75cc24fab0c9ed1cd5a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146c0a11ec3febaeb5798230e08eee17805d9d7dea08020ac9d9b2fca3872ba7b5dec935b30faa17ab36d9243af9fc2ede150fe8ec81e1a469d451a63f1949d2ce812ff4c63e6e1b13f0c58c21a399477fd4951343c51277ef98c8d6809edd41178204c02a09cd3a953be921eb00b344a4c40c7bc4403bc8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcfbefa1c9afeee7919117f27edf37a8d953485622612223a966d2a0cfb7d05c6f8e7e888945c2217a3d1bb2a3c167082aec2af47f10d37076e6d0928f344f046189b63c82fb127d28e9602b1cc1a3c32a40ceaaf355cb0fbdf97a9f051d7f256d14d2987b8575340b3febdb3fe801853b303560627ac38;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6cba5a961048569c41eae2d3b59e78d9b9496fd02560d3d11b5befe2bdc2b3f7ebefcc6974254c4bb15bbf12647ffc33b6914cadd970bb62f30738870b8d1bbc3ee38351a05a5ceb2f87530d147d36ac85df033553867251f832b2ddb4f77ae819827e54af856b3b75f4dc91aefdf70ed61f06d80b15dadf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13570d081eb541a091d92ec92e661d42f914929baabe335a616df38a2f30f5fe439f2242ea14f8bf4688315314ba2d0dc0abcfb8e6a5ea6dab93483626b18b6aa7c0c56686db4593ccde747f50d2ff3926efd5aba34ec21c39c214c4f0756ffb1ddba8d22fc60e0f8a4ffbc2b193280ace37e6b3d189f4fef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f1a7415baa6512836446f25551c8a0470d0bb4a5f8d5e0ac6d37f809422f150a92dc89f82cd13db273f45551fe69e4d488d60f6669e7d932da7e201c65ad281c869b20c0387ea20164ed640bf59ff90d6080440e3672e01d848cbb2d52f314d0117e541d3ba70a4f9d673dc31e418b74612af61b77343a56;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc86591f225d7a69439b511475c6fa8387e2ca6646ae1b3b86d73c348a63a7b17ba349c8884b98740e98f3b307bbe6660b789272b4945ef9eeb2ef8539b21ba6eaad38f6d80a74438ef7e4c0226682f8b749caec15446cf51614bae8c17b5a7117526008867fd873d162117e670b88b2885f94317d830e4bb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he469ec0c989616be90ce48761b9f2382c9f86e106482e851598489488426d23f7c0e12b0dbd80a4eeb7710b17e28744b608344479d5811bcdf5cd3260d64526f90b1283c387108c9f4410eabe3151c95be1334c48ddffaa1ab55ebb468a65c0a8699ddcaa5adb5eb45eb2c9617cfd7d4c125d4bfe4e913a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h67b5931ba2337e29ede3428b2e2eeebd22da0084a8314b8f93d3b68312dc1e392f9a5cd6efc234bb9ad8cdb513e594656a39b407da139e4ec624d2b138c94817146739637edb810c64550640ba0b57787f488102a7f00008982bd61c5e4c9ce13119455a0c89e33d86f1a385bf74438b0a98fbb560a96a7a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a126b3efaf356260759e4fb5a52ce95f5edfb1d31820be1d953385da7ecfc42703d10e09cd247f776bcad5354e7c8d982bb6c204847e9a59c79c08e8faa3a7c85aba269c61629300604f9a8ee50c67916be609fbf3cc04f5410b005a20a79dbe4ec50d067a2172641e277ceaf3bbf51c1e333a569cea6be7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1553c034c1688b387f6574bc02fa1d3253200a92c2f57e6124a663020137991c416b3dc0f20e501c116d205c1ca3eccdbaa6699a0dadc34be31afcde13c4eb61c8e4e8b4d95e9ac845598ffc2a8a1d9573a8a73839f365bd5527f121a01964a6106ab6b7ce942542a2180b6c0d17c1429b77d400f7d18880e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h268c90ee677dfcfb7882890cec5881f8967140131d60c4ba16557af86ba38ed427745551438bd4dbe0805a47a7aea2acc0e2afc972dbb2039ec6a35cc5377eecb469da665e6f77ffe1ad97d3c5ee310ddd55e865467118e4301c8f14cee8927acc51db3c4294421f52d87474c0952da45b0e14ad5422f49b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h476f6e6a2a1ebb5472f0ba32c8eb9760c9628230a204de7d6ad1fc23320140309a794140e037dd8402e44f2e3a0676d0fff3d603743c1cfe6e28b07ded3e41df43f8633f4eab40636f5268246ab7ce879687a965a50deafb1de9043bbea780be314b253d138da1c22600cee205b9f19230c290248beec0f2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h162a9acb2cceb560a34c65214425e7032792df664619b2b58c8d26e1e7c8b20b4d90d09ff6dbef061ddc9d987572f4243b08d470feb22d210a815637112426f129a7dfb71c70910eddd1a3b0ecfa5e4990dd12dbea3a8e7b01a5f67329205cea2b023d5319293da3cde852384aec5fd2e10324a43b1e92f4b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2096f4927862d8703f4ec308cd7bb91fa58d7171b9233ab3a1f53898fdd448fce09a390104909e41e434967d7e5974757699d9976a03636bfda5105f409195dcda29c2d2a6b5ce06a2d05a9021c0711954690b28ecc1bb0b4d8681103630e6b9102a66c2d8bc51a6d7d3feab659efd77519b197ba2fc843f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h212fd73fbd224c37886579bd26839a209ce0c1ad0d7c0a25a0623a9c2741f2de52c6bf361e443b7fdd4bf03a1fb8bd027c15182a7a35569ad9b1d9dc68d51f8c33a3a85c7d7b3adaeffcc03b711a8395b76ed84008c1d595e1a78fecb51b11f166bb71ba19639f8a9eae394e40da1aab2ece703238f0d6a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6e066b0d38a57ee18393391aa320ddc2dcaa65534a6f0f93325cdd7a5232874d22bd9611bf3ef9a8ef5c53f67e2be1ae41849972a752047e746702e2e727b34b5be311e78b947c38fc9a1f81990e39c1203a5d0045cf9549e3deda8130806a4f59dfa741e864a35948abb3b0343924dc827537a660d7222a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hea0f9899a6918cdd4f5560f82e43d975900e3b0552251409a87e6978c4d92f8c5cca374456e534c9303a923e6d988ec50a825b5793af3695b290514bb3ab60cfe94e9c44478ae832fc4b320678b26f17b67a6df6a262d5b2952d1bee0d2160b79ef01a9f728d46a630cec9e197702ecb1984b22acbd9f73a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1876db0128ed3009fb56ee5afb91e2df2e6f1ca9eac1aadc3891e95d47a4bced0034c32205118636b0ae6a5805a864dfd6fbf09d6912b5ccfbf7b3a854471426da222317715743b7eab6084acf931abb214c776476a9d24ac92219235cc8a1e3f16eeda88ce13c5d37c8b463c529f8763be88cbf8948a1cb1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19cc18c1dd78e62b6cd8b7f4af6cbb8ff1e8b2b025a72fa677a89af164f69a444f5e8ff3c01698ae21e62305b1f65e2bfe91abe9e3daa26c2276421b22ccf0c611eb2edfa83442835d5a743562dade3203f9782edbfde71a812335446b259f34908b681190aed07de6a790a35ee3a48a1076b6c931d5f3ef2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h106e5ccdd84161983e0fc5accea3c216fd04031e525b61c708a3d15c1e2ded692352041e556cff70ab9ad186802c074181828ce0772ad4eb8944f42c2e5e587b0e56b7f5d27369127e88d0f3f0bcb970d2d89726a829e523bfdb5bfd2727737ed8b5fecb7d5fe0e5a720f047c11ba59fcdae0348e8e48bc0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7550d738ba95ba1eb6df0a0755d05e2c67745bde101b02172f8423472a0eca9c1de5944b160c145f508d9dce2742c65d6c77c4050c41b91994ff0d20c904e44f194f23ed6b2ac32541d58b7ab2cbc4097d7975ea9cad92bc6e6196bf1cff0c60050a4582341228b9ad40a888bab356bcc6f479161e8f5985;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'had933c5f21d1f2e9d88a4ebd5791fa5008f62e0b7befbfc9b9ed7b55af809c544b28c316af7e875fa5c7ca8dbaabcd70358ff9602fc533782cf7efc5a3cf142cbbce40c4b91ec9325a9bc0e1a6e5b49bcd1b02e47e76246c52419889dd470d628b639c538a5918d134920c0702e949356029dbbef3195c0b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hceed9cdd9f34a04fb9038861108623a1a7b5e0fd9d9acb4956d4fc1d44d9c99f34d076946f31f6fb76aa44439a1fe31b5a754f7c882e9c4ee31464d60ac672cc89c8416791c05c8d1c3d7b7e610cae904fe5258a60ae23cbb955dcd438947c51a0b93e92ab2838cbb47ed8c09efa7b019746b75df57fdd2a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h54ca4c4ba37e9afc12d54f3f157d31edcc0a516e2839c6c7ebc09c2041740a6ae1e8db45cef1d2eb1e77db862e12ec4b1db7d236cb71f4af18910bd33a0c3b7a92b5e59e5a526b3c8795dc9bc5bcb0d522d2aad712eee2d1c3f082fc7d270e7d088b34714bd1502a257005962405c66424bc750c8478260;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfa563b319e7d48f9b2d412b640255afe43b058f626d1dbe80b9ed6a0150f897af1d96306541222b9ae6a94b1e28351584cbda251dc7f59d946dc6400c1f9d87faf74d00f53a59ddd8ecd21605a275206fef70e5735f37950d717e0c817fd0ca4e3a8070ef4c8ebf842803091ae7427a9135956da8a2c482b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf7a948575fa6df5e9ca1e7f6773c9a7fa6e2956ecd04febe55d9f1895d62375a1c73eb1e437bac7680010186affe44f2cf42275467058f0a0839999c6f082e308f1b76103bf5f0cf787edff0a2770ef810bdcd4a594dce1e374cc18a54e382f818539b530eda6d000c866fd5268fa4dbeed72ab9b4de8cef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1550ad60b99f0d704e93ad8fe5495a34badbc63be801d37b9d560b83de4b056f0dc36a1c899744876592006ce30b25951c095e77ada2eaa8b626cd290b12f6b228740c8e7581e13603f55e9a59f1287ff1213812dad3f8d99b65ae2a23ae67fc8f808e4c24f29c508eb26f0f251435eacd133e66636a20c01;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1efdcc8956051d78981a1b01369c21981db2d1587f6f8ddb1315c9be68445d6d2889564af103e285089cef3709b1182d8ce839342cdd9db99d4b4065f51c338274cce7eb648a64d457bca42c9fffcb93016afd35d5228ee61f6d7aadc4b8db3c6ebe0908cc4158811efdd1bbef246cc8238ced7a708432e1b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b4a6eac14ca3ffd2127e33f456eafe03a039b3f35462673c0ce798ce6014d977a64e4977390af57e00f8e52f3b39fcd9d68e4d29fdd7d8dbd182c0a20b67d5ebc5f65de807dd01fc0b7cf7fd2051889033ae9376b8615fc79a0bdd87c6c0b6185aa8b632c5149c4a94da2f6673185c1b4145db8640c96560;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h192b44b00b5e8a06ca5539be00287e59c74fdc5ca1b3c185890d102b737e597210795a8a4c55e3df5bb30c0e53665d2a7748948243970d8a5afa8f09aa843c3ee9e09b3d3bad083bd8d74a97001162ea14d3bf27ad85e37688c0acdc9d888028571101eabd8c93a126288d8dcb1a098ad862ff58c00862d49;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h68d69b1b573049025d0d1591691ce37cb6d9287d9835dc45217f47d5302baa51ffd7bc6d9cfe6606c6d90f7bddbb8da6c2b9ae502a3f65ef22ccbce8fbb5c992e5a9be15831474913724a6ac842117280a4260d561c2223e9f7ff86f134d468e71e1c4b670551ee7ad228b7eac3f15017f23ec00fcf9661;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a95b2131287fc58e573914bb94bd2a7b866b21d9e6266070af6716a267ee912a99d167479aad8fbef4746722eff34b27d7318e3a6fca969818872d532e5642583bfc44bc8c347d075d2439e2d1c2a25b39355eb2feb59079acc8275866fc8b03de653e899b2669cf2f745a024d3aab2448dab7c057bc4c55;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4e2078d7b344db1d7c5b3f3e08524e1872541196e52810bfce3e339828789e56cc29bb829b4c1ea7ac14ff68ef29070dafe460c8a99b68625387989a25e3a2cccfb62b4ff9624d39007d640ec46ea5d14889e7ec351117aa6adb42c60c7efc04b4a44e78d8e46971488673ca72dd0dbca2dea34ec89696da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb1bf2c9b14ce3fe282483165cc89bccfa7117c1fb6b902331c6d2afe68a3f0ced808a692671c2d9fac724de551cf8b46d31dc93f59bd5a36f0b37a7ab1a139c60569e9e13d32b5258f8e1515f628095e84ce05e1d6af82fc07c0b371995b85dcae731b11ecd6cbad9a7bb6a2374628c87d99ffd6fea31885;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcd892a2648f3cc5b52636d4b763e7d706a0806b1b0f683986e039945f09e4281321f7131cd4d12420ef0e82008a85a03621e2180e3c0716a7b0e44b4724e27f541574571239a42e9fb428a8c082d59faa8b8a2332af729d8c7f68af29da5a725389d1ee2a223f90847445ba8ed66b6a143c24015197a7f23;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h984224f6d64efd3ddc4ac4e988fa7c639cf3de12d9f50f9b95b47d009afe2aa996836e568bde72e442596ced1ebae8cebaaccf0713b7ab431a1d45a510118ab73c2bc7e5eb7aca9fdc4cae3d5ec3fe79df14a8cdfefa5b34c3d9ae09b98a8e809ac38ecbcb2da35caaa933d39a2ae85866e7192aba34e5d2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hae203448b663f000772230884d229caef3bbc3342cf4ca320b321b94ddc42bcae593c22e61c9686d7279b1bc689804122791ba56a34f16e0ffbf9e1fd81ffb78ec807f03446d63d662755ce23dd4a994a1db310776726353ff025903790a8d04c15ded6f6b09b79a49a9f9e55ea0741e5ccfb2b9c0209b47;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha166da275dc5cbe49aa59c4360866620679171cc8898e6d31bd7b3e22465a4450f128faa40c1e6688299c90624d920653df70db56943c52425bef54b2a0c634cf1b11128fe4054c451994581544df7cc01ab7dfd42fbdb0b02a2dff35bef67bf0fedc03612ee52f84f35948f701c8838275018e9c9f2d8a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1752b39d0f8379f35aa676fa870e5eeb3f41e40bb787295f175b6ced2350442dcf0135dcda084f4f0dfa5f081505b0ecbfc719717d89358c17aaef61cb5eae3df461d47b3ed801df8f8bddf95cfcb58fa24491b388c9837f41a7e14d46e30a547a98950ffd82c67f41620efa4a972f9d237d819b1d9056620;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h492a088db2deb6b2f331b6d34b3e38f3a1df8b6e8082020c1b67026fadeed95b267f1312ffd828a488c51065aaf5a311cf26308bb89c137476a253609dc31934a6a9a4bfc245ca389fafff3f7ef28929079ef506f1c83a5323034b6ec5c25f315c90e801a117966189ae336e8a732856aaf0751329131f84;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b91a0ee4c1ed35a1787c15c12aa862b208f0ada2379aac9e6e002b0398e7232a774907d6c0422c09414873cd7cc90a29b78aaaf9cb43e8ec789841779533fee5e0e9fce17549b40d4f6068888fe9a68469e8c4099e81574f810e91f7ff77ca78ccffec9b1e8de67b16a16b171fb91408dc9bdd0dd9abe063;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b99acd6f3e0adc1753d00b337a5b6667de34f51ca18e9888a0954177a5793436848c163d94bd8e3d494c6880d6491f7e7169ed0d8b6f0b296b5c38a94510043e1f8b44dd3fe7152edebcfee1dea0342ef5a224df7840db7ba2507aee5eacb35e4f1d6d4dd0a17e6bd3be5c4e937eeeca28e4d0907225c3db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h763c1530db6a9511e430a6ec669684b05d7b9ea9d4625ad6374ff23aa62d996242791579704eeb2eb4636ce9e8a2f00b4e64ad4071b7fa5c256b0c49743bef36f3992377f9579d4be959908572b5b1e2c55dbfe385a3ce09a1a49594bfd00733e66e064a1296f19022884221b70a8b038c02959a059318b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c2d03f45e0c5f4afe00d6a0937a2ace0b95ca02267314e169a8819c879a8b1fb2a5480ff2840e121bf316d96288adb5aef6b127bb917478a28b1181f2b7066b352bd3be695e69c30602eec0001271bada66ceabaa2e29c833b5fd04b68dc3733f9db24b98af746bd88f4e66faf7b0f6ee6e55f1ed4baf76f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15cd0cbc36928ee38702aff4d38988b48f89ec713deef3c1e9d4c58e9e9f29006943fe2fb914ea3cc30f2284ae176bb91b2172eb6575836cb7429409c21d8cf0e6c298c1be28099bf3036cc6386e40fa263f88c7c3aeecdf371aab2dfd953eeff4c346f834eb866579738b6abc07c7ae9cba43e78e0d3f0ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbc41c6b0d7feca92ca709c94e6075d220554f9afcf47e616db9043e030ac57e8b47d54e2cce51746194798cd06a100743af29a6c150d5c14448c2e64a5ed477f17f5c7035936053e2850e2aab4d360a56e00a13e4a605f5ce759477962a2f3c96720aa642a2b6ff6ede44c0f392e4dfe3ba92c1c6214b25;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2d520c7a17ba7e20f8bdfced52f95db9089991aa6fb1e2cfd4401da35244ecfa022b62baa7b1e71d651c662b88bb243e130315bbb624f11d39f7054d0e23137693c9d171d5bd2a2f5b5521de44a245119a8f322e9b9d89a190edabe275df12e7db6438e4146bce9a4fd18c80db0bd2042c1e84fda11d5a20;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf3210e19966723af799c226553620b94aea196f9e2073c30fb714498a804dd1da45cccfd84893192620b21a664b4d6df808a1708428936b82c75122c8ccb66cd83bd9b81c422f4a60d9913af5a5219b3baf981dbfb11a5def40c8bf7033ba970f7dab1b30919bf0be94f5d0c66ece1bbdc40c374898b2d2e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha55146b35b3381361614394135745fd317efe13b585346c421432c8452537f998142edaf2d402538d277f72216705e798151c8b4ed5d1169fb8aaafd1bf1a056a203744d00ffb12a5734562ff1decc997f3e1d40ffd0deb73ffb7687cd6020e3b843f8973296a451fc9a24ec5c1ab280d8a294b98332e482;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bcde70ad4b79bdaef1bc046512d86cc6a9c4fb1834fab3b24ad6ef5575cdee556951fb8cf84e42da6106617a527251f159952af088bdf7019ee275edbfdd165f09abc364a476d497ce70b7147958475ae7b203a3e57ab7d036186211b2aebb0ee423722dcca10667957cd3811a970e84af9cae3f8957263e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14fd573d99bfe49b2195a6817c23253531ce28fa6fdd6a5758c02ece67df39cecc2f83295d6e1d0e50199a651a96e27465c0f28b4969338df875b4f4192d61e064f35bd5fceb6f929faf419dd18aa6f20191b6d6888b45958c9c0c667225d99568884f6fd40e03269cf9a1290c5e11cea6b20a0949a6f8e81;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hef39b6c99c750c62d24875eef8bf7f789f7026fdc38ae9f22011d20b54e542d6bd51199be7054a1ca707c7921291dfe88281d4bc185aa28ebac6687cc637f1447384db48b6af2ef2b2766fb979eb359b7efa3210936682497d92b0757097e5f71895d22cf2c9ba4a0a4943384525ebdfa9d773a3cde860d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf2e891f26c7e3cd4d2a506fde6a92b23e7706e5ba21a3186559876d460f8d42b0de749fb814b0100bde2485812698e45dfd1e806f93ec9904a23e39a4f9433a149e573bf80fde85a1e23f2274a1633502337e46e509dff440a967ded3e5b86c73d98afd7f8acc1dfba6b81494e448117b92318a6e4c9f13a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8cfb81c598be6ce4c2e128ee0d540d3c3d66b9c01710052f21f2383cd99922c6017894a50ec04945959d6271b8513543d107c07d11d25bb6d20aecda4bcbbd606b9ea5e8b3e1e4666cf73ab47d041434cd69e0c0e0421c13b4d02859a24da81aa43656ed4faac8ac76a136b0c27bf6793aae2d95d6597cf7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16d34ff8e0f163770c62fd7b10b9ef416b495b325f6845e3d8ba76a7873599628a4762333c6eae229017f769184fdec047d5ffe9da7899439a254120e3c350cabb39aa5fd00ddd89f74ed79b9e42683ea3d369774b14531468bbcc03804a6da15d2ab4989c7493448b557d0adb4e66fbf8eba30c7906634a8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdedbb3607c2629ffed66a43601a43c8418c2ebf5226e8b8311e34b1d719a068d2980419029d5d0bb445ab00ac6386d7f565352929535712ebbd2b417a5208b5f34eb7ca29ec31911c44f605610c33fe0a67acd8014a04cedd8c9816eac0a2d5ffd5eec045bca292fad8f8b8b3c2209384fa9bc6a7cd2fe41;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1272b2d12e05c7baca3e31b0407a8428effb8adc29004aaaf4d478365389325131904c87c5c3183163a811c177a103e913157a2c240c2f6be9d031254867686082960ed570bf467ae64554f7efbb05b25a7695df617152ce8db94e03b7c1fcac19a12b81f79ade8c4fdd407949d93456282137acbaf25bed;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16141770c861eefb9b14428876532331e9113fdc3dc3fb2dab7b7eb28c7cc5c72bf1cc3730cdc822bdcd3a5b8708e8251738432a395921a5f5745afa70f195c5fe24aa9d129ec5b40d2a796f3bd1a48efe4ea4957b25f5d93a1e17e2d24a48042788984eeae64891a2e3eae0c6b5718cea8a64d32e190ca26;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13e17c6d6f86031e3dcc7b892e8ba3e62b7c0b94b5bc5352db917492ff9496732fe42b03a2395c1b9d1f0f6333dd58d831c9168a0ef6b57f52c59b671a8c79fe5b54bcd3d36f3268cfc6e9d75ab80b3c2ac04f5a49ac3996e922da39c631079cc64b1af000dbbe1b923300a0fba56bb7b38e2964f523d4b51;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bf8be4994ae4266212f39e568eeb54dc59706a2ebc1cc24aae90dfb795ea83de452c5b26f1dd49fcee9a8f11a68407babadb514be65df0b107dd4c418a08c5ad46ba1dfd25ba97567a79385ca0de12135aca4ae788cf6147ce04191219cfc4eb9fa304a43ce806e60b14f194116abb2e6a57ddf1a8d82e24;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f758bbb182d6410da05b5b5971b024812a7f7dcc6ef47fcd5f7e815743e676a865f6adec16df9f15fd0e39a3653845344d7e93be9e2516f515ee830af87db6b9cb8accbd8023257d6c4acebf4885de5e261cf5c422300f5257654dedc73c328d9d493c5327d655fd2b04d190dcb39181ff05bd6d219d4f5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h877f88ddca79963c21305af3b1a8e547f8be357e18a4c0893d078e4fb8d9b3398f2634d91a2277a287e49495607f8961c09a491e5ef12f9880aa7f986a3bb0460d428a283652076efa6f7b17d292c16c29b6b543088180f03759f8c6ca036c7920bcf8eb5b6306f8f70024b497f64a320cfa0b03a412c2d1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haa2f9856df12d5d3012fd8d9776b26918bc7e4a93ee3fc64c5bbffd139325ecfe2c49b98877bd5c283b8a373e0e3f5c5c696a79600e422922d390c319a3d525952323dd763989fb238bb02e010d407ea0a84a4e1db78ee82290747ca6dfc5bd73fe75a461ffc5f9c4233254262831b666d183482e7d7cc25;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h314da39ee4c5bd27036a76954dd1d8c0ab6f9707167ddcf4cab95445ea4b435ca6a6e521efbef43900faf53274f8eb015ff2466e486e84eeec202a1a4ff0f03c950426c09e54bc3bffeb1ca37610c8e3b4ea60638143a772a3b33e50bbc1a1e71913910d30b60014a9ab433634c91ba0d009b925de3ce751;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1969da37c038d9e88a1201a7d8719a17680ffccfade5333e5c750a1ea6d02618463cf2f65f1e99af90ed6ae6dee33aefbf7a94c6565fd8eac1aec6fcc4ec76ee0aa5b45aa1dcb0899705e5e5b7e6fdc1149b0a58c16999b3f1b88f6663b9a20e147b25777640e4d595444762c07ac3b16d8ba0a2386b43c72;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h188244385f1bad55a1700eb520cbbc928dd7e1e6dbbbadf7c059e58d85fa2f5543059cf6a158d22430da1cf1b31444e3aa87ce1ca87de476f1406b19830dcd9ba803d42efa602473946d33542f8ef4b8479fdfc8e8f2a4fca3cc8e9e172da8d83b46caf5882af51daa45f36f10cf29132936458ecefcf6e78;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h179b2a4d48d252519c6f98e6bf016080da0abaa170b896e0d083bb5fd304c151779b4c85a781a0d5d9e71bb0fe2833fdfbe34aa340601bf603d929336f931f48062ca5cc283b070d2746f2f3d2408f7eed890ad6942125ba34c98ed130c81e8fdcaa85e9b11cdfd3755acd8c9883b096f5cdfd7dd7292e4b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3754fdac5dc2e8019e28863062b998f5a58086a3cdf37d18c9703ccd5fff435b03583f5f0da21b782a75b76fc7d31000173d74061baf050c7bfd1884e1dbfb26433d1d929b512ee143fa4f8f81a8c47456093afebf2ea57c36a89105a74d5b50bd5170eb0d4fbf3c9ca9e7550df27daeec4a4037577caabf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h546c078be028a30b1f22e7681eb9e560a9e8b2e67d73da39d1d784da35f57b946f334a9c8fbfb7b4fd395ddadb2293878558906a3b41b437e7f73608201521c78a3c41b55625473f44f6f84951b7359b248d84b04e045fad05096ebf987113f6d2f49e5b9a266483b041a50f0c2ac1e3bd682b08851c10;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b5387bdbfba8809b6a53f920c9ae39987244d44055cb1d6a1457f2734cfa71fa17ac3c9af1c0c96783707cf3297387d8cb70b65ce580bc9ca45d3ac0f69f8eb175210d80099ca6a0f5def29167b9cd20c8a8fdb7b72e5a8f4f5fef72082cbb098ba7f9124536406fa850698f38079d0159dc892ee57350a9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14ddb05ccd74881a6ca5dbca871cf6930e6d7988ffa8809420e504840b2c041b208cf59767f601ac8b849254b75a1e31ac126efe38585332c39b95283a5fe7c2be4a8258b14f664db80862524200d31d1691e2dc69bf56c1aba2b04b800b93c9fb94861e1eba059c2eddd6cf1969f48386d5e63542ec2ef3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1580a0fb60e126649f648dafa5051ce29a167a898ea3f622eb7435066bc1af1eb89019b1f2b150a71ad5f1508d5fd5e6ace8af4e9059f472e1f9a2278140cf647f7e6831d48abf876437e603a87825410da8df6ba77f3a08574000220499aaa4816d1f8dbfbcc66fead4cca3dd919082691f7f3c8eb310ce2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h172bfda84b83b0ee42f8be67e70457ce250711d1fe83d479a9e52253bd48050eca3c1da976cc7986cfb0208c796ec3cfaf7cff5d1730a0ded8ec4d52ae4d0f5f99fb117806bed35625a96edd246d4a4b4fd6b52c70a44e8b1f6130ef16fec564689027c332d90a4767c454fd5a08ba5e2735ff8b58c3408be;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a483a08421b6dca81faffc69f60af070b2b98502644d0e0df6699698ef2586721f7329be54a52fb371bcb177b819fe9ad6d0b0b6ffb176b9dd9b50a89293c3f9672245f5773e19af2108d187b9b69c2e8f72a5296be5e4b093a234e512d305816e3d9fea8c6071f76a22936fdd86dc6f46187a599fd31e6b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h426e1f0e058c326f470c1f88d838c4110759ad5f5d828dd31420607c931d146211946d752fa34eb205c6d624257cea2ae2e8d955b23bc89937f91ec49850d1e2d759f6ee0c6c050ab36f18279f96a32b38e8e97081bc25d3d56c65bf8bed4dbfe2741bc9662e9f8f493c274821b14cc4c5ad9140b3bbdb22;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1638ceccbafad178e5f0ee1b13259b3712fcd13d453a54310c972ccc09412c87418092242bd1fe80e5d0409ca8eff46f42c83369e6dfe271502c3eee431f25e98c577f2ac99c0b874d8b522eade5d81730180c8af1e6823aed3f826aa402df5219dcd9920b748a54ab1a1564d8eb23489f3d989ba645edd15;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f67fee631fdc00cb5402c26a192b44840da939a736ab25cb586779aee1b2d097fa2e323ef7c57855f0927a6a9c55592968dea995db609e01141f3c982168ddf8494f738830301d6f538ac0b9487475c22f8815d3b9188bf7ea1403c815e06b57a15964ec34d1e8b3e2118cc2319a6d5221f071ee1b2631d7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a5040348e6be0fedb55bdc28cf73c31f8de82629e1aa886371680cb0d837f0ac775fcc0eecf74a3078edf2ff23fbf0a9cc917de6c6285ccd522e3d9a569883c686d90d426c7a19d3873b157d228ca4ea509550b68d87f33a49d596123a7d24c7708aec0b001389a521cf684759ae98b441390e0b3203f21d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h140cf609cb4e7cdc96d1a025da7f1c147087835cd23e57847ef2e58666f3272c3e9a1b46a5d2a4913c06b62c319717f5ef2ecda801b1d41334389a91f92b43d1eafbd8949e284865638217da6e50a47030b2d17c6daa56cbfafccd3f4eebe467e1d48168c3e8ca860b8628db3e3573bf56c0c54063657d0ff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e4026a59fff944aba5e4eb8245b1bfa77a168465819f5caaf36f25134fdf7d322fecda232e4eaa60cd586b4a75b71ada152314a7d017e9116f2c62163c401eecbde3088f76676da852201aaf3ab3ab6b59e1725b486e7099fbdfe0e9f50c1a70c68bc0fb19cd5f40d0dc522854efabcbb7112eea8fd3cb61;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12db32d57dc42122dbd9e9472423f3278bf43623e9de2f47735154c537fe8584c92271576d32fad77e1992cc5d67fa54bfb548e1327cf28c4fe82c9d5f8ec77e4f5947113b208a1cec8dead0f168ed94d7bff582c7c7146a55c3f90f02c647e1acaaf6fbd122a60d647d62e9f5491ef9aace954c82f5c9239;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haa749fb9d7acda272a135735831ba3c132f6553510b6e4658490c642dfa148b4637b3a427b4d9d41464556f5c122e61d0856f5bedd06929bcf1145b62448058f67185ba43ec010cb001d0a18fe5df58b3137f9386a9f08b98c3e628ff33afdac91e665397fd64debc0de510f666792cb6fa0886e1ba28858;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd0365f443236a083f2937be29167404d3f8fc431ddbb0f81f5465eb534a4553cb5b2f59e3e71dff4f0d957444ef778dd43ef16713060aff79fb78172bda28698344b391714f3eed89ee9707bbaa61c9ced428861f64144ba19728848db3d841b6eca77442cd7c7f7f5b94930d3053630e2d55e79002cfa94;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h180b6f1b77819cfb512b38193ea12882a7d83f7afb003983d55eec4a199294891e3bb3a33c00969bba28e4e02184174c6c5b2e909830b7f2411a9d27b40cfee7e7d59dfe755745dc13f6db6627a44e776cd55ef4cfc6fde57805982e49e4a9083ca9685039c493d5da5260658442b0ed6bcc6e0247992aa25;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2c85d070f019db91cc2c06eca1faaea5a24efa693699b47a89d17af84873a8fda438d4623f3543179d189e130290a9160e89ca4285d5cf4f70a52342a9fb43dbfa1a47c5eb575c41db6c23b6a964c2997d1709bb61472823e8224eb59110a733dec2141def0841dacbc405fa4b07dff70e4f2fdc812ba914;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h506421f0428cbd033494a638f6cbdeaf733202570c4f4c6d5eb846e945ab78f595cf54eba0f313fd15e5b5111223f98e9666c5b6408d5fe655229731f1d8fe852f54d33810eaa2aaff9ce06a71fca6bee1af7a0e2ca06d146ca4c70d2c4876784f95fba5684d8ee84943487e919f4de083d6c61670075561;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1435f52eee89c21e1957194ed42bf5a3c219a4356c5e4036a5d081db066bb6f1037e6089947214c6a7bd2ba51cb5a50b6498b823151eca26f30593273b43970c0b5195f9831e79222866ae9a99b3703d8f5ed94271647aad013eb90e20ceaac5f7f8c5dce3ac61822523e2b70d92568704a9ba7f532431052;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h156985e2895217e4ef1c57e332860b8c5f40bcea6ed147f6af2c041dec66f1cf4e1f73c12ee8ecf8e936e443d48742ca3f8fb57707408c87c6855ea6912406a5e1d0950fed66ce17ff15ecae0031500b49d2b59e20fbc1b74fd6faf637c4d30549f60b2b4cd19204712aa606da95cac540f5c6fe69665d0a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7285f3ebb06d5e40ec7fb17a45287f6196de609cb7f87d956bb59e3401f88a94d8c9dc5c4add0c8327e0edf929a04703e369c0dbfbe9e8cf5b9b64ef81fd061eb6eb02e4ff43bf369a3463bf016adb0edef53c000b595096bab42266e41859c4cf606794d06a9b79e3956aff0d3e54370c1a70c4e3ef221;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14d323d90669f2ba81d20adb2a4a470dd95273e226c8d6c80f888c1f5b56bf419dfdcd22821110b2006f4f2a039367b21ff86b3a4f5f9becea415e0cb60615f7e1d69c062c1d711dc40556841523583f4821e4b889621cf380f028a469972b04ee54bc7cfe1ffecf771e0a23f29b6577c9ee56dbb64264994;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h129785117e2e93c05c24845fab0c743223e2a328bfb6ba97221ab111dc59e6bd057e0b0e391664a5f19029d3abde6befde535c88fe48ef0010d9571ac43389c18f35275a1ab1d9392d87ef0ae06014e3298874c138d44cd053b2afb1d537e3bcadae0d54a5600603036ba1a06f1838387b31ee02cf6c67e94;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'heb1ea5e1d223b0f9f288f249376604f19e597d9a089ae64b5300ce1d932dfd7e5941bbceffa66f0aad2aabb295d0dea8652031924329eb5c03b6e4fa1fc4caa13a4cd2222424e8d9c0b3cfc7cf8f343a5925a75f449351804e056c8d412e3377fc19b63c13827a47597c2c6dd3dd0b9ddded6df309429223;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2604a9ea5bf35b20b98b1aa31f08b5eb17bdec94b3983ec2a23f042146dea257a90248f0e98dce66ad1244e764f38499d36b48331943d542439550db0f6beccd584102b2ba0ef53f03c6219125afb3e92b2b9c581d39a75d4e5cc2338e5795967f6da79d9338e2d0e9a724bd4cf02c9769fc89521dbebff1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2f9eedbb3e03df0d89f7a62c8c74550b46b2949601edb662c4288c5e8a8c54a93160822b0e0c6800b15f0d3512d9a6436c3360889a7afb052e8dc6c305058bcdc02b4a20435f295a51eb317fb85e082d8716cc2793959534e5da9842b361d28c683d4fd109ec989b90e6fcaa798291057d37dea1eee4a42f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbdd8d5ab8a5d982131a90a356490d0d17ee3c1dfb732d162db75a7444ae252d30e41a3c2c70cffabb5db4e7eebe9fb296a00d71c9a519502556c97ed46e0ae50f93e400eefcbdc0ab75beb28ab2c43ef372b6e89b7411b31f92f666cfcabb13494d48b31f00e89655fc5e5eb21fc96edc7bf719931829963;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4ca9055cb48b5b9b5a2bc8f4378ff2718b4c460c47822ba6a67df4ac6524bf1613793741a54f8c3e3516ef5257e08ec66cdee00068ced9b49df3ad7b64245f8f5493e0bf21534f3b01a6b52aa6d7ca6aa83b87721fff66497041e014721a5abc45e275acd52335433755b5ba94a0e22e2df36a52b83b7b82;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h56e9c2fe12ff9cf54ed23f7053949b1be323012b3f3b76b766a4344679e66e5bcc78e2b0d3fcfc4b84ae889daa3739f4522652a3db05cde3b3bda7b88eff536dc2f7715095119d066f2ec3ac83e3bcb1d33b2ebd09a90aba0733064bc25100517491fbc0ae8183972e554ff1dd2cd7c172b7af8c8afdf0ff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he8bc6e4786971addb4d03694ee4bcc3a4fd5e172bd0511835cd9c85531fb1a081340aaf63a32ceea61d606b3a6493ffaf3d19ece58b5d1c8f79cce0dccbd0900eeff03226823c7de8abd6fccf1c4366e5071b1037df81afc1a5ab28c8de7be6d16dd26b7acab3f5b2fd77289910de40d10e4c5cce114241e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a7de5f2e040044fac1263141854c6efe294ea412946fbf51a74011ebc5166357cddbec7f630da2cb5cd999a1064dc810ac667fed78a32d24450b02deb569d69e0fa1f6a707618be562b6479d60c5ffe66e1e011ec90634415d7c94efc39f90bb5508a6600212f6d67a644baec44f444ae02e7dfc5d14c54f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6a2122058a244dcfb0aa1fc0acdedf00758615225ca7e5eb5f02bc5444b6c2fc0a4144fd893e05a3b389aa03f8c3172ea922ea28702c5e655d17aa27b2ec02828baec06c0bd352928029abccdaa336f320af3ee09df1ec15929388ddbc446619cc1b4fc8b26a33652fce5a1d0143e15a17a934480e250ec6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ab0c1a12402c46e98872baa8463e8d9a5fcea69a20d5c3101186c393094fb3e2bafc114e994d5f3dd042195c052939ed60efcc125767368b84ae94bdf16c37be58543b40dd13409a1c9069c1da71f5893d34544e57dedf4bf20ef1e8479412db2d28761639186b1bbba2445079278b5be5a3d775a82c54e9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18eba87d0511c33cf1110e834696b4ad9c040262dfa206a74a9f1bad0d0032dbfe99287a567d0ef6292c9749598997b7d4c399cee32dfc9996c642d9e81bcaef7245175f2780466d2759f5f00586a9727d1642641358454ce22a3f01941513909be85e46d2164a1240e72b6fb6457276234c13955cf24db2d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18eb8cc694516045e8f56a01bdf9bfdd81a71b80b18f96fd7cd15f8fec6be862bbccff8e6dde49712952f80f94acabf3b6ecbe7edf3696df14806f4f247c4bf8789825b0ab87993055a167f0c0be7af2fe0eefea90086ae47a2e0d98465c4b97b8e1e9ee784fd76398fa3302438ee8c4fff483bdef268866e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h96b93b9cba3a5080e91a3d10e318538426e9fe89185e6cd259d18395b72aabc0542a0d71a2e6041b06e7e9445b109a7acde970fb03ce5d7e436a1e6a7d5cff2aba3cf7ab0cebe9351d681d9719fc74f212ac85e3da4b7d5af751e3fdeb6f36bfcad667c31c31266bfec2dd32e1d575e391d05009b1f9a180;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb3e65f4d3454734d9374beb6ce09391f891a9f50a512c07f582a64d8b712464940ff0aedbdeb98e5ef854fe37bd664b73ab5070eecf2895531b6836c8585ff2ee5ebaa9eedf0281d61c2b156c2e24244773e6acf4f1a24f22a601c8458097072ffe83bba2c3e9e57c0b3a037d79ca044b1d99c6a1888765d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10e7ae14444119d8bed67bd953c5d2ecd9f83c4c83dbfc763843ef8d09ce157f1afd60f3d40e8aedff09b4355add4cde297525e7c90d7e658e6726832e61fa30a643fe1499b35e848f3d730d98bdee9f9370f2b85875b07e3a42deb59469b306aaa372693161871e72982d6a5831627c6b1e5b9ac0346d020;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h166d55af31537a7e70d56b4c184378f8d40e954514e6a1bf60e33037e1895617982e5d7a5054d8893e493d101135fb0b511b300454a62e4cbce8225c50ea1e9c7eb6e0d3d8fded055f05218bf636a086d27bee566230406dae016055b70778eb8da5695728caa3d1296dcfd8de5d32ddcb987243532be1198;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9c183d928754e9bee960ee5e9f9b701bc6e193307d5d9b95a3d0b35dc2dbe15cd0b6390a4f7c765964eeb6bda0bd269c7f485065562f2dd556f82ce9116c27d27913fd3d0da24a8e94da962a552a48ed0b2d720616d8ca2df86be9850d4c3e55fdbfda88eb3c41830ed44bc5bac16b374a9d27939039615c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2102da30bd66dec7f823db32bc92654ffdd69fb4013c8a40011fe6d2784e15d0d69372cec0931d500f205739d6cb15d2399d8fe8b936b89ac7a9f3ffcad6f492ae39e8e063233c34037658d18e24669216ab6a7a5500e913458e3d047a72d580ddcf58a28221b8860f5b1d8a40fb60fdc8d6a3dd550484a7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1822645f9a0f503d884acd72c978f784eab9f6a667fad87374b4e3f4cee0ee5f056676463974ed1bc97fa7901f12b0b70c7d8f11a451b03550c1903c78f85db4c70c52950c5a870c89e2d7a3cdcfefee5dc99a90dca0504bac49a366c311599f6d92ae8391f2023ac485210cbe2a24e9b5110233fb0b17fe8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aa4928299ee9e773dbf08f63413e3374020b457a5fcb56968f9a856bd0187b5005ddd73614d871c8b00e741b009fe9d831edad65ff4f4ca52cd4facb8b891b39760aec99413fcf09f0c319bbe716cc6591c9449190b1c43e0d90885d5a8d1e5734d90b23315636ef8a72ecbf1aeef5a9c2b7de547f2fe9e4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1863caa7ac57943e05115e980ff4ebe6dfe23503d49ba020a164423162efe9ee841267c4a0f76aff2144b8ff25e87070030303b85bd6933c8d355aa5678c789d6730229a46e695e00d06612fb0bf1a47357421c647587460fb106e482d05afbbad8b9e4492236440a4fe7b33c67b86decb3c7d2d3045fe4f1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbfc17783a7693047e692c8727bbcec87289837bc1f59b59d2afe46db3098b029094686c5065e40bcb5cbad9d93e05ae2028d9cabad0bd3c934865d2620b853dd2e11bb1f9f7e9a3e8e841692c84a7ccac66f7f1aa1c811464b65bdc302891e1de2fcee43a85450414cd13dff6209378cac101a883dbc13bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e9525c39c5faae9ee79116369649314a64d6fef6feb46aa042096c520963812180ac76dc327a95b1e524a27c8e4cb081b92442ad6cf7fabfe6cfdb2758955bf3aa62e283a5ddf605f4aaf8b6e9654745beb7dd87049eeea69b4cf97a28d5bbf82b63c0337228fbefe5869ef6903c5f95b8cfbe18b6298666;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d3729e057bb77a8bf701d7e4235d93f32f8d6cf5c138bd52463f0f3bc4513be91e21300193ef7e99f7a796356400ed30ce50608ec9d85440c48a5e8adb7f0902b124af5c5512e4295f2b96532e551773a7a8cf4e907cb3b45f2dd390f0046919e3fa8296ad8f4382f5d30f9973fdb1ae589709f934eb7bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16ad5b4f35a2c2e1bab81730e661f75f36a97582dd7edefd81a6a043fef86ef0d0812154e48c6d9ad04eab464d126bd87b3c3ec4b56d73050cd7df14a9121d1ddca0bd66ac87dded7a78f32930c6938aad1c71a97407281c465e20d5e8fe4deaf182ae8a1ead8d68f1610e94042ce65ef7c8bbb1e7b3e2af7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h74452e26622926811c0dabc0c997d7cf76a35e8ee56f5608bae09d0d144657b2b3a1fc8dd57ea93085734e734c88216e59c6b49782e40b89474df1df7a076a69c71b5a6221fc1ee6a885668f6d3801fc44e42112411920ed62615041825ca52ec88590f1ebb697cd1e14f3f9ea7f2824e83ebe0c789fc7de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1789374aa28f90984ccd4aede7be4ce42997e4fcce680063eea91633903af2860798f7020fd490ae5012b0ff80fe7a808ff3944e4456a166515a2d12ef6afff02ba768d76848b58eac9122810fa19fff7ceb24d775af17f1efca8993b2a01ef9406ffa9b2d72b4546482a3cff0cc40f96a47b5dc8f8d1fa40;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h141b5d4c1064404837418212ef505be0401e0985fd08025f681a290d03b218ff0826f25ba99ef6ba3d118d695fbebce4465cbf1ad399d9293cefaed620c22ad3d5dd565fd7f97c73c1f9cfe7896e2b62fc8894960d89d62b1012b96ff35f24f774bc06abf55febf6a0c4805ebdc90c2664004086269730ee8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h98de684ca278b3b7b2c0bec5d2421a06194853a3fef4cc35afc7ad0583db9e15bba09e0b1e092eb751a2029392fbb8dec16afdf365dbcf0c7c4d6ed2818f63fb9daff2133cf2c097354a22a7b104e84655628ddd3451bff651b9c79ada0020794a93b5bcc7177425ad28a4c5af29cc4f3b4fcc1fa7a89ee9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha7400090437156a3ba360ff9ae6592bb17c3fbde489656e9d8a8abd7b3648766aadc98d6d561dae2eb2427eaba743678f31b69938f692204781e5c7eebddc2d18af434b9f44fb4f6f68865f23690bed4af3ec0d496549fffba3726bc794b61ce35152d520fc082ed7929817bab317cb33c990551dd5ac25e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc5115f9e3debcd5d16d5e4339b6ce983928e5678afef6d71ca10e5db9a37f99f7f9a7ba19299cbfe9ef3b203119aa659795c48e7709bb6400af6e6bfce864473e0426ba3c45bf255dfc42d7921f411b85ebf90ce6b9c6954b5ad6d76e9215c1de9f2daed47cb2d00ef4c4c2ee7a5a5c10f4f040441b609a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h65dae1c5fc99694cc5dd25b5f62d926a65d7913a32ceab946ed17cb44b09dd06acb8e5cf17f8ccb688775a3eda3bacc6873b4b84c459bad6b61d60a1a93e61d1cfed90df1209d077d3fa2dabb8bb2bf9f72e0ef73e2bb155900aa6ba731933af841011e6a553ebfbffcc5f2fe0af88708021c570c65ecb0b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d3e66dff465ae40793dc7bb2953203b427575c5867c9d3b7be77ed2f33ff36504e57cf7a6a145e5cb75319d92ee5ea13d1acc1864298777105297545c846d3c46ec26aba051c91ac61466c5f674d90a366aeedfc0ad63bac31e6d6d0f91e1464927dfe97cf7f4b2dfb8783c1a3ed62761118c0ceb7f4e152;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bfd4fda5ec23b765370a75888499a4aadae5263d6a2e00ab555d21d0492f6f1e71014ec0cf7746e50647147805b79f100b74906c2538be769fd910d370b49beea4af4f42a273e4b4d14c39be13635a5e857184d79f9ed746509de495e35f699cb5f2d6f0423c397cb98c01f92ae2bc82526d79871df48d54;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c27da053ec33c917a0c9d8a7040e191a60165e6c3869022895a391f502389cbbf6954b5bc5d643864442204de9cb14048cae4ad8976c72c6104909692705bad6643a3af3432c8783e5b28a13d569fd4f4f635bad3467f2aa970c6e98d7a4de5125dfacbdcfb59109e5b9d867568f3eb62d6e397110b4880d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1343e580c81a7a69f7f4bb04cc300dfaa5cd14f31b23361af604f37c70b4133fe749bb676b36b30fd17c5d67fb8a414b7cd832550b429316c0e3b474b53216dad025ce17b04a3133c896bc6d8ac10e8f4c1cb2c156550ec0d577857485f3abbd8ea75e9bbf03682e12e860aaa96b2304d1609642b8e886267;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7a3269ba98ae8676720a920df0fc50162b69e577f0488dda3febc57b21bb9e50746e8abca176623986a6389941c71f7033551477fd4d73317671d8ad964d4c13e7c778768c072e45d60d11f5fe92fc48cafc11d21a2f6fac63bc26a70ee33bc31a7e70b3ee2fd98e4887bd918128d8275c5784608691c279;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h105072be8df1780b54dd49ed7b2c2f42431f9cbb702fd0f17101305bbee816da30dd52214ba71b4320c6e78890391c598a102437d4ff9c752d4c64e4e9f788ee9bbf4e5931c8166f8b6c73c015a65cc02bfc976b7e8b0822187a1b13de68382f4f8ca0e7329b53980b9879991643b05b24728dc15cf2544a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h485a562281862e48558dd89788b17e4ad81c44f1e4133b0940eaa9c888d5e4a996499ab1faac3d25e224f89ddfd721b1e2a467512b421fd3c52a3e7fcaf067af396dfe7e81371bc45bd8af6d807912640fc9df5dc70e98cc9350d93eaf69ae759ac8c1a97de7cebf0b881008419f6b65d37a51ca508d4724;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf263697fc357153933cdacd10e33f57da59409450b20f2fb470f593b45ae8f1d72b7778d7dc6401f263dd7abe8583af742ce916b8615dc1828bd93eba41b42c762d88ac90dfdb5a6062c1809b9d3c27fdb54ec613a3a02cec4d5f3a14608d4f36812a5628eea68f38bf7c93a99ad7373cfe2f4bcd0c8b458;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d0eac6493981164c96c821660ffe8b9da850b4dbf82b7393630120845537f92500ef6c4c6fc31d2ce35d56f891444c39cc59e73648835b299ed011a14592a41fc9390b1925788ad0fd256959e3a61ea6851579d32fdc3520def3088ec57af0c0d584c047c0d12cfee9150d4c12871d299e7ca5b53864eba7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2ef94a10ec955154a09c7894674954d08c4a0b33b624c14b20f23f82548319a541fdb42e9613fa1402c2eb6ca9642fc77dad22767547507894a87c18034d2092495a69488a2a1021c1e28a8b10dace93f1283bba16a91a80f19c89acdf2b174f07b6e1099ee30911b0330907dda0d5305d53eee4024af10;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18730fdfb6b5528b0d15f8b6c39e805c5fa3e5c2c227f368e3c2d369e3c2ed8de2ed8f27d4d16caea8e7cc2087e3df109aef8cf418bda094f1e7c1c941cf3653e0d9c19049527945e592ea752b1c558a5a314bf33c69b8d45a1d799d3e7d84f935590b8019dd9956919fde7eeee2e23f9b830dacf63db5b28;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9d41a2ea411f626372b6b4a9846d922373483070610ed758e7050a791b818ba45124107ecfa1b2fee49582b18b700be0f203b3b803821c78ad7ab4a248cd868763dd8700f305be715c151ad507b5c094ea5ea6e2557ba779fec46c0179ddada64e31fee5d998b2408cfe48c1c3101a408a85bb454ed749e8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha964b808ffe4c7de3adf06f575144ae12d20204ee1a78c3560c7d42d19036a28db8d64faaff0aef3fb3f0364a858b4aebe0175753bfe8adbcd3b4d28c28b1ddef328a7c3d97f3130ffa617133a197f1019d0ad2a835d3f9cb5341ae42497b42d4fd50fc601a73f38dcc8255ab6870128655d7ed2c9195a33;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haf3657a73607e676680d14c0703bb81698784c11c68177c9bd1f01a85781df837de64898372372e2920a7ea8229efc06eeb07fbf09a60ac14297f1be3ab099128c0f56f05d8ae5fc6e33517bed9ad4fd2e9ca50a2dd2ac2d95f253d91d11c6c4f011ca5fd2c648d5caee8a28f75ea6328b072673523bc3d3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h38c7fef81e7d8b7c7a7cb90d4b3392c300b09dcb9c1222f4dbfc6824d809445c382eac145829fe90906a8fa0f474c64515c55a3f580683308246a5d948341481250915cd3b5f5b706fcb47caad8276bbdb89ce21bfde5cb25ce0449452d47a66d4c3f496595a002e5b37f0af51ed9a6f437602d9491153f2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfcabae1ee82db51d92908483d0c9637f602623b06cac93b5bb5e0dbfcd2b5bf96653d6be4a142653a811d73ae42ed68e27781fb64e8f68425fc591d3a2bf0d8480b424ee358de278d5ae91c65eae02b30aa3d94cf4bbebd65be80c0ea14fc86e2c9b7c9f5a476e8902c1ff8f89913364eabf9fcd61c919c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11ad84019abfcf83dc2b0c233c29f67e6f542f74f367deefa5aeca0a6765d26bfd415d5fc0047dc0ebac68191bc072894f80f867bd80ca7ee855c9cd35ff3e1b0355be3ea25d82d82e2c1b2830e2c26c94420a634538dda8645c71966a6de56c7532a111d21e3cc10c7bc5710341de391e4de9209123eeb4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11a2e676a42be6dad119beae258a20579e1f741459b4b851a013ea7f4a0b134a772a9d09db6f9c6b99a7e8116ae1fe44a2bf5bff02c9feccb61e6b1daaf80735a632a5f7e7873133ac33d34435cd1dd46759dac8cbad78ff7eb69a9511ada20790fe5b8990ce1b4e281d88b75ebb947a5f25147072be67bdf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b5d3c2b667e90f900de1e43c3f3505a83dc49be1a9a20ed38fa3a7f2f433d61a75ac310db6e44eebbab03d552215e123fc7ff21b19ad45d04d930fb7e842ddd4bc1abd7d21d3864cdb2807b6a54d4b698e848cd7579cdd453e8fd651a9fb11d67c7939885c9af625cd1567ab57200c94e24f4a88aba15cdb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he8c762454792123e00939e78d21b01406b3544fc6c7092f37395817e494fe5e9d79f9f06195d65d797652477d4adb56cf1ecb85344f9781c3c606e3932923c3d903e9bb620b14f561838daf1e7caa201361bfc94e6bd3cd447962c32e1f7f8dcf95080ab7156f39c43e91ff0dbf8eabb3cca1f594a9db0b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf3bc00ebf125fc2c3fff07a8b6f3f9d3df7c9dd2151d7141294bb31b782f850e0411bc9d5341e9079f3696c5bca4989d216cfd1b651df1e7989e0fd6b3015ff5db60b13ce29b480c86abad263e76f8c6a8c041407fe46876d50612c045816df9da87a812835a86edf8da2e6f7c399d403063ad3ea8276a44;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11d253b6437737d5a8f6933be6ab013db713ed5df3b664a6be27f26664ceacd5b7e1ea49d8222d07877c6786c052090625527637a681bc585e097ab6086e1e2415a5a28c76715f54fd6bc825b895d1a46d4cefcd24c399945cccf0c4b26a7b2b3896020e2d35b1726e54eb97dda07390f99e5c0bcd0b05562;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf658ec77a72d97c7afe58e929e463b0089e772f71b24881140215c49bbdde4864c65ceb09eaade70eace5cf8282968087442f6994e017b9eec54896001923ce073998a79b8c72885bda5a1caaaca3e735a20336299ab1d0ba9fbcb490fbd7e58aeeb5ca95ec606a3bb59f67f51bb9960a631c6121b019015;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16b824ed7d442765bae5d24f83e9e3e446f50bc9e6a271bc952e814ce079eee1b2dfcfbaec15cbb9a595770a6166ff1ae2ca1c94d568a6d8d3a877ef8945ca3a99efd4ef46b4ee03eef9a34c1c259f695fac120ab6d90cf08a5ebf18f1d5bb08bfeb9aa923a8f3ce216a660d169a709b5d9b8820ff324365a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h33372c23407ac6113ffa2abcdc89280f0fc97ebb59d167e28f5829ecbbd7ac13a0d821df6576513dc0317110a327b699ee2f192126be2fa105b1bff7a52a1fb002aff9a3a33adec3e2f71731f83cb445fdefd999e28e8a53dd80bc96f0f8a95fca48d2bfa2253776416e297ae56d6c0d56cc510af17088aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cccb571fd6e0393b54dafa58e3c6da4c060cf1b72c8997a49f2513f39891d54fcd6089778c2087f9d7d0404111101e6d9e0b3ac7ac2018f1fc88f3520f2425b13980f5e111c31e5147121b4bbc1fc11544e1ff2b150872a880237687de3e8487a749f26788aba55cfd6d2737745884cc387ae1e6fda02fbb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f9ccf58185da83abcd49ca3113af83647cbfc85ffd612bb8212a8a640545a5190db2541bfc89945f5d81cfde8c9c2665651e38b756f58c0da697979c9e48461ce5e9160241c2c2f73d35359c272cba7271e9e65eef0630e6c9b675f55865bbbe697e73e8142ad95655e8f9dc4758a10c303094d4d2eb390;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ac6e76f384b9714f87e9663e523c73117744716711f9a879c9c576d67018ce61900c84c811bb53473ecf4fd729289251a2d8062aeecd30951119878b1a5a33c49568dd62f97b996a8ccd7b261cfc99af58567f823a39de4ddaba77487ef500d99891a735047ae9dc7f426150d75a44bd66c15388dab850aa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ad82f6748a7dc82ab03690ac967b097ac025a7b5e117d5e6f308864908e3ded48519482657d4402148b0a3808b314937118552337391347f68bb0e888593d01d9e73c6497cd606daae66910993cb686d08940ad02bb24a46930bba01c75f393f1febf01b34b2242166c1542b887a8004335ee83accef6c65;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d3f80f54e1ac5ffec4b3039404e72d354069b466da3fb2177f89a7ad25f567dd2eac5dfcf2f3c5a231bc1624ca9115360446113cd72a543f36404dde050c7c7ae5539487796b0e990c64f95ba61a517a0a9c4b799575ffacaa55473f3ba2b3a4938b82b6adb0227be5518ca889c2113725de2162e1536880;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13862d7255acb8356573e5b62d8a61eb555eb575d46bfda32a0ba3299b7151414275613d6a2cdbe5b29a495e3a2dae6047616a8e674d010c92427ebbe9d41b79ddb91b6d4884409a70e442ff9cf4ababce7079f6370806b0484e473d42cc918ad422f4ba95ef509af4a704e62b959b91c2518115177dd6d13;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bacbc368254170e227a0d869a10eb38a95fff6eda36be9cad5a21459dee832b957bd1bb7a2d007a10a218b4f872a3ba4e15fa9d09e75d241b4083621229d9e42ece4d5471d2e4626851e511271ed87b87445e32816264773639fe6c8888c7b21eaa9ab4a545a1cd315fc3ab6421c53040b78154f88b9948f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h833d9b6bd92bd476430935fc8e8b9d5901ec18ec52bb4343f7e0d440cf7129d6e02a331b11707d47cf545fe6caa516790c71a29d69dedc10c235693602b5337805938396288d170598112719f6ffffbabf4358202879b7e8e7a33c38ac9c61c152dad91d58b53698f0e7c8d94e93618ee97e305c2e973b09;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h66564ee954c48f6f15049b57fbd91d639b2ab7fa12bd6d5bfd6544d85e5d06022fe5d54077502e8837e438add7fc66bccc950cca89f9be1996f20cce39e6e32dfd03b45729be9a868afe6af84b9312428572a905be77575cb4b74c9a77afe343b743bf54303dbc9d279eb5bb4a66079e334835c7e1335a63;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b2369b8cc50e43ba74328ccff3b04778a2007e272293c3bfde2d1d24d248f9e6592a7b290ed019dae2c3a6075e25dfd37c1b131037dc4eb23135174d8cf6d39d189e33a333cd3cf267bec1096fbfe3991be38eaf4a75021f07c8dacc6d6478b1548d3502694b2eb8683173d78a2f2a565008061c8b783e4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h119c826e29d194832e24046d49fab44ab37b742f222c93fc93ef8aff87264ff2789847760177b61ff1171bfd94dcbfef96001e91341c1a1bbc94dd3aa19a7de62ad9a326f559550661c0b86af0b591ef0119ff18e1ed17e13b47326c3b68bf639364bc82a81cfbce1600bcf36cd1fa2bd004fca86ff2f01d6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b6112047a4ea8e61977e2169c52fe8c49a4e9c1ce8da7b7ad11f255516cd2483d1d7b11af8535d4114208bf60ed4c4490c5680b50251cc44bc7655deb179745277e9b05db5cca244ba2ae2c4b9e40d46a64e8ecd83b547dcad91de9f0788e7e0086fd5e04795109237727d9a41cc5833710c82163daf07b2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2cc077339718c724b029f0aab273a1384e20cb70d82fa629b087c22bae2ee7aa2c56d06ef44c0d1a6f1b710f2b1b8b758f2c3f22e7e326d2eb2505203fbff92df1dcabf7baa45a1e5a1461874b1626493d6c331e93c6fd9d6421169f0e770bbd87b4c6f0040a9265531c4d9d038f84d57c5fa5fe8353c646;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b944bba7e90ab0dc0b6056f54de099aef7c1b785e0f477a8bb6a3c32256568bd408c45d0aa28f69e713ffb7dd95f7b03fcf35c98f82abba868ba6797749c29d4cf04d3e48678c0e83c1f14e893100818fe8b1e68d17d37629654a05dc1e1f1fe3aa6d0be0af981c5eb217cc0fc2c7f9d2b85179cd2a599b2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d73a4ee0dfbc551f057b897997f155e78d6d8939e0e788d2c12d8fff55f721800762160d64ad8bb184c8f98ec98925c65149582d51b21edded6a243e0be2d6b971370d1b29f7abad86455c5441c358d93958a75ac9dff88795abfbc46c015397ce40637bcff5790f89246c6c5db05f81bb40c3b36702ba5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146d3a896f6c92f5c2f7fa49f0cd81b593b4d3c61de03cfa6fe2c42240de70e23fb75409bce9f09ee8e3674fe1235c5a87c2fb3181a640d92d5a04ec9ea389540beccbfe23a4d9822bae3a63d8f4ba1145e8195bd4b4ead1f29f77a4cad08d64c946a257236e156a4f191d98833102001d47dfd17f27810c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h118f75dba41271929b37345f258c6dcc9be160d8d80512e5eaaa24e5c592c4db96228f1186b72d9682f2b6c31cc0816f51b1f053fa79bedded5767f521422985b8c526779154baffc3c0ec778a3872b0c82aa7e024eb59529cbb8f0bf66a742badbd998968b52c64cbb13206d2297cb26fb099e2c5e50819b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h84822de9b4e150e67a40b28c6bc68888f3bf09242caa1a8a9df54bee7f913a1ddfc4dbfa9eba920419613f7e440142f68641fdfffc5624b3f91b313fdf4b799407b7acbe5e6b6412e9ab8c89284474cec9ce08b519131ffe969692e55ff584f93405e1a4d32776f0427b53ac0bb0a3902e27133f6baa7263;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h65babfb7847327aaf96d9687ccd155d9d0392904f1766d06a370d1637a9e8cbe64187d2e4158616a44732d03c93fc6e3c7bbfa7b55ae4e15186cef11402bc85553e5e58fd37619db70ba4ebe988f82a976be70cb25ce2f63387f3ea219303886d495eca5f298a98dc314dc444c50ed24ca00c2fcce158e4e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9a69c06bf46674d593828ebebca2570a9e2e42f17478caf13f3e760d96185e13baa96c243ea6300b5b931594abc261f42c10ad669c9746e8f4f1b31f7fda5c27a2861233dab4d31e620ca9dea5037940192036643c5826ea188eb1bf6e301fa0487a405a730453840569ad369ae457ca4dc6063f70525dd3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6f4060974c83831bb3bc04330282ced3c63241cb7237e192a1667f71694ed50ee578f6813ee6d2394ae62fed7d8cc0c2dd21237cf1dd9ff123c40c0b3610c6c3f384e49a3a68be44936b7f790e177702781342fe20d97577a9b7237a51f51cff521b85805897862d594fe4e92c3708a76b42260813521f15;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1daab1b2528159bbca671128e0bdc8dbbfc642c3fd216e54ac48a0621f9d0d17ef5943d839ab7117230f96b94f53e5d0009a779eceda2c4a85510eee9e8a3f187d094f08461ef1bb3183cebaa1f7cbf79e7fb8eecf456e84efd81098077c3d2447c0ab4ceeea6f9abf4598912b2f79be11110b13f801beca8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfda87b3b09dbaa5d22d867ccdaeda1cc5291f47fd63156a4094937cec53166b5cbd57e9b7d3c921592074ec4ad0720f0a4d8b48dcb879338429b36340fe1343d63bb8830910d09150c49f9ff3b8915147d8607ba42f67e0044e944d65db7479b0132a615810e6fe2554c4196a281d96b3b491f6318c0d5c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1554faad46f31341ff00421b480969a13d29146e970bdd12f5899b023d60f576736c53e57ab01629bd4323eb677559a070cd51e92eb09944918596d522862b8aebde26fa21de6135b9b014446f2d63d1c4c2ebb66d37f202e4c88abd61f65c7d60ead563726ea5e97bb0f2c2676a91e3df53ab065b59c7c2c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ff4c20d3ffe00eedd3bf92685a02f8379399356a3ba2f72e51b57b5b91b3a85f9be88617deb3ba12838bdb999720efff784081e06fa1f50d75ba62266cb63be313aa5a745e64abe9845c909919d5accb452c48fdf5c7a31cab59c89fdafd9adaefd05f40d30b1b27e92d9350c295c7ca4efb176b9023776f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h63a96362b162af7f81e582a999103b71c9aca2072c55deacdfe114e0b88ebc734f40415a6dde925c482ad7a22cbb2c36ec1a2f77ea1504336c70c7af5227ecd972fb22424cd1a54ef67c4f79daec5d8b91c5addb74911472485f0fabdf735c5771f930ce053cd17fd41d697318c9ad8fb6c64d33eb8f1642;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h341cbd5d53b8b634a1f80364553bd08ee287aa6a13f5980ba648842cc30aec2159071f8885fd4cd15b5305152bfda60301f2d6ac99b97d5403c56b147c014cc11d2e7c3cdff0bb89802486c27d422e51b37053e25a2a9059806d4c24bf88e3f4bb71f62c247c4f59f7c1a1e2eb9cb41229bd6a4b348b1c19;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf29ad7a2a3871aea00b83d53c1fb3cab256cb032d38b28f79f3fca715fa681fb1bad38f6c037c36d4ed90bd76a02aea88bcfbc609f3f9ba8a8186dcbfa18aca93273fe9ae0430a804b9964622eebcea9385f54812fb661c50f9084521a363a8ac8d85620e845ab2bfc3e969d9f02c8591ddcf22efedb990a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b0523bcec9754ce55555954f2760f0a984ccd6d7969fdee71dde17182c641da59b73608925162d73539f2bbe691750819807ff39306795e3cb3747c69dbedd0c86d375802346ab09d215beee1e68ea8f260c105169816ad7b11455da85b86686f405263644db5fc588ec85fc72b4f89c888cd4d642d093a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hacd4a5321a1f0695663233e5bf2d73a73f5ebe23b4a98e6819b0bfeeef9f5284f6ae8d172c09a302e56bd1f6a3d44d648b2776237bd810faf94d8323b51ec113a878a9aa581e18c2f484d9a93cc857f543bc56f4245d64835312c30c8fa8cf1f2a0e8677659df216f4bad3108d3a735acf401f6084acff68;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ae503f0c4d2cc1928e7700d0e9d472439ba2dba5e4d62ae790b6628d981975aa257ba6c65579c26c2058ebdb945d078b2d5d15b015b022314b68d589e554aa30e2b767565c96000fe5a9e3151fa4607bc4044c5ff30caf031b43c0d940b015e2f71ca068a1a45cdb917586f70de5d82b31cf432d4f60ad13;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb2c02aab1941a1055439a125e4fea9b30048f3fafadf25e62d520bae55ee0c2451908d89ab9a804bd2c2cfdd808a7dfe6bd396d18b4c830c4e36725aeb1d22b8502bdf886b0646215ea949481dd3261b0ba4168ca0dddfb5fff5dc7a083c6f8cd9d5e334c51df14a95db401faf0cb06490cbc4c91781f909;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10b57cc5a04ecf6926d4d45af813c576564c19ad2e51f5523ffe55a0337aeb3d746790508812c3206dc0c2e6daf14bda851d3e6ca5bb50bcfa8c47e97914e43609adf979d99713d969734f76e745a1d3b624f8a2b9ed22d7538ad7b8ffda899f9e244a70a9a54a1c5d5bb997dde2f0149d386fc3b4d40911b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b45378a23e49c9a3b95dc9247e21c71b86c4115e4be53e2bcbd8aa69c51ea20fb91be8e8ad864eeed743cc22f022cd48000dd9e1542f3863254a829f75938de0f1c66ea0105f12a109037700123569b0e21da685556e2979c0bd8ae4ab32eece4d35e7047c41bf3583c5964f5de2033e02be6b82d4a00108;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12c3f97b36fcad0b02528883d83571afcf8fd37a2af55ac9515192481479e6370c3c2553a1653c2aab71ebdb331e5e21a624119ef7cb5ad5343e858b92522cb9234e73cf7fd8364d48d02a8ebbe1bccb7df24db898d42540ffc29d014dad6d6fbac389b60a5c6abbbd0e88499dc7ac8175b62a1648dcea83b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc029282452cb8708e13643d3a963358ab9495569686e6b61b0869a28321bafa8f26eafcc7a421433b030eda6c5aca5bad1539b47b6f9385d205ffc94e69d28743787744ebd833818b9af114aec3ed1251241fba2f4c3347b3292cf48f6ca1129505b93a9d5348dca776296165167f3ee088a79dfb812a7c3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12f5fe86cb87ec4c30441a9e86e3883ca3b7af8ddb2e38a46372c11578e2ca96f6adf48783713613528f7be888e222e1ab459b1715006a58abc959bfeda747fdb86ec4e5a7070c05aefc6af1e3cf4bfae35084448f90e04e469e3b85171d39d749842661d844f013d1817618e6ca690f9d5c1cd428e4856fd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hfa046c44ccd1686dec7dade48260ed01444dcedd4ce0512bd814e853a598f077fc203cb6448f91b8e8c5e8681e4e8fcbbe99bbb32196262260bf64b9df779fb2c36d0815b703774674c20c316c6cb8ffac1becba9113f602dc1232e362d6cd6762f56386d0a92a581c53ba8960d9e7dd931ff4c7f8118406;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11e4404cfaafe35614813b8315ce53e18e9d73dbfe3eb406ea54cb92dbb6a145775abc4d5393a26f6d6403e23f27f39663ccb55b2f781f06454a5180fb6b4e06c27793f34282da880edb4648cc4cc4169daad29306e4e1592ef20ab5341031a8cef1d33dd96331641f29950ac25876c3e567336aa176cb6df;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13ede675b52a261ef84e7d73cd1b3d92f6085bdfae513af1b31f9ca445bdd07e271528a68cec3ce0bf244c2c92df2b77ca7e0388d29c8cff5cad00cf7121c811a4ee1f25e8b6ea2c38b633651d6e89537cd9885fc0aef449e32e6e66535f02cf248336bd930b0e777dd146670bd8361df442fa0361f6222a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c5c24025008fcaff601a9cb8f5537e3494f7f833185471f313717e155a5d1a76bc2290fc5a57c867c25f5b929c564921f01a0cb57fff5ac21af058191e332074a5bb17071e9f58eeeeafe03231cdbdac0fb2803d4f880b6bce8410e48928a14fdee24dbbcefd963692edf8b89800e32f1b3b96c5f01cdb64;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7caa4b29282226516ffc238ba04a738aef4c0a739d281ac3b8a7164e207c8ba882866197e5715f30c672f6f24820b0b86c6411cb216c6467de9fcb8fb08a58136c7a7134f3955a4838f69692410204c4d0d69860d047d4713431672354fec5347929d0e5bfbcd22e9f306a58800d1a1ae0bdf608421e92a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf9b28a954941024b6b64068e17235465529a7b3ace6a0e1ce7acd67687486e5fb5dbf2ee398c4f8551b62a132b1a23d85725bd501be0b5ae732e3afd53a36a5a12059b0b528f6c55a5b1af0bebc47cd54f75eafc8298839f6b11607560e5de813113c81df4246d8a571c11067332fdca88938594c92b7747;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hedabc53ad7c5931860a531f11ec32c2fd25fd4fb57dda431da411c55c2c7dd3e4ca79a989729e281114c2069ba6c4db3f95abcb003765a8bd02e58aa41d5a8696f3a2329b84544ad1a7a8a8a3315b19501dce3cc7efbff20e0f5df3d13adc61eccd0bf3ccb64f4c720d4e623a3f04f9b4b592b704df99061;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h68a5866ac9f07afe8f08f58f54b4635fb60df40c8927fd43c6c16c20e93d41c88190f70ebc8220f811fd615114de2b75f7811a146875c363f0d1c1789de1dced939465c362e46c5393c2c550420acd49c2fb716015cb68de571889ce53bb553ae92729dde16dff4a525eb62c8c31fa0be4bfe012bc622cfe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6bf0f186393d2410739d153e4c16f4203c1793176c33f4716b38263ce0d0ee04c45e2d9f2847fdf6b3b59d98d45fc0fb935ef67a7b9b26c00e12c7c40f23664ca8c8e90a5efe14b5e4699b54664ff92c26f902cb656ff727a4a393e7ff1db0816bb648a0642d2a0234f8eeb5ebc7d744d7e0b2c620ad8208;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12e1f41b2ec8c5f79abb8f8f914ba5883f7b00ca3148acd2bbe17a513f4708dc6129b69817ee39733630724df076288da9b82f4272bcd550c8c02c43d4e6de8364643f84d06d49188d41ed1118dfd9e1c39efa852cc6a4309e4febf3d00e177833d9e7deff56110cfb8391a9fb2eb1898cdc9dae16112bb65;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbf4938353701d7bb03e8e4602bb4394de23802bef3363629902683df98c117dfccbdbebdde9c298a95b65b8e7416a466e6cea0eb302969473b451b0dd05bc66cc9b1cf49d79dcaa5d3b161552bf7037d189cb19834f50cfad49ad1d9f27d6727bed3660a8227187b5528e50819a9acfb564fae06727f510c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11187cece5e7d9f525043d38bcda50efd48d832de1ebfb1962a163c8f7deafe5294095c121ff71c26eee471fce1baa79de45d2b844d009eafa021190fab4a4f1e68645a1e5f43082f84933f310d3af1a5cce077361fc9a79701f6bb3cf0ef046147126b706f5b3dad678e7146302b54be4cb8ddc575c46dcf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3d3d27479a07b3aa30133082521c749eb0571cde5f8e4e108a0b5bb60153751d23b5f87bc3b66c5d07ea16383b4baa7b526dd32179d4b11dc1454ffd71c1b1d315989625044168d966295234e866cf2f0a8e84854d543be07bc0b1972c0ee25513a5c5521bd2f9ff32613e82598b3a130445450de0b5278c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha33f2820882b30597b6c95687624faaa49821835ddf413ca5946a6d6405471c03780c7bef7ae8afe2afdd6a8b3a8d1aa0c6be7eb48db32e92ca5afb20ebb7b2068a379d3926f1169a92c25e5d331b1398d6351b774e6310797646a68f15a6005c166dbaabe65f8f39ab85767767cb046bab420c5d559dccc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd835b87913fc5edaf4b31e198b2d488c216fbee74428d79feb5388243e7ff7108d5ce5e8531fd4ef2d18300a67924e4cfbddb3d076cca1ce20fae7bf7427ab73a1245bdc73b79b3bb466be3b523c95b8ac1dfdf7f32944df74db0f44a0c1f454b2c6e975afc337f3efbe22abe7f7f15a85331b2670976f0f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h739e212819d2e2e73577c0920ab915b4202da18e8a6170472e95f355085bae67a34054da598955a1949f605aba92e5fe3b03ce6c14a3212c5d2f2ffafb7d98ed1025fad39619f894a94bdb3f1fca89f632cd826e8a385b4e55332e96cee57872205c32f4746546fbfe7878c809aff353457f2b3855dcad20;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12b8b6ca155c7f47d40afcb086ae98e33683b9b6cdeac1835a7d28a7c6ac7333efefbfddee483f9290281f4c85afbde980d3d8a2c32320d175fc54b10952a0172a528cc1d6862c075c9b9376fd90e33864dbe498d60a5753ad611091d74ac78dd63b304dd3fdb2f6fcb288cbcdbbd31f6e08e14324d2ea17f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f005b81ddc604e37807869eb5b4c9c59eb34e6a225f7e18e95bbf241fc1c6ad5ba6c24afd859ce0a19af93833b7eb0dc268f418bbd8d196f6ea0f4d701c955a539b9c77d6c2aea412e8b58cbabd6dc70c4828af9e5d331942321a878c6b0ad2c1dd69df9010f72967029aa1b304014c033f386c6a753a65;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7504ba88ff0c18bbb3f42a172e44121f2d1e3d9480b1fb4d2e1a076cc5e059d032fd378c94e740aef7bcd001f94365188e85f2c25e2ef67a413d6f9df2736508e319df89e3b44669d43f321cf4c4d2cc8b4fc5d9256f326a0d70eae697d3ed8d3934502269b7deebc79da8cad712aef48afeb20aa42bf602;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1620c89c633be41f780ac305fb6d6c805d922e54dc2013678eb6e95ea935d8058ca2127e8bdbc2d8a50bd8368dc6029c082d13dc01802215608062b11d3dece06b53e522cb957927df728b5429f37ab58b5b5c643258f84326a9e6803841d10120e4558d5e325e4e469a3ca7207a8e6b6ae7d0c989fdbc325;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h71118936ed9bcc4375bc74a078a8be0c05978ed3d73fce2cda4e8e65fa6c285da2fa750e2bbefc18bba1989e140a979becf6d9e9940cbe321fc6700568ff02d7794b06e58d823a0ce3cfd75b7601c31ebd4e46101cf0b713409df5eab8c2b1b162249da6d5fa533dea4d880b05d61c8ada5b971f6f2cac08;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4ef02b61ae4d013bdba9556ae20a0ff446f95b6626fdd2bcf3db710914cc6415befc318741f6754333244bf07f2053b9705f1b3282fe5303a03a285698c35f4ec94b2f74a67a97926f8602e2046bd9a659e761fc7a46b5fdb556e0d4df1c08a8279d26f40839583a8a88e0eda91a71ee90eff35535f61e95;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c0d06ae1bcd8038b8a6a541e4e7e4de4f7ca4bf0e319eccc41dc104e891788b24bb4dccfb9aaba8ee46b67e62ed498b611fc6cdf252fc796522a2c797bd28729dad06af220659fa9f270fe1a5305f84ddaad767274ad47c745fc36cac2652768f158358ade6e657c9666b0d05c9c82ca9efb4754d6337ce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb7eb4e7b95a17ea61a8f86653604122a8d8e7d790092562a2c28471e5019c1d464b3ac1b39a535a2e4d9e0b49f6ef8c25a1fa81a1dd58f13948219d663e2bc5e6d19eb1ff34bea0bebce1e99b1759a6d9b62e2aa45b4e65b831cf862ad1e30869b7c634bbbfb7f6bf8e95dfaa3aaa34a32b62b8610bbe713;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10a347df09b36336fc1f2b5f6baf56cc48a21944289da25c7758d7910b884d1b495ec1964f065e7806bdb144ab5421f6fbe97d463d8b9b2067d65f118c0380791cfbc1d0a81696a54a5b970732e743b7dd18a56b9e9536416398543273c517d5f83a0bd4ee3ebb2aca88aca558f6148bfbc71e9ae9985342;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1022f3207c09a02529f020c7608a26497426a0e87b23b28baa4c9398079fee58b3ad9c9bf12d493c680b966ab2cb3f5a274a490780044a5b743e472769bb2094311367b27d80e2bc2c83c1c363a2b18d2020e2635c46518600f3a9ace5a3fbe94407e9be18fada02397942452d369a6a36db55ee714107cc7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h191f9980e80d32420b0b8f84a33c8a374bbe2acef9f76c7ad3276cabd8c102a012d00ae284d1ee05cb3808260f9f20953d2dec84e1d292d472d61ee8db5e06308b5a06ded73dd97e9121b753a867eaa4702a0ceb2b087bda7763386407f9da913aa0ecc72234907f46ae4161b88e1d16dff52eb6a85732e65;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h708403379aaf727e8776dcf4172b14def3ab6486c1fe8841453c089e07bbda9451bd775a1fdd55c52c3e0c61fc2b50890a60faa5237d215fd0a33f29fd57f6002cd3c04cd1933735fabc0af2124fdef6c5e29f41ec13cdac5d3f80c515c470a504a4c48146ebb08ca01911e462bd22909541e2a18d9cdd5f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h83b2703cbd1f7cefb917d92839d183edea884a616cdb7dad7d977c8ea3f113f406ad8f5e37dd5cec78bb5832ae4255d90f09394386603a9b0e13e72bf9f9206c375d483fdeb3b9711c443e9c6177bd1ebc00aeadbeba853deb9707efc6da8fbfdb21cd64a19c193e3fb6578d3ce9c16af1246090c2a8398;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7a86e2843467d0288d1f936ff04e5ff3986b9c213a71bb122e7696245c7a7fceda2ba88298f82d2dbca842b31df911e43146c5cb02d4b4d608d7d8984c7824e1e707f99fdda05a8ebb7eac8682bf4b38a7bc4c97aa6965a3ef4f4a94540244cac5efdb29e3f3dd952d359ac9dde6ca03de4f833ea13c4d13;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h37392a0f341c33d561394ff34885fa075a2b60fa07832305bae95165094c017362164dac404453b74c9d25c40c5cb74d67e2a629f1606b918263df5d39495acaf6c4e2600e7298c883bf778d8d3bbc55e0b8f5827981e4f461aa1d94e7a2cd3d9b521b3381fc6175f7dde29041205ae8b04da042a7acbaa9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10dd6c7d3e3d74923b612f78eb485a523a00aa23fd14e994c8d35d631b13c7fcf51f3041b103a4d2c9afe76f813a451d04072bce7591ca31349bc55a08dd0dee43b28258b23db8d5ad35d0f8c7620fd44e2478b491d6068da2bd91f6751a5cf18a799968491e7e779c6ab88c5d0bede805cf4b27bae242cc6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd780281f05facd66884b5f42df762baa662e8da2cecb9fe4e3647fd050d7e72d43627fdbc59f392f5a026d06ba22bf434bac30a7ce632d38ea6122378948d768016e762991bd5feb52468079f7e9529ff94d01cddc398864eca1b9eae01a266944c2c99e2ed48055bad1a208fb85bce0f8a57bc428952d26;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h771ca2299efbf97ab98a2206c097033086c160eb26a720f9e4bb0ac08e31de32d490ffc440e53666c35518877aea2cd17a121e3618f7e2b94ffe48b9d57daa0c269d0d83a326d91155606f132e6a1fbd5353a7e4948f429f6a78f01b3b9eba7b6f31ed1ac43d8a6e7b2522b66adaafb1db9bde31bdcda2af;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1566960351cfbb67be028924990c4fe2fb5f3bcba05cacb7476d5e38879fd3d74d7a37dc3770adbfe8ba044d9a444250bf06a9458d4033c11a3d23838ddaa62b29b755f88747427367ae8778c2846300025c14eda1233f16404571ed4e2ef3d7fa4218c937559c04a6bd3a54ff622955154ea3dc45c671655;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he5503fb71fdb4262ee604d2af5d6ccb46d24135dd459cd5ed12ebdf9f06c1927274736ae61ea86fd56a30eac756ad10a4e15425d366a233778c743eec9f3556a3fb81aa2e9e9fd8f88b50b221acdcf64c18b83afa2a2e9f9a2000e1fed142f2722d3aac5ca25de9a7da93d11b4d215216385f3681e4b4785;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d49c8970d7d6395d873dbe7862190743e0c20d585ebc756e9f8035d8418083b621ced2f49f0c077f745ffa5d459cd9687e526fbca45515ed1d7f8fbb39d4b360e2330656b3ebd242bff8909688907869789f94da21c533cbcf17b85d7926f45010b6b89c36e17c7caefec23ffbd2cf65fe3f9588b6735d85;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14b06927c4ec370ce58c3b769b7dffd38ce897266caf0903c5d9c9dbac1366eb5cb8e6f13888c60158727f226f59ef84bc33ead39aa7f9199c976cded943488e269d9987a5dcb0d048ce57b2670bd0167cee36fa57c210090666c3b9a0351fcf4f53d20e56a01cf3883864495a4e408065815625c55a10ad2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4c069ead5505bfd0fd3c1ee590afbabf0d917592221fa102c5e5da4f8d756cc39b38cd3d6b5ea07887352b661fd494695d24db73718d7026007fcfbb5a513d4b274d99278aff982c6103e3d2389d4866dacf081c09571da6ebd88fda085ee3ae180a63d3adc66d980843f27c19b57b77109517ed4d709e2b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5f51ad786ad8cc7efc9759431bde729b64c6e641063f0d609e7aa3541c16d68394c0760639a232ae81f4eaf0576ae3eb8569954a632c4230b7c568fb1b2364257fcc61bd9a5c982839435498222bafccb42da38f09217e5a14d59aecabe59ba86f1675f4896e004f48afd11f9701e11beaf18193058a88e5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'he298b14d69818a6cc1a17681237f72f4ff1426f9fb23c4d02d41ad699d95f3f1d36b83a15b10933d248eda0bcc2c1a86ad514e631c7225d5cf7bdaf34f5fb9ffe67d8a857f6e853de3787171d0f18a167c15205b6987246798b9acfb4ab70aa3523037f8dade35db4c33ed501a72f75aca01279ec29bd468;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1829a2c7eabefef6876db84e0b0aae97f44cd68845518e0464ac32ea660045ecdf7ea2a645d6326e7580dcfa6f3cae6a3f4abf15c1ac499974b63f752736eaed3c586336ad28e9a07faa0aac9f83274faabd8ddb599d68180d3f29da479f822362b852e67f64f3c1993d22092c26404782eb81e0e678da168;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf9d6851da30f8881d1aec05141ef463161a48f34b610be329f3f765c1f9ceb9d15894a9e786e192ba5d6d3e6c635eb0a2cdcc3d27e8e326a0e3f3397c7726bce18e8c840b8fcc78259e121e128adf740fb7c8a0b701aadd3dccd275a2984e28e9322d7eb0a15f0c626f4d48f29fa4cd7b05c978e1f09ca12;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f03e0a33b232953612ab3d08988683c6263e0d9dddfcddbc2a8f60954de82429c2da0d8add1cfb636a0cbabb8b2e00ab42c53f690db4483dc8272bbc82ac4d7d534318091d8c7efe376577d239c6848ccc75e12afdc7b82b9747384cb6ab86f477df8ad2ebd3e520e7d9e9732920460f035123a320743895;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h176b3c50d8d54f52c49eb1cbff8554f75dcb12bb4a46b1cab505b5f3a3370ff6a4c68d9220a361306e151458a132f25dcb05ff4f93044f283bac24a7311cb7a80359e77c6bc2a6661aed0e41b807f8179e85a8d40d357e9f4f15456f810a6d69a86a0c633c181bb679fb46b3d62b961a276f86c6faa67612b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1727c24736b460064126d984248b3ff3b2dd7f04f1a5393cef5ff75d811c82cd258c078588a9f89f6d7990472e28eecdb925193484d44c495e374de591a134b5c33df2ddc8591e412536afd0f99a89dcbfcff2cf6391e435c9d42911fde8997b22402b0edff1214ceef358da15b18ebc85fdb9353a7ed2754;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d3e142cdac599dfc5c39eec0f880c5aed8c8bbd355f7070c9ab2b41a1e62389f5b759cb54851562fc3d9f0956feceee12b168eebb549540cfd4cdedda857a6a605f751cbbbee5a80b7f37839be7ac5e01c3f6305751cbdd3c7f5077b1ed68b65a6f879a2d5f1ba1ee0b44dd5711646856a9aa25cf4eaea0d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haa3037f65574c58e7b39d852001252a78841d7e8d3722bfca4c424816ad36ff5dd14f506c0e8b8e015238a82ddbcbce55e847b9083db95a917202c9e86b05620c4f68cbcc2799397d5f55a140bcb3d1dd4bbfcb4647a6f20882576d28d100031622f7a2ab07ce60c76ef71839b3439fcbef129d312c5cb80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h541a7d0591179af5574a0b35977488925a3de83489f7b185d0e6d1961a655b4f14d7c17d4e7d5d20247e8cecaa27028437d388f6c8c6dac8ace5c94ed3d4b1e7dbb7ce3f7e3f5c8c14e90cafd8dbaa0e7b36426f5acd48f7d98ac2aaa96a82fc43a0d2bba13affd9bb0355a85ccff579a4c64c8f64eb4e24;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fd302f797127eef3047fe0a607aff764e1b6b76573a0b31c7e043aa751a9555cd5793d7402bfeed14b3c45b05ae0857594cd001006df5d585c3298acb090c2fbd1812d7bb0567919d4bbfabfeccb6e6b2371dc6b58361f9eb02949e78912fe6aab435310b7d39021f9454df2d77d81290ff857ce147c8bf2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2eb85fe3d431d452d2aecd6d14dcafa3fb6d9d50976f041afc68ec0231a74faffe0e79c44086c9741a7c291d284fcd68a1e2fadf90cef1691adc0be1dff8fb90e2d2c57a801599a08616311d21024426ae25baf1497c6ad0bb93e638037a53aff7133dae26cea923b99738938bced1a8a36402c73c7da982;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h255e6e190396a36c2a2543b357580a95b5165f566f7633edd9a2051e35d3d4008d59c37734fab9847872763ac8f71a470bfec499d0eaaa9f062c44c3b5e4f1ea0cac8c1b0a51683248b8518005f130f5af8e631ea1cd38ccf1866acef18e0b572605257607333bb405e41ac40ec5a444251f9ff5d8ee1213;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dff4b93d78fc30bb0f7fe37cfdc9ba597c45920f8e36f5011b95446cc5152e5a14f605986410b399b96dd618f6ee772c3cbbb88d4e6529135cc679a58b5dbdccaa6709cff99818f75e56304f4eef8f2b54674fc2e2668731e78da693e653c3430dc14630fdb426eec97015389e326c8ae3924811cb73303e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha3ccd39e31e2951f45ac9c69fee60c8fbd6583081b96f542695d348fa5376b68e54b0cc0a9ccb514b6257f96097e40a2522190cb90b1eb4d1cb094e0df192c14cca5e84d268da2bb4c5ec7e841be5ea059864a1a8aa0c0aa10907c6b112a389cf9a65f6223773ab5cffc4674776bf295a8883e97a8995b92;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8f8c9b56df8ec9157fa7296cef6287ff706f95e7a6067b3c9ba9f950394e0f6c410278cde58ce03011549bd3625f781628de00bf705ebbd9216926a72bacd4875a697103f51286b934140768f90f2c78747ff1dacd1ce13f88053b65fed83531431f5507af431d952cde42fd7e41ded4f14915197a55feae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e3117e71c91386765b467d8f46ef50dba0f243292eca465db389ecd8f9522a979778b78147424e9e2bd7a64c669d83601ec5e85c0e55a127fd12311293d65ef90b8abd72620236d487955bf34b8fec1900e39e4316dc4eed18b01a15bcf5ef4c781a67e3ad3446b26cc4da4050879237287d703547f6ecf3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bd190a01a4c54993fe4e7b587160460c332c00b56fca5ec540a2181691d230a4909aaf2fbb8be3269e377a55060fdec176c3145c7789bbc5a3a95352442141136eadcef9ee7e52471282482174ca9fa439ec48f8e9a9e2bc533d80fbab674be60c9edb621508ec345be1ef078b85e9878364a6635dfeb944;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h44d4b0a762b494dc3b0a687d2be4241f5f0bb22797c62930ce2558f100e26b0cd4557572e8e575f548d1ae1918add633ceb0f191546469a1174b1eba1747ee55ca2deb5267c3b13a3fd7065b5c61dd985af610ef3f78cf90c2290aaf999cd65b43cb949794014fb34a5c06fe9391cb92cccd01a6d04f7e53;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h102dd0308bf1cbe10a968014e4c83119a9bb1d1f931655fea93bae0bf5e15e74d33e79e3a8c8ef23f4f89914f55db2309e079a47e1095722f6944c2ec0db61b6f7520c6137183c0e05b30601226084890840d3ab0635f6b082ddd2752cc2f1c476bbd5d3058009795b474d0a7f590ae9afeba4c1691c56448;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a584fde8507e30b6724c15b5a8b4e55b6ef580e24fda9685b95e4f0a9ece4ccdcbccaa092dda3a243f14cca55402cf842b469360aa359d3ef7758f4fbb3aeb5b613f507f9e981fb10a182852d0cc846d446c3d21b7b0052c63a5901f68644ecf8e855131dafd0febb83989f1b5c854b1c88927dc131f9f12;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13437142331c498255838c1daf3fbb8839ce6397bcd161f6b96c1e583fe10354605149796a2de57edc2fadd88ca51a1f121a64dfb24a923384555d5eb3d219cfe3f91f1776aa761633500025247018aee7002b3908d589ea4ba363a67c3e71780566b42a37dd90387c36676a915157bffd3c0d0339852ad89;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb288ae7fbed002c0af298b7f1eda0960af5fa729a67f233c624daab7221b344967f69300d3735281750cdc3b4165218b4d62c1b390f9e5f5c8a076148d8f8b5754e0191c35d1b6adf7a45ce6b185dd99c76ca6fe3b2753844094d5874cbd78a554734c55227dcd1aff0da32d28a463c8276e7d2d9fb43ca6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha1e2c2b5346895dd31961ed5a3f75e5b28a9725f355174142851e302573d761bbb4990fc91ade4187e48f79ecb487e30fedca93ca499e0f0c0613d39a34b2ee6bdfed173092d1cf46c8367ec945e8d24d3c778422bb5cc9087d5f56663445a59c27e6b37c25631f7d2d39c05901732acbfa9790203de0e3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f334951e028ba315a1a238f0869e1da6797361555249bde1a5c0c92159a305de48a83023d59dc199ced70007edbb8e279500fdfe638d4ed7478f0bd56d6ea3a35e6e00f36ec24818f7772c3a19fc71d7d4d8dd83dcba4ae9a4575c55c550ea6797016213017577d98f95bedfd2fd7bbe06356ffbf7477059;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h137948e9c29d533386073ae4344f9513ec0d0ef0e8afdca3326a5806ea8f72dca93520af235347978c342a9c2296299ddca0d53cc986f41fb103e12d6dd2f269fd92cd33db9116d9a6dcacf31aa73e02ceb62412f1eabe827025afe18ddff567e22877e9db275d1ce9ff993bd3f159fa9be128167d97d7a5e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16236111dbf36f94b505eab718b0e2700fc238463b9d86a70db5f4507c82788535ed28d8c9ac2b22603dbd3e7aa3d3e767a69d0751596d624e1d0c8d9995404176d7c1fe071f9c3809caeb32771fc20567e9428ecb8690b47aedbaa4b0fa68794f11b2ed1ab0d177c66664d64545591692e1abf5edfcddf04;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18e8f2f0e554e4027c03a1ff862651d8839eff5c0f1314f625da992a8f3db7b608cb9d0209108390ee71d55a2e046a7bc9ed7ab0d9a0f99ffd636ef2d3d83be3bd0edaf26e902d86ad7d7446255b7f3cccd78d26d3f0893f688789315b29dc628b14f5aa9c34fb60d38cad99c1151bf017533f81fdb31c1fd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7c6d135deec0b297b2c53bb26918e5914791b3736e61bd5eeb82f5d97755f1370a98614d287484a0dc65aeac40374d9ddabd9b9e2c6a9ae814d149832587520e07b2f8d027789e7e0c8102f6fe1757f4ac98484531ae3b2c29e961c742addb2a6113d9400af60d7270bacda30ea9b284a116925daeb0e194;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h155f8631e9df0d9df53144bf3a44d0b1db88650c78b0896a2839a5cf05da36d0640408811dd5efd7f853ccda1ec4d29577b5ac7d2c1692c0a26944652a646f4a8db651a7c826daa6a70f896bdf4f888c4ff251f1062048f321a998dfc179c47dbfe5c4b3d12c61ab2e664be7db1a434e70d61cdd818c85cf0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2593250bba8425f92dbe0f5eda92293c47aad4a646926c4f9fcd48617b73fa39c5b71593bc5c803e9f11544dca8ed821fc81cfcfe7a79354a3aaf718ec5c90e8df12326757caa246737f5f37e4b9366556dc9c4a6fedf56f472273340f6c87e6f2bfc6c7bf459d96393dcc785dab396507d9e4a4929c2d33;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h39013d616acd5329c7b4e9cc0fb976f3071a1c1c56337e5fc68f07e4b84593d0e988910fe1b495a8762b798a4bfdd262f7739d3914204c4c3272b2194f545981da440d612c5dbd6c6e610057b40b0b19feb1223218ecc9066bbc44d3080f17cd52a1d806b07ed9ac007b106166d4f8b12e3d9861846d4621;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dc0be8e79a11426ca002a9a768650ddef310d7dd758ea3985c1a4f5689b5bd18df421409732c76ac4903d354d51ff550351b4fba596b345b71fee5bf3c4ec7b69c6bfb5782c508eeb9f316f33f59876f99cf359b5498634f52b29f8c63985b4b3897dca4f0d5e8b77764ce7608cc4e144dc9f8b2202886e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f984e226eee325f029dc684f28305c781e5d6ae5df3abe85282ecb9ab4eb938dd9dce540a351d19df3d8cff12bfb8aa0efe546a1921e844cb2b05f5bf15bd816d4de338b8a7d4a23692a4f80c1efcce17ceca8740e266980c9265a9610de0aecceada3b428c4eb4469488713f68e727485aaeaf35768a8a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3f6ef4e9952035cf4c5f7bafa16f5916e609995ef6ed0e8cfead21d089c749b26c15c86bb7156f8c44234f7695eb2aae53d29437eae90f1c6807fbfbca19f16d09c803b98249218d12799e4d0b5c038571c1fadbb1b708ac95731a62e3e5e7828b7e89b519f24c0fbe364ea748cdf2d8db6eebc734ee5ba5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h349bad0bc330398eea4e661b437d36eca9ae31881594f99d9b0683ee31beebab28561a48825135e4cbe98f7b67a35f8e78f9a5fc23ac13a80fa41e6ce2f4cfcf3325d708078febbe50a97917139b02a60d1fdb9ebefd3f6928f9af3fbf9b1f2d0128299e5ceaa6947b284b9880df8977e8e3c91b7f50796d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h199c0c11a6dc95185477608e1ca9e9fd48ca4511711cf0f85bd5d0f1f4a420bce5dd538fb2b2c5c6e0d41ab30054e0806906de24f0fb4a464db3a38301510d216e28c879ca41032052fca9d7edbf53dbfefd8485ae1d0348d9ce06ee9c8e38d3c1023cfbdfbc647f7678857d92b47c8238f4a0c3273c2f26;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hedbbac09e4b828c813a630f27742c5ffd4f9121c4ba12027929ec928d1f2d04095db16c2c14cd0d1f93950c72e4fc9a10a4c5092f83a10738dbf6f88a253eafd69dad486c3246b42ebf22ab3772f85ed5866d82ec44b083aa057eba54fc7e085c09cf5969a895e4f1e47cd3d575a5136afcef2a8e4e19d7f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19657bb8f50dc585161854944dbaa4b60345a92ea24eccf167519d21bbe659790a3bbe6aee5fda548123064dd13b4a47ff078bee57215716cea1d7ff5a25bc15e5853bc8f9a807410e97a2aa0aa9d7186887aff2e29d91837b34fdc49d7ffaaa81572f6601ba35f1e2949d38965551ee1ef823fe5b88e2ebc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc5cd59620be0e3a196c324a9265e2dace371a89080c34f97026490cd3c15a0d14ef61d2b88100c93318bcf27f5fa7499641f8254fe413e157dc1c5cd41f540a239d4a94865a12685fc81f30e5a2cca8d93a1ad21eb14f18addf3cf183d3b7e644169d7d07b0ecd7fcf946118f63cb5a2d272567ce57beb5c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e69a11a7fd27a5b19f76d7d868fa13ecb39b12a9d5a614ea946624016fc498419980ab4fae185f49f369270bfcaf49e6f07b3ca9e90591004758fa9086e7ae0e9f3edda85993a504a93a5b273962dfe624e3713cdb8859185c4cfd01f7a6d49ee7b9fb167e7661400361d6748f0effdf2b9f92f73480f96c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fe375a8c9ab5e39986b2b5432f858b1758f7c137b864a2011c176e66cf7a92549ea6fb64b42ef34a8aaf7fea0a3e6846817f8d6275739d4739ebb86ade76c22a15985b985b2fdefd7f590444d1511dc216b3f0d933c9f04ed2b0b3a15a01bcfef9a329ac96d94be66e3a189cc9ce46e087da31fcdbd744af;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5510821dae1446d9598710ab55c65c352eb8c958357b2336b5bdbea5360476651acdc5612792ac5e06541700a74ab960657436fcc9291469289eeac4bc045756f4ca2506ef945b0ade7f9cdd94740d607fd757d647ffc3611fed04f56106c2bb66a4e1944ec124dc30a5c9b7f7db1578ea974011a008d868;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16bc0b2352f64e05cb27354fc3ba60174b5b9b63fa9206242d2b2190661ff48a3895419cd78cf0e2641807cb1275c02ea8d1752da2ba814b93ca5cbdb34bf1f63e2d17b756ba52f06566f7a6157a4c1cdb603757b4011db9604e4673e294644ddc7c9d2435bf4f51267338919c1bcc2128d1b2a8660918aeb;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1366ad2e93fccaf666757c22ffb29ab149c8722e37277d4fdc9d76e6cedc53c68c3aabc0b0fc2ae65a0d293442daf80c197b19fd7f015639312dd19c5c8b3dce932d84848eafc3ceda3e4d06d547e376afb6679408a6a4aaee11531c1e379d424a524944312fff83b70f69eea55c13ccfda7c69ce791b15bf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fb65bc2447d6cf82a8ceecabb0d59d340c70c22ef878034e3a6ef2bf9eefcbf5b27951d6e838c740487c8dc777ef855bd6b2b7c5dd09ca32be82312704a27d3b80930d21a3a8549fab134c7c671e4372f612e9419e9d447486c5201e232f365f2846804a8735872deb7578d34e923577069b24ebac0032ee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h84bf13bb6b79f6549b401d19690396fd4232fd73044f31367acf6be04a2ef6453e76c1e7da436a4012ac67ad4e43263bd9d401dfcba9adebb23a1f2e26b4dfbd80777518a43ff9eac5ef81db23fa46fc5619df8e5ebc5bab09c316d2fc33782d6fc28f8129c36ad2a45b19fb9fd9f77676a0802f9a9f994a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7b8ccf75c81ece692ce6dd4fe011758c2f5e02a1460726c138d0b660f0fe9b5b8e1da038972f91008311b18a55d0adc0c018cca01cbed65e091e7f1555dfb4c068c1b503f53c99e30dac5df1ad76043ec5c929c8e1966453585967144ea8fc6e810cd8cbe31634777aa5ea01336fd68ed2601487f0d14e8f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14d41391a9cd966a97e39d6657b0e6c18d135416d29677dcd0f58a2c9caf2c8dd696e1dcbf6a3e48044aa582cb23167dc3862da893d162cf5a79ab587416f88681e1eca258679f01839271ac5db7bdce9a2d9c599718f6656f20d24068468e8fff54ee5ab7947c8dbf047224cf6ad321e6ebd27d0a16d057;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ee0ec13c7f3cdd8c9fe68758dea91eb5d40f3e21f47feebaf5963283dc11ab95e24566823e2735a8e83767172cf4869e6e1ad6f960f6d122d9e7dd700f4290602e0e8e436d79c64211d4a16496255efd6c883a0be51979c12694ae96d8002be7129ccc70fb53422ef9d00a76a1299b37370503aa64f461a0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h168840e5b6d34bb8ac8271442c9a548529426b075aefde8cf38612529585bcbfb27eeaa71aa20e668758e24977678d6c40ef4108efd06c87fe54134fd12cb99691c97506d0215479b57516106320140fc9868a072799ae8f880dce76deab80a429d0dd4e43f42c8d372d022ec71baf3dc68c6c75343068d24;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1591b0438da025995371e85bca6886c59cca5a9f879edd9c37984a366b21b1e70e589a3b6def0524cf628bebfb51d2a2c30f57e570bb794da7cce0ba4e74f86d404ac3ccd343d1b07dbf3a864fb9003bb011050fc1f607d3f1d1a35c6b1624e6bec539e80b77ce7d72b8c4da41d9cdc152d1c00dcdcd2fa80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1cbb4952213b1d496d2e12689b62f7fb547eb3a1d32733af9bdcfe4359098a727e7c9a73ff0802f4e5e993dcc9f0c8048c257e2cd69b76c5c3c41476ecc767c6dd503a3e9c0a236993f7d0c4751ce5f54ddce0f7019d0655fca787b3b49d1854cd5f2783025669322ba22b8dec9c7ccb97be126be46a1fe33;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h7814d0b3460f121eb40fcc7a082b1b34da876cab76d6734fed8fe433fba8b64a6097e43898117d7a8648510ba23029163475f7feea47b1f069f1091300fedd5486ae5034faf26c826849c8cf8ea714b92bcdbbbebf1b53e06890f6c3d08775a6a347c0cf0b48a2b1c641eb1933a293ef2a96ed127880bc77;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h153b1fa00dc76b131b87687198321fa793206d44dae40ed63d35f07184b3f9dffbf6f07c335178e0a60908338f6bc18affdcd1de8b9f769d1e2cf10c31555a7e9e256b78fc5e701868878a8a02dd429c8368489caf2d214066855c6b159d6785708a073e57082d34c0fa211f995773392d4ebf8ac3eea5b80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h53530a77921cc9f9f0076c2bb659738de5dceb71e1930540764f3aa825e344a9c36b1dd8918ce44b28e31ca4a29962156205cab508b8cc757ab3aba3efc223717a91294eb28c510bf21654427325537666335e16b1706a395dde9d9899d3470100d505ce79e305ac2c4ee759d367972c2ecfa4b38e552133;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8124af58a5e4f8b2ea47e47f167381d3c371add0928d6844e355ff758c302733b599476370041930c6dbce68ede8b4b66d064db3aca6f734b3150e225f26f1e56a27196cac822d47d382571ecfb6e8c893c4241a5265adf2fbaeb81bb07f489adc3cc65ee48e78b084cb9642b1a2ea9a757611035d65af90;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14008243f205551e89be145f2b71c959fe508e7921ab33261db1bef4ef2ad4a194f2b170ed5540d27dd20a08b80e2e78acc1e15aaaa6b7660887c9e618c01492b2c05bad68a66ec1c783bd40302b84de45cefeb3dafaf75af10df347a07e70dc3a9907aaf2e75b1b6de84fba4a0674e444d7b36373b0d4ec0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2562b3fa06e67a06061c93a4aab483eb340d48890492f4ed95338fae42e208a4debd18c21085fd09f0beb58d13cf8e8560c9e5b955d8a5c13ec0a0ae2a1ae657fc99ee4124aea5e1dd7ed654748ce343fe3eba6017a6171350e69c61f97fd0b215b3da717c817fdd59fa9d7556ca89333e5e6fb32a091e9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f4b260f41fd47bce7d46f66a30b802a8918ed3e8641e37a439094bfdaf0e821bd3181a6b469b64c87fe05a223a149957d3e0a00e2a570aa7d4b8eafcf532f9ed955c8d7e097a6105c868095e8001597289cf713735909f96a37201987bc2f89421a41c74ace244fdaf5525fb622a6ac39a0054f576630e98;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h68985073b65573c536b9a96188278ae7f2c3f4c71ac00f20c53d2567365575a4d2774038a93c316a3032d659131eebc44713cde3babe2740eedf1a9ae52fd5d894361b3f2bb87ff213d84ac034dc5abb6ed3e387ce8fac952dbbe804f4d19e8a61b52ec994500cddb01d84c1627d5e39ef236cfab20cb665;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c094e186b36d78f6b98ca0dd4338b2cc19c912750ec82a00bd208135d4b339952afa5e14c7ebf663c2788734cacab89d078934747c840d6fcba5b140f74ce5ffa7a5023d4a166645570b4a2c1745a091e053fca6222cf9f808a40d1e717d6e525ad4626d06076c8449bdc95ca34d810df17489c0cd8c127;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h473508635adf57e4b8d2e77a85c16bb18976d894891df9c6d62ce01d03c45ad2bb007ba8e92926ee2df650ca773639fa8516cf433b942402f63f08467b12b100029960cedc57bb031a5a9a6d75e2e54561c8ada29783acbd9adab47a7270e8eda890c114edbe709121f412c427ec9d752c9707bdbf202aaa;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1aef12fb5e83446c9a1d8c3db3a460eb8087ec2b1a2279c42dee0fbd59a57eb07934e3dd27e1428105eac01cdd86f2efcb73adfd94513be8b26ab90b3cd24effad5a6f1fd6f46eddb73fea58fe4d200eecadc19d2922f1f718ed2e0d09a9c70beda750b8897fd23d0e34f22198d7a68daf892cc32d6ada432;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h69452e7d3687a48ce31a571eff7fe0ec5538f50763482ba3dbcdddab7a540e46241cb49785f7d017e8d92b5b25cc57c98bd781d949095a74f3419405aaa599206810844c65bcc4c9c730a70cb2e9865fc762f3240638fd451d9b5258e6caf80de89a9345530f9536ce8bbc2a83d8e07f42cb0f4cafea50a4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h175978840849ad918bfada550410f2bd392ec6bb31dd7c6b8717cb7e24a8a2b5fdd453800f891acd11e49691b8439a512f71328fbdbf16ed18afb9e9c4f9680c06315d7a35eab839d03b1a5fb13ef3742f4a3f31012eddbc83573a093c0e0aa9a87475481afc3d414884e7f241176940ec59abed483ab727f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1148aadaf88f5e5674886709896441219beb0523bff38cd010c4a841e008ab808d2051292566b044db5de0b68091e7d6daea0170f322c706748668079397b4ccba92cd9baf0c0bf63530101ff95c0e6c41922577bbe2f25b28b200cb28a1d4da1acc3080562a226bb8f6bc4ea49d04bb6204d030d1f7f99a3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15352de0d9c9c94696ccad7ac2b779a1bc243f0fbb5db1a448de397d690425726dac3a74d15de48783e3364bb7b3f5fa1abece7f3e638b2452d321534d3b25a310efe5bc214b79726ab73754568bf1839fda5d877b4d961d8f4ffc243c78051c244610eacf3c56f66485e3289fa9f8287021d85643699db33;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19dd56361627ff39b271fbb2a5e0e6d07a0947d816e41d7238675a052bc081dfcb66a27d9fa7515f8ff1c35c255a778c095736aef46f2d97f3db8bb24937ec868a8656087aa45c58af9d92e2c264ca8d20e9d9593030c99b3231a8e5d6b6a7c39665f809aa120af685fa3a6d981eb42e1c75485cdfd912b5c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h558325c5f8701dfe2340301f7ee25f6804bab8dbc21c276bc13217ef2bd2aa93e937691d477f5ffe74a46f9c573d355cb6d384c03797f2e13f0477b906ca4b3f6a86351b1e9b61c902995200769fc99c1b12d3a4645e849dba9314a493f776920b22bb9a7b5973f20aee07b3785882538deeed969f95f984;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bb11d25e2fdd59ff9f1e316aed97f147dcfadafa20b0ddfe9e95dd3f24028ccc705d9d96808b4d149d416dd2cdce366edd4d45ad1880014f0253d679d9bc9d01e4c4fc7f41c0d569fbf476514ccfc158b90f4307798d7d71823618ed2b8d04ad9e19ad7c893b05f9a17ae8666b4acba1cca0a4566975c4c8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1876d4d0bc3d7b449a7bea61415f341e21d29ec8442210b88ec034b532854011f3bbddf298aef36ee0fc179137764fc37f81440c2e3629864560698772026da926ee366a59d2e1bfd3ef15b0c411a6e6a3d0280450090e2ee0493bd611c1e178f6fed618fcb3d196a61086e7b238837249317247c73281a72;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ee0ca8bc9e3f358134ab494444e8b7d433514e2c19eb365bca8b660194c4c679dbd0c959b1274c37ac14a3cc7190dcf9c33a38565a41d1821407e5bfa349447c05a2624f9b2851e0c5338bbc9b83c0fa41a6d5f4e67e406b99aa862ba871a1bbd2a864fdd711d8802c0790fd2aa284bece473f28eab3d695;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h23016330dbadbf9a35eec2e798043028f4a354ef8a291c7d4ca03fbacaa604d7c1648d1b8f4b8234a68d40f4b9041087e2f8bd86a41aeb848d06d26fbd0d18aaec34909d5385e16b045ee8a06e41b8cca3784260547232dcc74d52aefe1b51d6f92ceb558876f7d033cc12f7e41c05e418a30b2252c36891;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h146b57d89583acee62d4bf49dd69485cd4a2563e101c1778915438c3f179c70ac31147c1803cb753d45ac3aebf94c8b192fb908789f99f1e5aa56b594cadb2ae2c3b7c11e5952a020d2b3ae943fe44b65e5c7d49138383bbca32ac9f3ea27a577584c9ef21b446dd71a59fc8a16ddf9dd5fb4bbf0c49b9993;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c9681fc7446f3989cd8882e96cd914bc4f0c57e0492409a2876ffc64596bfed3e903f85f7bd990ad7df3d457bbc6fb33a24cbf5cbcd008eeaee1731251689f248ad0c03b3ff8193fd8c6058fc0195a85b17810de6f07e39fb3e23a7416d41c2bd6fa9ab72d0d944412a2e54342a9c6684889f9864dcf1915;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f08a180a8d206eba29bafb3d226d27ba01ead405338a5d00defe86ced1e0e2f00035ae4774fcd522acc2ed85ca974cc1b38aa29aad0bce1c2d3ca013b94202265c2696f49f6790f97ee1cb1950b06608e5fd22d60834ced8d0d6fd8af29fd7ba0ba18c183833340f57956ac096171af301a3cf90425ced6e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h5d6ced987e8ec8d461ec1084d23c22549856855927f2640d5222190409b9f112510e00d7de854ec0850f2cd53706214280848dd8310c38f25799d7b93f984f0bec407fbac2dd12dd6dba267921aa2f15135366219f2c1633140b228bd21d49a25246f77dbf4f0f46ff700c46b9ffbe8fff970f888abb16db;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f0487c941daf64c8adff3290a1de18c7a482a7ea9cbf1c7a06c10c5cf67384f4e4ed2dc7fee138f101496156ddf65c7c2e221a7d8faa1c171c972469966701e4fbdd1e71bac9c0dd5b5afcafe37d6196adef1d397c2dc80b711a383427759758f217f4430356dbba8cb5927b762477e44fc9b7a38f176ec2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf23b4dacdac33b0f921c947bc8e7673b6a2b948030b30c55df2309cd7a48b4403ed92a3bc8bd2ae29ccf8d1d8d11b1bfb698f39b74b48b3ee7dcd10b6e4f5e15804b76ddcf4142765ba28990e41380c16a6fb55f82fc6c692aa6700aeffa13eea8f407f29fbd440d54fd0cfcddf7bce5e60c294e1e9e12e7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a9366b4eedf24c6d252b46d7bfd66748cc7c95317ea791c96a13ef9ef392dbdd228274a451a63eb78ba51b3925918668991ef2eaedd2c727bee854688527f43c1bc4a5d10ff686a5644af565058c90b946e44f1d7e611e1f75c89b44dc42968126925ce71ccf80703ff02a5e0caba950cce672084c493622;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a7ca1b1191a2962e6ea9e88a2f69349ec19cfc3a7b4bb30d689d2c922eeeaa7edbffc24f66da4123621c7418b19802a9cf0fd0d463b26a0803cd9d683c37f208896ec365d2d9dc21d30e9957b7bda0aeaa330bf65a1d414280cfab607734741047dbdd775f3e4dfe86a9fa590e8f586bc1a0037cc1e4fdf2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13f6bb9b602e504d994ee119fa158fa2bd2322dc69437802335fd620bb6d47851a05c9cb2db5c640b10c4df54194000233dc60e499230591a682f71c0028a2aa4b0eb15195f9c5a65f53be872ded7657855d9a4218c431b19eb1f52f452056cff824870e6259b0ce92573b4156b5b3e31eea7089e09cdd751;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'haa780726a8dc71c8fcbe4c3db7ab8aa87df80d5f4c203bd5026ef9a2ba999fe496b85d50af4233b09903132f486ae6e8e0169a3554ffcff3c6893b5fa17dfa862ecc3d85f99aa6ac2584b35ce41d547ef529b7ee6cdbb7744a74e0b09b7c01ee536febf2f547cd6d2753dedde84e6781c920ead9a155b95a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb225856361f63e4e0ef3b0216c9ed77919d66f6879e28e9e032318b40db4f3f1701f6c388548ea07912c8787109964d87a8dd31640b59e1b37aba84297e0b316d784b2cce24dffeecd5c52640c53604d03aede757c64a7e7538abde848bde4e7e29f6463c14180415e0273ea7f6697c385fa575538c21b45;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbb00c5905d47bdf9b782d63e3be825be66a5c137b2379da293847ab5044b4c349afd825c73536a7f161f59a34dc97fcc5400f3ded25553cf91bbdb34126ad8f3c6280926f5b540677e37b835401632ecb2c0e79e1783d84a994d0fefbd168b3ef7f62431bda0f595b2fcf43600ec59db83e1bdb7c2cd0052;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19504b4a02c6273ce8074c8627406114f168dbb81b7a34e229c38494ff94d948edf873de2970647e96d139d83c5a194dceed0c46b2a9198d1fd1fc01da55d8836b7aa4f13234cd9152330a40d64cc5badb62c7751321d9acaf945cfa65732bd3363632394e62115bf1a242dc21621226ff0b14cd530f5f247;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h199ad7eaa2ea4f3bab1b8859dda07b0a60639cc7a84d4bdec18bb36ebfb8ecf8dac5c74da0d5c2a9a9dd5a8cc5bb28dc2874634b8d1fd2d919dc298b2e2bcd15d9435b96783742a9027e32c2e1f9886fd68dcd2678b3a61e9750fd0397a4b0c1e486290a24410b19cdf080876df2ab4c5310e63cd8dec4c61;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h766168c3d960221eed55ab909a32947e07909435d76d3f25a0472049e176d55757dd70a67d234333101a902a31dd5abcb49e4620dd7bb45617fc69a5642ffd62aa84fae652b01287d3df4f7631fb54e403776a595b47fc8d671c69a493fde855e9440e9976d777b11762aca55b297fa5027a9c8267b415b0;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1ac46d6c4d10a759db2448a8c9e60852e43bf8e6985d4e487ee8d50cddef52ef578e99d6deab7e615b8696f5aad1ee61023260feb888327bb7a71cb2c5fe6b306bde9341138983a337b37f29f713e22a7f7b266aae3782ab23db77d9d3a4201fbc5e5dd7581ef8129dab82ca42c921f0527a25b64410caf;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc6ef3a4ed9d83a482df73800053330ca0ae153b11ac799e65241ee3836810c683c7fc676720710943f070745e672c27be373c147a2756196ccf9c744fa13038e9b23ea7df92490afc2d477e48b24eaa3a35169e764aafa8c35dae79d254e8fc0ae8bf49e6768b57b4968d1466822af4631865b53310bf2d8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f1df30b632f98a7e08dfa3c992f4d30645a7c484a92efc94e4c5f5706bfb1b672c52080c86785b5446ecdf4b76046e2c58e37ffb874463642db4a501a2fd1832b94565a356080e99f9ba9bd514a274e1565d34588eb3f4451b334dbec038e3ace023a2dbc1c6b15de26baf928964ab75b8432f6fe5daada4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19c98562f081d3f0aad0193bcd87f0ed5810e3328327f47055a754eb0a4bbaef532c43acb70d531fcfefd9f7f0dac1d3c9b81c911e068ec2304c414ae4d222eb225d29ea116005cd1d5175a7d0769690810ae3b1f1e1ffd96c148916b66f4b097ffb4444b63b2d7804a3cb6c3903818492f5b404f254f3aa2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h61343618637f6c4d162c7a25509ddd5a5c23adca2ff0f46271893e6cae378474231f7b2818c10f657d915d0af1eec52a712b418fbd6070d67f057338e63530915f2006f093a0cb74508e2236533e9cad6d05759111b89b131bef040c43969cf01f272df3780e1a22cea6fb2e48d513e7f812f8b609f6f9e6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f0ec1a95ec006d7c953bb06025e19ea0f1e83c61dc48d72457966ed42cc73a2ec674a7487a2a089daac5d268c96fd4f14852b730db5023920e583d1cf68a3d385e29438fb9ccd607752cdf5813e16f332ed0c85d43e642152a161bd31c846bb9b686cb91d09d6edbc21751c2e06ad6df3097b9e9bc277107;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bbd963271ae05445524ba93651429370d0901269e9c60b03f366631b01c72d548943c112ad0d0792db361e2d0d4799cfaf0e48d4f08c2c53043ce7395833e77e6363452c62eb7dc4ddc4f0af88c1e6b49c7ac13c1863f474d85b9fa35c15e09d09a93ac60036b62e0ab544d78343d121227bc93bdac289a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc0859a97a73ff196bea6b15edb3fffa1718329975fb83f5b33948d2593ec1ba0f4e8eb6f95e50ff820bf029d27428880338f73b675a07b6e8d274d81cf77548a3300c120f65b7ab2d65be395e40c2eb539c89ed76d30439d3fdc01ba2fdd10b25dc8ba0f8b8249d3d3c89aa1b1d02ab4104cc283ac23002e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h746bd96bb1eaa7fbc78f00c831bc7f9bd172980f9d2e6c9b01c01e3922e0c0a6432511afa296f824d1bc7c9e73471a2dbbe0729e1303255a1d56652a54b2b27bd14de62fd9fc70f4bfd18b2299c117c09a2fe51bbf934e40c6e26db5c92ccc58c6ba4d87f50a478ace27b43e4816f26d1bbbe5a6452d3ce3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h143dfbc2bb6f9ca47113fa1274ed28cc2a1833b56ae2627afb49baeee39aa0fb4fb306f743a6e8b24e5caace1d426b15730410607b4b5bba4fac079f5a1baec84315f9627b5eb70bb2fc4a87f68ece41fba5c98faa92c0cb6e1c1c98be5622b7baf047c4846b9382bc7d10bc1c1907b0e1ec3cc20922c8592;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17cc9ef6822f11b67af94a03ce1e729d058f956ebdb8ead13e216dfca98f0866c213b7075d735dfeb69880d39db27279f44e04f6fd420952b4e853c1f9e07012a6979dad85f4c7d369890468727c547dda4b8aab25921f87aedeb9b50ce49cf02bbbd4b1043847bee02409073b2eaaf396d1604821c44db1e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc471c5243fd262d989f4e764143f41a44a258671be6ed96d9a598ff75313e85619417670e67dd36545dacc805eecb9659474254f05b6c8ce16607fd449c2a9ca784e0d65facd263fe0bfdcdfe69a1324e738e603525da3e632eec8f7fb1150b3557e642b490c13e1b3bb646747f20e1e8d4feb23001ff09a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1b99a3d0e5aca3a930a647907519aa18ed9563dfcf1143bed6e7f80ea879f57520c2cacef18c25c004fa03a3d93593299b468e65e630b1f063109cfef3735dc169d4bd63f3346615b46a207c344b219c84dfc093ad74cb26ff8e7313010dfc2368ae65d0ee905db0618090c352f1695e3e1a19113e38c1dd6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'habaa90dc4cc0a76f857f71b27aa5c1e7cc1fc6d2615c1b51c663a5f510fca1dfff09f588084d4e558de6c511681cefd3fd87d1b0cda5edbdf298a5917849ed8e355d0635f0ba205facd7205919c3319e545397fdeed451ee26dcc8a5515090483d385296c62505765a8cefe84908972dbd9ed97f63049fce;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h104fcbd5e130c6fb453589656eddc6bd6f6da68ef9c41caae63728b86abe8f826ff586c73295c506b6d3657be4006dfd5a257775b6c3bfe510b1bf939eedc4b0b2aaef8ebd8a9a05ff3f8cc631bb5b4fe46eb2be11b4397347caff2cc1f75f911ccd94018ace90db19c6765975263d124f471b14f96258bf7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fae9b01f66ece50c11c8952327ad394f168f74e86d79ddc26099fc03faddece5f8568317087466da76fc052d9902b7070361b43542d5a8b95c6a602b1ac186bc9da23e730646017a09fd2f4660c18dcd9007638cbac3ca7a88bed8f8a4ebe5087a4e1da8a5b2c93f3ee4e83c2e5c1b4c9b2fd4520999c835;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ba364c97774c97c08eb28b2c50f38c4738de89345d6a2783bd11c7b07ab9ee0e9cc81817c685d5f8ce466236a7947418e6c80c7abe9b1fdac9af2225d861a73a0a31af201515f65a301dd401bcd1828283f99685fe3eb0cdc798b24381c1bf830641761b0cbc3d55a8d9ca08e3ab3381ea75b8a7cf60d52a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h74bfc636e3689b68dfa547f8f5ee754c81c431ee6bc09268eea94d2af49263de187b32c3bc3f4fa73b0d063eb91d9d1b17cfc357ebcc7f2023e9bfa9b6016587fcd005ef31a68e7af28c8478e6b366d7290987032190e219f95c105b470d5f17777e1670b35eac98f6f6aba46119f7cd1b67ca835517d1fd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h158aba4ce53fade9aca77b6eb163df3ca5bfca827525fcaba90def98e9bfb561fbb78ca677d02208076f9c7331e5819d9f50a49059df20b88ec5e9715a087be32e5df64101b3a5163df4417087d9f9632843c45d628391a3892e2c4213da327fdaffe3c464b1d807f884575b4f1b9fd477f2d69db6f51fee;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbca4a0a42df04d5c340a3bfb457df3d515c39508262bdfaa61efd9abe1aaa6760161bfc2dfd6d3868531f975376869da19cbdd80e85eff6dfeff2db096ebd574baa99a9876f89ba2f2a0ec4dd7cda6fba050925ad15357974309ee0e10017ee6c62d69255299e0d2ef53fb90f445c41e8f029cbf7c49c319;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e4b500f469b880a86ca4e2b2a0d6fde04d90bd0eec38f4460ce13b94d7b46f2ba3873106979942bae170bca4bd0f2765c7e67437f743bcd3a3626088a379dd6555354661c3d1afc46b4c7588b102299de222ad521ca5773b1aeba35497c50200f7753e19cfad05e8aa34e54b215eaf20469b5547724fcd4d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h6fe9e6502cff469bf2e887150e5f7548d0c0a781baf14c39df4f1cdd8a76d347f31d9097357cfe942e36674c51e3ada0d20f8220411ea10b0bb312c2dc0d7f47b2800ff4c0e4bc92c1aab11407e347cd589a39643cbec592935e985c87d32352f975d5a9f71300fda3f383b72fcb68cda59a9462204084bd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2dab831f3b3be3498e01913ce2a2d9492e065020d65bc82aa123fc4424bc0671fdaaac4c167112abb2bc4f7abcb65c711ccd92afb527da03a162d1116289e118687ddd7352c569247c83fa91a37f1750858d8522cb1406e3ffe9c80fe85acfff34c4914eb733b739d81624134f6633b325625364dfcaa501;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18fd65159b6f16a89133199c5aad796761ab0ce6a6ccc8ea4e04e9095134d44fde6165ec63c2c5de3face7da59c7068f977a10730af74d04904ef219a9bddc9b2c3ecc57e915d36b7d3102c43d5104f2090a5714fa43f26d20e562a2b4d57325fc5f7602129a611bc3bbf1203fda1d0216e38ad64b9349462;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3d4d92caccb850cc03c898cbe68ed6cbe3d1df493757ce480fb552dfd397e1a9a3bfb7e1514ddf19e0dad3b584d41a67aca3889589c4b6ab4ae62084c266e4372a0557a6ef555a970b172460238fdd273249ac79df397c0c16cccb5fa3ff79bf09214447593e1058887c47c45b9b9035e7f82ecb99e5ca24;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a21c3b3b3d5140377fa7b654fa82da9e5d1b1343e5710e1605d60cbe1b7b04237f2893a23c003025eb740d9e7617378150cbf63d08da3961f5a13f0439cd74c5b8a06120ec4b1b8067af2b2d618908de28124fa01c43dfe44f7418b5ec3a006656e3ecb9cf1987d78a1b5ff56c9c47402f51a1d1b8355fa5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h104cc06fd39ae601b7b744d0f63dde1a6ade7fad02040efab87a1106e155a8543e06c31809d590ea6ffcc46b4c9ad51951937e5f7065d9c33c3986165b24499f13dec5f9ae7d4fb19edc3a3a963d537e498f37b3810b59bed43391f93a64a12f0dec38d7c3800ad3a346eaff49630f9cd01fa76d2fd599421;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf2d65a17b3ef405f242fcab630fb3ed0492c37f3503d58d1081de4a7bd1889fcd17a8a2ec34420510e6dd3c3cc21a572a89156c2b654b349c9872a3b5b4435ceb2175e7bed2933fe015a74d4aef99903ce255ba9ef6c9de206bc3adceb87a08bffa5237d71cf5f06a5a79b2c77267ef498c3e77c1283e41d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15d0c2df892142803da28a8818288de61ac362fb408f321594cce8763148d73eba1810438b5ebcca0c17cf83eb54bbb4390c37c17350c77bfa96bb5569bb0f3bd0683e44b457c99468fcd5e367e275443b0f01d12524fe3bfedbf3b97c2257538c48fe60906126a1de7aa433ecd473b4ac09463ff8e13d446;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h115cbac861e43bd55a8d0b1c8a500cc00992b3ff43acd9f529ac994709dfc25678b202e42be0472cd5dcf34608c9863a614edada755ea81911787a20dad82e07785154e33c761a35bbf3867af53a1791f8e5ab14eb7be77d55077b3c56ea2073be8c7e7f8039007e369eb29af5cc94d57eef247cb03349ac3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1d52b828f3121f976d827024682f4da4337e818b86d4ecee807c11f08d6202a86edf4a0784b3a936fc8fe9c0cf10a491883b39ce296edb2cfe7bb264da80207a871ce53afbb9aa0dc2df2b400cbfa6a41ac8e1fec90b245db317fbf087507f76f387f52677d966aa77c3c2c8ca665dc267bd71a1e6773380a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h16d4a29a8f49a5522ba472d9e74ec9377f250ccce724b7b9f678d6bc172e2275a512476a3d343cdf2f21001ee4876228eaa417b740ed0e9133613cbe8b3f5092bfd7d644ed19725db4b5450793637458d051904851871cf9a59303e346ce4c994cab6043d278d3be837a3d72abcbbc854b6181b0dbc7a8c1b;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1af165314bf084d2632311074731951b7796d4b0e31154865bf9e15f8725e3d33523f28f9bf30f3b113c1f04fb721f6fad57aceac5c58740b96ca38f2fc11c1b4a0acf596987bf26814edc37f70b20ac8eff14d3fd91a5c19d2b23bfdf5e235397af2142242d9f728699828ab738f7d90ef9b9193630022f7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hc1b746fa546a43465cc2c86bbcfacb91a0d4a3711d7aa0891a39310254113e695ea165e858b53f92c653e9d6ac7e339ea743dae95d239dabbeda4f2ceeb3e109e6393c05756c6fdd7b21e4bee18a4511e7105040b7c636713f32fce3ff905de2bfc57149b65f4db7d2f5415224326b8b6c2009eef98d8f29;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4c779ff0eeef054987d862486922db477f3d2ca53d6bc9ad8302e3f179c06ff24593ee45d04466ebe0c7db89ee4961db70c038080b051d67af3e73261d34326baae448de6cc51a092a21ed189fabd835bd3d2f9466baf437f5307aece7cf3c23aadc81fdb842b2d934a83cf6d3662461b01d4e27abd675e2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hec4aeabee3813bb1bcd48d57f9ecff2a9b347019612bbe9f06dd38b9b970cb0720e5f60eec7eb36725ab8087616be19b0f61f51d63da401586a6c918212f002363525b40ae5240b0d0ee34e3bbc352928cbdc90f3e79b34bb15f4502ed25385311350270d0604b97f0414eee3881e460cc0a7ee6249c04fc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1df47571a108a416cfda284d8cde6f5d46c0bb824e2a55d722a786c3e70ad95bf7370474628f70a291eb370f4ddc596f6cbadcd6a97bd123be75d57319de2cd5f86c8ddf153511c2c4450987f31f95d950a451fbd8646af7b404df830784eb7a296c6812fecb43c395e02bf092ad1ce224d8cbdfae681a89d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dba6fb46e4fb02a5b241f1ed5faa71ce63699f9887eadde9bacfdc792103959e072efe0b50079c3d7ad10f71bd8c423d71d4affd572131b8d60eb7b62f779442ebca4bbfb423b75dc28c7c45d4f4f085030dd3bd19740d3c5becdfe06bbcd436a614108859dc313368723254225189df94dd1f42edfc4d12;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10838f5b9dae79415bd1fb13d6ac6a6699c5464ab5d2b73ec656ded810caeccebed979d0443e05b87812a175bc2b5bf0bff42ebbeb4b0a645b02e79664a98d0995fe9e9bbb127394171cc411fa4abd87b91b2da7178ca958693607d7dbb77ab5cdd4994e1d3969f69ae96b9c06f2edac25a217e8f20911bca;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h179da7d7a8c3f0aa8b3a5bf0517c7d767eba0c70172cdb6892647be66a61ba895ca0808e3733d171b530ae00022b11f9a6c9b6479b52bb95bc47283c29eca5ca5a46e666d068be2b8a7f407a7b70ed86d13bb4e3d8bf0e12283a2c16349d0a1aec60482a89ab20daebdfb148d3da89ae54ce2ee6dc6200ede;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h138180fe2a9d501ab983464681c62e711200f1c4a6b162b8b4233579c8d989791b28f975cbe542305bac2940f618071934b1d5c1b53e1edf8f434eb33cc0d9c94c2fad69d9ce61c2b856af64de3cfd85043a84b1cd457461efbf5b26c5a8ed23d005a2709ed486aa27f8c7a3ea9b6190bd1051d5e8e603402;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h83a8cd03910e740f74d0634a24a8ba8c60b0349399dfb2ba9e568aaa9d05109f63bd31d3c54f14321693af778e25f69d666e936670a16f7ea71ea8862c4687f6f0e14966b03193ed26636170e25e589186b27aa64a4ba18d05930efba97ba679c0e9007648e1dab4da884a262255eb03d017323026f14548;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c53a8cc7e6e606ca8e484ca0c2e9c8627786d21cb8fd3dd07272230ae86a0a3ba4ffe3fcc4575e3902e303d77774ee4d4a0b12c4f2367f4eafe58b3d0dde77ad68fea17f4c9fc1700536ff8538fb42d1bbafda287a549d2ef2e4fecd41625406b1d6fee23cc5e942c913ba8e4755df52fc89c54908422edd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3964971372d0f77fbe2a51629e861c8004d23fb291407ea8c2f6001c12760d683f92bbf55f7141c6c9bc94f6936a50d2e8f22fe73998d6648fee47ec2035b8d6c1333d0a6435cadd1c11f9780fd7bad59148a4159e1c2346fb7e4b258fcad9307365d88c2519a41fa4a58765722f3d90fa9991fb35764f9a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h137df3468b9e87288652eef912e16c8e1e5c7aa602266bfb7d5d213b080c72a12df73a9863b4fb00bc73d5e13d9fb48cb1512c318858937c3bedbbc4f6a5a0e20a412c7250a578b8aac9c882073f43d9c34653932bc0f85dc2fe8c6e5bb6b51f4384175a5a74b67a04637389009c0aab9e3c3f4c18218ba90;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f261a692ca2e1df023d90b947f3201e0376005c4e1d80d074a188a18f0b3a5fc3509648e940ea5347b80ad1fdc3fcab1abe7c4e5ff47908f3b54e8711dc293ad734ee52b7e6fcc69739706410aaf75b5beae82084df9f3b209c9e7fe1ae922907f9467da14495f759c50548cd75b611b83728d265d20a0ad;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hafa6ac81dbf29033b5f455e09b378cec3f2d4e10d01467e475ed493a4d574d5697f2c4be4d4941298a347f2fd9f06741241459f6c4279efa201c0029a8431ccda9d6b108fad2ef936727d5e321952d8d80ed1d60495dcce8c4b6710b3559a00db3025ef663ca39a3fa37ce0cef883380ef04f0a62596e324;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h195ee0dd06523ca1b83521030f33c29ab2f37c4b53c874b237e429b9cc6207d156c366c71120458deaeb23e84f890e921f8931dff81b2f93af08f71761245b92158e64c3db0bb8a96c1d8a49ffee254c858106f49455218380187a714301655c3f70474b72e7e21dd4ad640b6b51ca576f16993a85c9de213;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h535229c1a7dc8ae5a8d75d086f22dbfbf02a49f1e1814806ab0b2a39e6bccde7d3a4f96e91eb10d0bccea9fa50a7251899a2e28dbeb95563354584306d30df47aad7873d6cde47f71a243a29920e1ddc558ea120d6c33bc636bac82d2280305e3511f54d0e50e25e8f9b5dbb52cc7f32ada6b426dc250bbd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h24e51724de992f40fb83771fb37e76556ff8ace37621fbce2700136bd5aabc0168c5a840278cc14ea7703e76e9fbfd9df2382f228f2419f4abca4b70fc9aaa868139881d64e11288499bf6596a9c02b97ff1e95995d5d7f85a91bfca80c92a018b1ff33e3d2311dbe17691bfe3e933c23ccb82f2bc9bdcab;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f1aa2df3fa26fd7dc503c3b46cd6a4fcc1eb831f9bc85d287a513c4eee26cc823bc53ff7495066a37c96894e1664ac330dfe3aea20e4af6be2f916d0395756d4e80648d2ae4ce3193292f70952416e9416c5d0e8c72b579b57d6756da2a8205b77936dc397f246a01d22142a2dec65cab95c2d39538a10de;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8a0fd72f4422b8018b044ab640ead11d8df62194e8b022cb61c5ef567a4cc3b3d5b10e8af20d69fa3099bad51d2d5bf9c5ab2e3b5afca19c5bf9efdd1516e98963507eb08e8fdfaecd710778abb5486a396db88f87facf7942eab3e57307a4f0b39c32492120a044cadd4933c9025b41b983cd33cb5df3ac;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hef13ea76dd391b722a5829dc9a7faa97788ac8f473e413f80ef3935bfed4cca909ee860aaa47fd13be771f8b0fed62fe51db20ecf1e25399c07f1f8cb104a50daf08aacf23a4818cc5a6dd943cf2c4144beb1e77a21e402adbb14cd53c731267079ef8f889015d8771b02ce830fb65a57a0b7744417054ef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a45503856d59c3a7e04b369a18c3ccc64d2a4d5853d76abaaceb73521f3cd8e4af804edbde5a0356567e1fdbd2fedbcea7951ff59f37fd08fbdb097a4ecdd554e71248c4b5f86eabf4557c2c30eed55decd721c804973ea4f0c88be74edf6fba2eea36d9c5e29fc655f7e27cfd20285136494687db4fbaf6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h84e03705899fcc7de2419506d10e68d273eb55b9f7ee56b3f8784766c44eb40c498fc62708b965e7b0edf50adc54cbcb58428bf1554c495c1234d936e5e307b0dcafe786144bc332bee695f9847e0aaecf89a9539527250fc5deb339b60f82bba05df9b1da1b7ad7c151493c5695dddbafbf5194b4431918;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10a1e6eabf36cd2edbec2f435e55373615ef68af3b5963b9ba72285c7720bc54e020a1e9244d1f65f10cb629114aac54beaadf3fd427948323913122b9517b3ceb69112d08b42052187d8917c01306c81b959381bbd3093dcd24ecd9ee84769b4cd40fdd509926accd1e554d2ca25e4e1b4b8a5be6fbef94c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h17132ed60cbb8ebe3d944bbb5be3615978ebf501dad4f8dbc74e54bff951e7cf6ee8585be15a5cbae0afa16161cfd566ad316086b0e16ad50d9e091b6759723a3bfca195dffbc70aa7ceae8a53a68b0672d3d2c1151243d144c87f071d94b8e4a0a31054f0ca0c694cde59998fc29c8727ce4e36cca88fdf8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1695e4d2146fca6cd98b3e774babc06bdecd7b78bd963b218887fdf90b4278c66124ca47ca9dce72584cf86a94e9cc575f90d78be7ce306048b55ed24dd104ce0a8935cc6f3ea59db9e95b81e716e2786ae3e21ca19657aa8d132b4b8739ef9b675e7785539ca459e5fdf4462e64f7836bdbc80a73c3fefe4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8b9cb133cf17ba89430c8760915e622f98bd7b873dd33bd9e417fad05b80d358cd0d53ebb2ae8eff4d2770dbda98609ee9a71a300cb91caefab8c8e490c2bcdefb27a0a76c80b39100efd19522c2a694063af9a8afb1261a6b59368f3b12a7e04923ebc085aac9db43c9aca9025765c777b4b0d6ad5a7ed8;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1ded88aaf42d61cdad1148c7fad8f7a5a9bd9fae750f91d8fa8733872142314b38177933f69a6fdd2a559219f1972f96a4f575e62e643e0e2b9200eee93be8b3bef6293d4419314b8134040adefef29908754f9c1edfb99ff7c77afc78ebf770116fc90b2bc8305ca8432f2c2026c5b0517d9ceafde38d86e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h912e8c755cd86116bc18f5dfc6bf8d7eb8392ff3412467a764d19d243fc6cc6c806256bf1d3e6518f7bfe5cab85adc505f2b3b3e8661e9604f14e765328fa6907de4f0eec509ee0bb43ad0e74970e6fb0da5a9b22cadbe9ddd4b5fb87f1dc31236fe0cbd94cfdbffc30f9932169add50a8f4d6bba42c3e67;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a699a45ad2cd871a1b8203a5614c3e9506d57d2d5f0fc79919c224291bd9c13f875317b9f17afb045bcaf4b23ef3325f7c3518ca4843f608e2799ccf604137ec7d65ed6812c35ca430565368756877debc64cee00340160e946b7ba5d75b4b5f0616f32baa1287604355756ebbdc15c73b5ee3347c4d764f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1c887be7ce68779bad60657463506fb52873a4fa797e96f4dc3e4806a9b17425f31462d0f67f342e22afcdf316d30488502cb6b71bdffcfbf3a46f11fe0bd672ddef7d78caaa91696da835abebbdff6f3b67c69288046ae9eff9638632d33b7296509dc16ff1fe9a4fbf0af03e33ec54a7b8a6fac75ebf678;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4d73635a207387e7398f195d68e3f5b07dc83920fd87bf56bfde46ad73a0e27bd3f4f5687854f1fc5280be09da41149c50ef8cc13498fa78ee37b72ccd36e8e36e561db1645f17a9469746b029e776731e49f81b1fd05dd569eeafa3c744736498eb87644a583d369174b40e1ff509ea13830c280c2e2c0e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h80a2ea9d0481a5fc5a7e4b04528771565dcad4495648f5fec72263f469ec1cd257ad750808ad72ec2a1467c6629fb3855a2e6368510119dd5718ffb5fa0560c0b9dd7fc10f9142be8fd0b70e49fb834c3fc1132150658fd724fa851e36cebc02708419d8cb63bee99f3bb2021b955bbcb9c162c794baf468;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h61fe6ed87e4010c7636945683223a719f280a1a2848895f9f9d616791e52a9597f167007b966f0f64b64b46ec2b531881ff38efcd689ea687c558ba8f1d0f89df7d1b0753669bed2e2d96acf398ad5ccb2c338916cecb307afe8817f5c766ecc10d0f63cf7782cf65102d85a4d7b9d3122e11f90dd76f47a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e82048ac050901d24d8040737074cf02a0e07d1792ec650b89681568efcc34f3e4e940a70f197a254f601dbc82b276b7e246e8444654a83042336b905f99f00c778a5ce046f06c411811245bfcb0c8bf2e7d25924c934e34c5e1b08680547ceade91b6e0f8d502c1c9b2d6f57da3940095a8dff2eb3d8575;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h180862b7b7268e80e73f8e0835c7c873efa1f4548c38639078f99cc3534a8b4d656978cf9d4fa1b5b2d1578e35c3c43defeec2558db3c245dbb767a63bcb64f7d3f21b24dddd26d5513890a0a6da1dbe2c9635aa0d44f0b24762ab12ced9e5b579672461fd2124a610a558151e9a2de5d95a331a4643da201;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha72e43b85691149177028b3ef79a78cf28f32b500fed3ddd0fcfad98b0acbd3707a28e7b49f2fe055dd89434254d830807d80590b6e593b6d10590ab884fd87dc839bc2a3ba846aaed644d9f0c8165afec77ecbab9d237e0dd4b49197e8e8f08d9aff42099087b5af1e53a7183c89ce79c8d0469466f1e2a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hce965a60d78dbc47f0343d426b9a0a19dcf34c485ad069b92979d2b61cbe4fe756dac4e5080abfa899c4aacf1e77389e549e477147de5dff6fc0a4acf672c62bacc8a3355caa148ba110eb90acde2f8c52013e06663bf7ee72ddb176c08d5c94281cea78b24c43e135a0079fada30b6ccc299f784c6cb8f6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha194d24d2def135ef6e470f718bd40ec766b966702cd21ae6098ed32c9054b0a3119c2d6b3f128cff7d5fe17fe103a87f9c0c5f0c2f0d723c171c4ba52313279267dc3a7a6262e8bd34fe669c04986744d179cb79c9878fa903db01bb4512bd74c96f6bc55eb61fec966eb62b2fb927ddbd492c6400f07b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19f07c9ca7e61270b1d95372b6f789a6570d866621e84dad25c75b6607eaf4b897ca88e1948dcb0bf326eb98b5d89246dc6be99130ea2fcc0b57bef65b3f24d7b6085a46c07d3760e75ee17ca2ed3fcffd3c1c15163d97963b812b38642d73b45a15aa7aa8cfbf62057b9dfe362eaeeb3228100e7428fdd05;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h122cbefb43ea81fc9b7fc0b5709d32bfd1a405b65b9121a8e64960059e1795707d39e9e710b32f00eaedc9beb495c6db7e826aba688bd507d0382c483baf4124ab69c01b87de7b3cf91c3547a9904f8244c80b234218e19cec1fead6535a8b79511ea20af2827c18f2a5bf49ed28933ad4fabe8b0e2ca59a4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12dc5fb8396161e93fc2e7d1970b90528580d3c5018198b7c7767604c095b780ead67ce13598caa9019790127df16e8a4f32043f945094738948c2d8d995c6f4cdc31cdb893114379ceeecef26a3921364e4e09e43106f37a77e207e2de9cfca8711008969c5d8cf137f2616c192a95903b580985b8e307dd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h390bddf5674d1bdabea2183e575cf41185b766801f2b70fc926ead9bf433843065d31ae2156de63a89fccb5adbc91b2347b39b7f21324207167622c172988c08bce9982b6e82500a751979090166d4e4925aab5ac427ef668975ad411816c73cc801c83454e7076a8bdfe8fb08302d88b1e5df4f2f239e46;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1fb6b12033711059a694a5dad72fcdf3e8f300977bc9fa163e3525b4fc76e70b8307d96fd0aa6d6feed2fa27e64720f39f33537b95ddad4eeb00a3db6195f042ee3e0b093a0350ce6a622e49507d0585424dc3c3af2a9fbcf8f5631315e89857ea7baf3c137f727d89ee7368c81882d06d3ce28133368ab80;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1719d14782a60240a55acc6404aff2eb7b5bcb8b47175c5a3848672cb400f8f2f79881893b8cf274a0eeeabefd656829e70014e5b9d8f128dc586e49e426a24d2e34033c7d9a2c98d529c902752ad2973185282c4a84da01af477fd470cc3be9b654a9da65aeb0b917d0ef7c6e37eb084a3df82b57fb9c479;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hdc3a4ec637a540c437a47c19f6b7570cef15d4c2f26c467bf30ba61e0fbf482ac3f225805439164f6dc88e29e29d0cd973fee11d9531b08a3c2306bb5a809ecd169e0fc5f77fe7dc7c919d6c465aa9950cff77ee5e40c90b00f2bd97c75d7c8955872501ada0c7d2688f16bfaa73445324530555944cae53;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8d6c6bf7a03729b9fec0f1ee1ca4909e6d04018ff3e604d71d2ef6d41f8ca2f27a5f840349129f8c0a4bc47f5f11bae56b2304b637019c3ee8dd5fb66178c9d169cf57d97053dd9b293255b1a46c1953b9b899d0e2d755186cf8e32e4d03a18c32b43443fc5ede4da5379049f6e3e99c394f22ecbef6698a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19029dd6f42193fcd6c056d0681d7958d5e4127da212c46d5a2915bf4a54108a10308f3f7f2cc70a260a9d5a7f9f7fec74699276a408dc834b64e27a566098cd317e00141cb086293dfa94c9851aecce27e98e4660b23df29b945183e4f7788cfdfd0876cd8c9b776dfb540d6e10def6732a07ef0014583dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h181408ba018578aacc720052e2400f9219bbba053a739f68524b3b22ee304b89b5e21c7e6c846e51c52ad6296b19a527a54e89ccdcfbbe163cb65393fab5907d203c5d82494e6a1e385cb128ea98ba4463e9833b12c1b8615269cc401753447af4eebfe47e8f40e82c9fec2d3a0ceb74f3d60209f265da2b4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10ace166a4284f83177bd395a9a8a534b5ec9bf15c6b655ec79966b98930cbf53a2ab7ed6e9669b8e77ec14c6d27224a0e6d2ab913c0e7b776fdd6c122498817a6b34e6930a62b26581ee72e06a96b769c8d2bbd3c9c99569bb285538873f2bd7a479e5ed711fb36ab26a9be7b9004cd8e8e33f74c4acdba4;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1dcf35dfea0120e3edfead9c4ef7769b0e1899373847e919b96029398e6d76a79d8ecd414af1b5b057b596ef96758250ec018f20a93608305a0b55929e90a1f66da708c7453c35d7b41aa997c455feb079eec9ede2ee13bd72c1b7b8b59aa465b555afa3b1f560530603ef5c1286ad5a3328fafeb55646e9;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3e4d5b9a7d501c973b40c71d5776d3ce20c522175b6e46ff3228bed09b288c923d9fce1a111d4fb3020cd997bbaee9c8bf29e333925da56b9a6daacea94b9bc6444ba36348b8e705738ffa6f57cf12c7d26ee0a1fe76216468ec0c3c460072ed7d6160b02a5aa36001c15be0624a3b21c403c67b15049504;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4a4a65cc19f882d423a87706f42eeb06254c4662bb45e79e2c5b5a3382a46ce8cd09c216630b8226f6c31442ab3a343ab61654bd9574c0771b40a6783fa66df8a5476baa39ef72a88290d99411c02dddd02b40c8a766b1616c17f15dcfa90e38148547300d6ba39399347062daf433761f3aa4d37be989f1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hf67505534a522b6ff8093e411bf2317816cd11f42ca961bea2368e8294bcf537244a7cbf69bda6c4e9b97e6a4cf5feae0dcd4275e890a9bfcf32796b1a4e116138eca9ec8c305383951c2d7e83bff33be5c775b75e1fb4823efff90c25da51c3b6b5ebfcc99a7fd2cc827dd14be9ca08db541294bb9f5fcd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hedfb9b4ff74f5f59bbb65bac6dc9e0e6ca1811182dce0f4c8bc406adfa96f022bb8c7ae05ec7937fb971b29c02caff6553ca7fe11f7b0a86ac7a04abfa3dac9f551dccaf14ba7e1320b494ff8da04ddc6614711a363a19eae30b48f8e4f2b08f4cdea23b3e295595cfdfce0d23e5911d42eb3ff6059d8716;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha4b307e6641172b19161dbcd1980062797b01ebe75b8bab2f16c9576442e1b19ae0cfceea1499aadcaf335d5826f05a1621d669f281103c79fd41703efc7441be181d5811fc175f604ad808b2badee0795ec06254ee0e70bd10d895fb7c837d0af1f9e6fc35d68c5db866de8e555272d2f3c69be4c5e0088;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1a853a84173ec61fb895e93c6d0d4ecf41dec6a86a751d641562b58ccb9365a6ee6976c0aabf40d44f1ce0c2ed0eaa095a2000f46478f89877249a4dd55bf8ac32af29bd5324d2ebf753721c094edcfbd2052364ece36bbe48d1fbec365e072eb53f0ae7378e3ea77834844bb11717f2022b1033bd94e11ae;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h39bd4fc460d39083e79d90e6326e11df0cb3826fdf4dd7355fd471a7f47f7fa1739b62696062e28d5e750d75f60eb86b4b6c85f572bbe98495477fc83e0b7e6f597ce9f835a873c0604cd083535295ca1a7e3f7e92393e915dccb8d83afa211161ccbe04eb37bf645d9105fe710877abf9fc76874ddf35c2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1541273ce264f20ad898ae5756c91d5f45d5ae1ff1f4204a9c32e9a3e4d45eb8043eb5ccbbef040425dd58fbd13a3b2766647ffdc0e390b1ff2ad9e13b70d234cf6b586ae429cdaf64e72e59b2849e66707c461d6429d438c2854ea847aac7a9b5dff43cf09b492daf573c359fc1915880e816587936cebcd;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h13ec8cc529dfde6130ce0cf8acacf07ebf6596c7352fcccee35ec99ae4bdd3a64505c88f5eeb67f79e53b97b76ec168c9067cf8e84972aeed606e1d7af61dfc287245042c5039a0196426a64303810ca7602482481dc4bfd7343062ae857d533061e976eb6438b6c748f399033322ac05902f4514a91243a2;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e88097f8bef44654bfa4e10aaf2d630826bdaf68df1de87adef4b3aadda7f01148a7e327da43579e12b79f3df2582f6e4e3b36e24db6d195ab8f3b324ace74660259a0ef1000c26e8a1d3df139902886302ce30e48f9d4f91f9c0a4b07bdaa5d3c353289a1c8682ce090e6309e00a632cd36f1da63c718b6;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11d20395339cdb21f6de91199b3cc546032c0bbe6686e60b82cfad8928b23ff6768566e06eedf76e36bf1c587bfe390bd349ddec367722ce4b052ca9d8a868af7516e9f5dddd0c4a5441db8486191f3837f92e01ef625968d26f5609a4d050f1240a165f387ba451d9b259e9df9b631217deeb9f2a33fbfe5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h20f125a7a5114c0d49df3fc533f38726e1d6a4bc86b6b75fb14ae49c0099d6bcc2c529d41d04d093cbcf9ffeb701e40dd1c81aa321f4919090b17a93e50f638bc3184d4b6542ced36f6dbb7084f45f6838ae7bda3c4bb74290f77315ae6338dea7e7d533a9538629a64e06b2a9b05364db0c565e2907d69c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h4a826b0899a84da6773424d8958a376c26c88696f647afbe6cd3fe26aad30584f648b83d4dedbb586c1d56c9eb87ce6b4097d71965864b89ec058842ea383e0bb22ac4cba5b4c8ec1279c3007f06ec5e024e6fcc7e937d38c25d471c69451ac619639e75ee68998e5cf3f6686a76fec52ed4e4db882cae56;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1be25156e799defb55b9b04cc1adc453a0d7a325613c513479105c769ff223cf2de73df00bdd6761f58794d518d3836eefa0092d932934d5a07c15c4eb92f5fee3a3cc97e93642cc2687c67b6a4ef4ab996a55c4f663057d0840d8ab33b718b376c7aec40f285bceb9794bd0981d388188eae35b7cdc2289c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1321a422b8406034eebb86b895df7435c7305b626e6379e4079aceba8fb9e497e2148962db470dd08c75b7d12e48cf289bea7fb238d850c34d4ddd110a91f09a7d7e967e5a66c45634ff0bdfc427a37afe1e4aa28d6694c2b748bb47e09968e87b5cd879e3aab5dbac80b659193120a275dc482e328ce580c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h12fbaf0425a15fb2481fd69ffaf3d14c2271a1c26ea7ad79a552544fd3cc7f116e1b7d2c7092fbeb727ba5dca9eb2930e91eac845e160a4b1aee8a65155f7ed73616260ace618a06e5d9d07ba33f602d70d67e99729a356e3dc1b3a47397e8c335ea8b3b5caa6c690642e741945bef103943ea3a948b8c40;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h8374afe783f4f1da70086dff63ebe6a62d011d5bdc289b71b8177e49e177a2c48139aff97cfa49ec46f534386065dbecb175c281fb0ec99616a7db1762fba987b7a9951c0bc121c4084f34eba09a5df0aceb8c57216244306d5c5ca8872ff7ecfb73a978cc75fa95d503313d36a224a751363062ea31ce34;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11b07a4661669222bb4d136d6b172bbf1f76e218c09bcda57b47fc4b350edb3d071bd309e7ef1836c1fe9374e3f3d5cf766960c660d92765ca91c8684f7cc9cdc8ed17286aa739dfa016544a961f9ee4dd715862c9bd0db51fe8fcf0101a92c1bd1e7217efd4895b3d555dfeb1a3d53d56ae0bb8d8da06408;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hcdcb9d0d10a8a0cf345fc4c9adba4d407ef600412bbdad46037fe621806f66eda6083a8f5768d9c752ed507b4160359e8de635d1b3c61f4110f31d7b62a56ee3552175814bb99754b17572874e12ac5efc63e6855a2c2130d68f4d6d77b117df486bf8441180e79011836e58b9666a28ff6d25c139eb58dc;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1694ad1f3a492507ebc45420eb0da887a7ae7adaf4c303f4b9d40b519c44afeb8a8056139fe2fe39b982d9d53a7598d7da5f496d66924cf4de7b2777e32a4718821fe6a71cc2d575d65bb9f0e558014eb5ce0212ae0a44e767356e16f322ac3b574439e7682d117c4b046ddf7b23c5a35add764b35973cf83;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h11b3dc46d39a10bf50b8d247bfa9e9276e8416d294b247c0cd07d218c919d1f9be1efa4245bf2b70e8cf5b8b53cad2823843620a261ae93ec2d680b3422f07cad907339ed9f4464b5b355d848f415003e7c1c20f7bfa59d72d50a6a31e737f985ca75725143de8dd73845f2ea45fd0c5aed39ebfdeb3e171e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2a8b01dd08b0de3c777c44f5786c563323e83693f0b2d51fc2c87c77e40e7b3a9f77750b25c08626696238bfacb1ffd3456c1a76e732e548f88c582cd4ef26022d8b8fda3d77c8c49d2f5dc098156416cf6ea27c740ec82ad642906af7678077c463926400c70e3a6aa675a21a8d5328eda431901df56d37;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'ha72a2a6174c50b3983d149143b69ad863993cc7334c094126fcf99ec19c322824599fb7490fbd49816db4d91cc82deffb977820b757f2e513784f322cfa7ea1620505d2ed4a90eb9573d28a3d5e907d47806fb65a48094fc20cbcb20cc5338f41a258b5682b6e1587e95dbf9a16a6edb6b022a23c3d3c07a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1285f37549a8ef898c44d5188987f1b4b8ab14b473705bca768e370224300ce3987cc4ad721dd126c17d3d62df6e82b7bb9f84c84b00aeb53b2caaf49e688a428d7b5c5a06377443beaa24af5bf0dfa1dc482c0605f2048099ef318ddd451068697541c8625735d501bda20af12a841992699a50e71fa29ff;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h9325d5c600c2a83b6371e82fc57cbb7b0aa656f32d8c792ea6183d7a755991c2bb46c792312cd1fdb658fc3d113c25e2e5a1b03441b325e72c1814dc9a84b3c5bc14947cd257b597ecfdc64241fbff0074732efb657a4ad5f9f5545972db965132f6df3859052a7abcbcd00c6ab76afee0b2d4ce10ff5611;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f75e04df720fa1d2a6661494f0a2c30d34c93c2cc4e8ebad0964c8144ebc35d236b78698368413a6783dcaf7c7a39c642cf6ca3e1a9b45568ac47ee2bc034f706bef94c59ff22c2e3fd5b0abf906b37978766fad522676c07b6157b572ae3a7c89469e87b1401de53f17acb3b45ccebd35811a6c071d4bea;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb0069834ae7ad0b7eadb291ce3ad6a1ec9fbe548be71788ca41a075940a912324863a097f0bebf523963472dfdd2ee72c5d30949ef7d2c106752717e509ea3b71a326ded2913076b2c9ad260e7329c825cb2052c3e03dce1375b60e342f1df426600324a52f02afb172745cdae9a703624ee8c02498dbbd3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h10267a9b384e3d01ca3316ccc0eb54dde845496ba84cd1421ed4e8234ed7d20a2496cc0402476d53239adaea4a2eebaddfee9367e250bc6cc1ad9aa2098d25c4fe6598b734d59c331db39272f50f81ea6cac68713e2258e4ff10cbb2a6b78732c3e09aa7888dab4781f72780d80873a963334d3fb4a27d6f;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bad1dde91d21dabd14c5973885d852ec2866f9f1b8732fd8a06f6e6ef04bf56f050c96fa64b93225a445d3eaf78bbe19cd7f8fe7e3c8da464d28bb5c26f5258433c9b9a784f77d38c2018ed970a8f9ebb86962981f4fb24e7d1741b9fea9de0178d4db8a58d168e068e9ee51cf802491d8785df9f91f3416;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h2f439c98de6dcd0476e7ff16626311014d2c61fd31e18ea6e9c9755920f6b8140d44529ac2fd796c7146f730515c3f7e389a034accc4dd1f224b1f2706b7133fa1988a802c6991a1d39837819a509d9ac8e7c06b6c7cc95409a1f209ef140b5ec7e830f27d8413a53c28ae2d7359d7d9c6a1b1039b481395;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h93955667ec3589b314e09d816202f3c0650ccb92f175a0e10ba365b85d45fec9948c3cc7fbb3d5d72bb704cd0bf270c5331d832a7a18eb42286bc863277fe0da78a667cece870ede24cbbdafcb22322ddbeb6d2063a23be8ca61f25c60eb19a4131036272877afc27aa3410637b1bbd545d906a07978e47e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h18585f1ee31a8c850759e415138eb148f1eb0246914a631c9f29e43af42ba4285cabfb5635b05c1f76bb08254cb2cdd841b7b71bd8e3bcfd0a2e14927dfcf79bf08383ef950ac1ddaf9b32203fb522257d3838d472ed3642d36fcab26af66843e713aa40a5f1a59bf477fccf52f9e66237f6e10b61efc94a5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h167c48654e8285f5669577d6f153be89b8e959a94aa3973338fb6b33a7399cf28c293986a9c78027cfd4b2eebe7e5f9c5eace7f0ef691d2a6db301194d136101a216948023a4398a5f5baaab6660661214a8843b23bb6e808a46331d9c7201ce0415f7385b54c9f36d3a39645558e9788f7d0cf2ab99df373;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h19a939064b3dce0a906086badd30ac58557679e6978a0a07cc4e7cf40372788b62aa39dbf3bc9b2e54973ea4e4ce685edaa39524dc7c54424e595559b90366d0f397a581e7cbb302e4839c3c08451ea387723d224c3c252cbce64e8fc9fb9575a6fa25ae91aae11da83d5b6d07eb722267574f9b01d042d9c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h14862d56da825f31dbd2d3a7e329bd5aa7c57d0b594e1ab418c1793c8a4ae6e6aca95c67df76a3f4bbcf5922db0ec39fe934a316f54da1eb81158779b047e651799f9d7d949b00d3930995b1051bd0f552742a9bbf9d6e3e97775b05389241637ac28d9628f9f446b65cb7fe43a1dbf70b7b44866c844de5a;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h3a307f5ef4c68323a96c4afc291e8f0d54438c339d482a6cee50a13989a6fced19b201eb327ec19bdf51fa085dcaeb3a7b20931385c9cedef1963e365257eeea1f989a4d8875bbfa87560bf195efa3d7f38a13add67d63a6ec6fe5590856b126d344678327bef75b978a339cfe6e1d3f8bef6d937f7e482e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1eb66c7c16d44e3c853e1f7ddce1a175481a131e158e1e5aefde346691424a44740655e3b2a12acbbe4483365487dec9ce3c0761be5e35512e36e9f0abcc619be270ec56b7483ff553e8913c59d88b72a335869b16c23d12665cee0dae28d3f081b092d2957a5b7db22b93b1c1efeaf4ffd3fd963460d5bef;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h15046df80b272a31fa857c8091e9a67967b268d4f6a5d543d52451db10a9d4670fbfdc277b61be71e93b16bb896cbf8eed900a83d716f308ce0ea59c28dbe24a7898659a4b04c5fa8fe502421bfe38c526dc3aa441c10e1b0806bbed27351e173bde818bcec8d0af00a3dfcfb56792f11f56ffe5cb3703e47;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e0287870dc051902ecc2faf8229dc8deb8db7b443a470101ea61b02128c23f6cd5fc0e69c1d1c4fceef1d6e922d5ee19fb07865526b2d62df55cd329dc302ba0804c2ed0e15fccdb1dd49057d6f808066e99b61fcf8bba1482b9f0697cc9ca5d0b099f41ba98fb2cd11cddaeda887a39ea383589677aa2b3;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1bd9aa50b3304b2e042bca97d9fa9e14d6f6c689619975745b9f144cfd345b6f8a874301d76fd4e86de256408fcb1d54445b25ee30961d301b7e68be3e7af2c2edcf20a0f7463f5b250e8019aebe8f2d3e9a6a76a1d73ad3fcc458ae927102499888957a673c270ab5c387efe56889983ebfbcd217c6eca89;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h536abc26a85e9cf1e1722afb2814a58bbbcdfcda4ae133b04d2c9c619acab0712f56d7b6b589de8f68e3c5c4705f6119ae24413a612a53d1e2758604bb6b86238323418572d9ab67af41ff552070f123b7a47bed3a2536f8e0dba0dde1b1035f7c156262ab0477a7c88fbf76632004ae90bf6ce68fc5034e;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hbceb64addea7a92582b6ae8dbdcbf3712d6eb29006ae401d5b2f7fb079c9ce082d9f2bb8248f04e9a23dc76f47076f10220885aa2777c632ca105a10d8dcbf13e3bcc04b414585c74965df934cc3212efe32f8d1f43b007d109aa64deba4e79c53ebf4999961ed5910153cdb732639aca32f678e26d537d5;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1e45438e1e3be328fcb0dbb2102621f13d7c8e3fc9917f6225b5e8137aab578e820de0476ef5c8b7971175fc751dd298bba6500e5489bd1b7339de6b52bdcb71d2152a31619a9044e7a3cf07c6acc69ef557e019738a27f09f2144a67ef9fe544c5178f63c93a2bc5b959567c4cea77e80d93e2771df950fe;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hb562dfb759c08db63c536f85add6323a030cee970c14f57316ab87d67bdf8476d706f41fc8c27ae523efb6e348a587cd7053791c6ac9d420a71e5dfe561808011435c619a5d1f7add42dbd41a860d628d952064419eed388c659bd243c112c9e18bbcd1b2ee7e0b4197ddca87fc4b7c78ae204aea938ad0d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1f577a43738cc1a4a5aad74522dee66aa20d7eddf6a048ce7f0534f3c93e47d59a6e3a2d28533bdcf00c8f5ea53514d246407773ca9a4c28ec1899eccc84285bdd7b247e52c65f0726e43e1667e13d50c92a0e6079569bcc46043ea6b86f1b7f553159af1721b61d0f1e4444105230ca13862a40f9e5ece14;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'hd4ea0d9c09490a6e7daf747e726114520dbb4e4fd239cc165de707f708c2f4fd3b4a5c6a45b5e6af946b6d8690f744ec87fb06935fa3dd2a4aa480fa4de323acf02c7d12004cc978efaedc19eea8fb039ff048e9ead5a07a69c2723feb28069ceffa86f227ee6c6047c3c3d2fdcc86c6b464bf439c6690c1;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h96b8a30dedeb56905d2fa7f32b6925ceb841c548e2dab5d43d1eacdfad0bf4817b51c17199daf7527062a050fa402772062195f7682f1d3f1ee4797bda02170650c4cf6b663ae7e890c51537ae8c728f590e730930f7e926d441930c513e4ed3f5382f2136696ca641fae1a68a032d8dad5ee0324253475c;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h77e4bddbcaecf1b9ce5f3d3937464368a20e7b0fa0ace484fc8a887fa47e2019fdfebf2858f8cc21e02ecedc8736bf7c26eaf05d1a476015a2af44dacc87b32784e588e06c21e2908f8596f3387ae09f04f0960f5a12958b89b19e6c9565e398588d7869f63e5167f14e4dc748e52bc0ec7c42f3fcca75da;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1433faf953618a9b1a4e5e6b2312b7dec4c0021891fd46b46deb6cc6825e068128d6cece2bd6294208998a295299f3d0d0b6c509aff3eb0caeed615ed1047982c87857bf6779ca28228d98ed7570e088d7c222538b20ead95da7aff7e0d1241adde90e74486f93e42aa86d5b8f70f9e3a7f9a8a0bb3ddd7df;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h54d67862c58d9cf3145c0613952683ce13f17a9c7f6ef091541a174e9aace15f9689de9df60aa681f86ec1a3c467c02aaa4eefa739e4fd11bcd814cd3258af2a7ebc29140b069a270c9a1f8cdd752d6481dbe2553875f1d13651842b5a4e20d727647758e39e67c66c12c46789cedd729b6e63c495a4770d;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h91067d3ae64d438fad111f468bd10d5314ef472a35bf7adecc8de66d6aa7a59c5106d8a19c6f6e1d43f086d1b9da05af6a37e0e11c16f2c46588da765f8031746efc5df8f1916836cb9031b4e5fc9d5be465f26ee8473043ba837cb1f00827828611abf75b798998f07fdc1fecdc1b4cd600ff56cbd3bef7;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h1021d6ae77e206004f63f8f5ebeb819321144c35d167f94a21cf798f6fbbe680aba2492152bb3a4ec11b6a2b1898e21b194043743e222dd71c4fce84308bd7f03a1cf4e77e526b4f1584ebb460c768d80de285d43e11696ec8f543773c76d778d193026a55eb13f46ed5ff9b16983982e9163bf07f48f6408;
        #1
        {src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 961'h129b43327e2e4551dfdcc3f07622ec8838e209b0de8f40d4d46339c9d158ec70a48a908787046e5715c922211a020afc02766397fa2a6fca15615bea076fed809420d298ee421973ff4ae342c6b555ee00bf18146f0a4b4253560217d0ceb310349e438840fbcff594a8cc224c947439a6fde75d6987f67b4;
        #1
        $finish();
    end
endmodule
