module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [12:0] src14;
    reg [11:0] src15;
    reg [10:0] src16;
    reg [9:0] src17;
    reg [8:0] src18;
    reg [7:0] src19;
    reg [6:0] src20;
    reg [5:0] src21;
    reg [4:0] src22;
    reg [3:0] src23;
    reg [2:0] src24;
    reg [1:0] src25;
    reg [0:0] src26;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [27:0] srcsum;
    wire [27:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3])<<23) + ((src24[0] + src24[1] + src24[2])<<24) + ((src25[0] + src25[1])<<25) + ((src26[0])<<26);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce93c434c40587a8aa8b1eff5252534140b99367f29851585;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4e6e389cdbf31b7095b3de7419c22c35dbc1ad807bec12;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4d6435609764948faccdf63ac26f8fbc637dd805423347db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13f70395081176e92c9f95f70dff399615f2feccaaf79c8c7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c551b242661b527debb3af013b534c190b525c59921bf64f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27f46312153918dc5ea7936314c5ed6b57f6ba8a230ebab10;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d60292b7d0ed203e411df4a22cd390270a20802991e77a73;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6fa9bc932a316ffd8d35c138dcf083162682db76420e1b19;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h80ed345da50b614ab1c5f8ddb1b9a14bf49c09db7440c989f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45852af7f67f5294e9b18f9935df6988df71d07f2d16ddeeb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79359055e3753b9756f060a0508d02c8937a76cb7de25c35b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he44581fc9e94d89230e96e66acbfa72e6ff461e61e471e9f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57847730da4a1650c680d44383ad6055681446d891a96a30a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd60945f0e31ae0a9e766c15f82fb1a57bde336cd05d2128a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7489ce181b4a8d23d1115a6cfae6e1c06c4a920ea8bf99ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h583ae8843551488aff44cbf24d9f7803d522e2ebce4aa33af;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hedb280eb342faf9795192a68e341fe1536d13a8a9a4e88420;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc72d710418d6e1d7f29aa0d35fd5434ba4bea46cec7c48037;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c383d1bf90bc1f980ab6a010b93720d64287e0c4c47f15f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3570dd1f263e0a8b8e267a65231e7672d70a00b1935b4f167;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e2ec3f62007fb2d2ae150f51f04cab4bcab6eaffe5b98dde;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfbe616ab5eae2a057cc7a7ce88fa5fb25789a67d06499d18b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc9991752d30236a9fed50540ec628ab4147fc2a4e2ae2224;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8da84bd0a4aef3b51e422a5bf5465b4587d4f4be2898c482a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4bc5c74b2f7a5290b7ae2b697c8a04c84a2dec8471d8f308;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7661646ec0ad7d3d6663c56404c2329e3c2e2e382cc3b787a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76600d54bc6ef190e7f3604d2235f9232c2f1e1bd58246fc5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab0aa129e460124143f46cade44ed5b4dcf32dfcaa1f83815;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc28846f8187631d99288a87ff67b633d7529e89efe8ca8d13;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88ce7dc2eb09763c554a225d3f92cff4db7d6dcd0f8771c01;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9616bc3374ae001c334bad70fee341e4b6192cfe94c628557;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac50e87bd60ab30dcce6eeef342e8a69664c000236e0d8b24;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he240b62b0c3fe91359c093af4ecafdd876b1797a898672004;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf899de73f73f53aaeeb83f71875cede7ae814f7a69e0e782;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9813adb0974ce394a36c0be34adaaee1b1bf6bcee61d4f78;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b9b6465d0c064afe460bb88c6181acaed1a2fa4ad5520327;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e5e42c8849df5729628df9bb298eeae85e1212000ce81693;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79f2e097803547239f0cf8bc1f349338a10365f6e99f572b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14f82e861dc1945e98511d41bb59d1de877bfb8e26ed9d48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2c7e6f7d2150c0297973a24b35138ed36c46410fb0ed7777;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29aa672ac5007335bfc66ab342441a27a372343f927bd98a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9729dc28576bede30880e7c6f1a9c0d2f2c63170b91bab8c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7307a582e5ac9e03fba0709a109b22457e2a208f5d8164e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa643be0f32efc2959a215d9fe70ce4c77c8c6cf31ab287f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h245301dc032edce39c082cac9cc9bd194499c8a7eaa83f0ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4fd8dfd85b98cdc42526aafcbb7a7cdcdcce1c0fc8b30c738;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf54ff5f4282f47b7356b186e2e658c0779aba52f96f1e6dda;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bafb4417211f88183e2a28c8aa5f9f66b82543074c17462e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he1b1eadca6a5706e4f83ddcf1d4aeed11c5fd95e7f65ec846;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67a3d59089d4dd10ad213d4fbb61a04585f7bceef421b42f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5140c47c2ac8aa1d2f75bbf93a4fc17154fc0d86fdf769064;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6371ce371d630f06070c9558836fc79e7ba1e2d4b9ea72877;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7e6914e9a85e3ecc7ff1d7c795a2cb802cfba823cc37b1b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcbc4ea663a480e85123d6c3dfede09cc588912da4a9a33231;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46534a6503dfc7e04ac8dbc0041519f251238230463535cf1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44b07a8d4c6116bc2a47d74009e549fb86439daec46e5d74e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88a732ed49e5fbe5e90d711bf160e9b642e62ebd906c00bd8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac7f1abc281913e5161c814e82e2069aad8add7b958ff3e8d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5456671ffd70b9a2b66d66c513e89a9e70cc76a0c1d9e5de3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd44e2fa279f54387fbb39a91cb047c2a65c3c6dac8250b67e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee63934565fc5ab83a459bd2c46ad335616863892dc3d9f07;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b20ffa24179c3dbb2b2cd5e40b32bf9c7e270344c7a2d271;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hccd47fcfac39113c57928bc33f3ade5f42118cddd4b9564ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc225017872bb53f2c9281834eb981795cc8b8284e53f960cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78d8148c31e0d4533f3a05de0456ece336c3004642d22137c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5201b1bac733d95506a707cb522b6a88800238b214567c8cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e628779e6c03e08112b897dd19a2ba9cc7a59ada0c03f720;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b9cce789e27dc8ffd840a12ef6000530f323efbb56bc32ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbfc4ac3230e073ead99a43875b5cacae623b973cda033c01e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h349b1e5f28177bec54f67081fb61988167cea161ea0240120;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a6942431e81100e15dfb2178d3da21770e979e06b01104d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haeddc9202582cb01845b8d7634ee36aa01d710528d90e616f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h15ccf564ef6e431c53b8d84b17b85d416cd73f31ddc3ab486;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63ed22505f065839aeadda5fd72f72ebf8e2ee5f6ff35ddfa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hca0a91dfcb0265dea7a0d955fe2fb0d0564f0b6b40fd84b65;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d40a5f02c0fc71193128d288bea57f0ed6be2e28870a4f23;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21a8c91c9a7361c77fa95469cf0d6a494c236d8eb1832e403;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed945e442ce6a99da07bd3c3a908f00ee1880910ed346fda0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f07a42694cc487257c4846c4dea53f73c2afbda31140ad38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc347207677240a79a37f839086c014b8841768d0d4f01a63;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a0144950f100c5c332cebfe8185a76f6c48c1ee4529e9d50;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda6ed293418298f19a888dd2bf3157d2bb0d952a656ee5d7a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb1660f84122754ff8396f9ab1048c6e35baf1bf9218ec4c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8116f0b19a4072bc98486e3b59e23c30b5c77ff04699bd999;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcee957d5b7da6f2d442d12e3b6378212a9168305cdeda685b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h868979ef49ae294104fc58545920637207dedd90391f34811;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h923ebed7ffb94500f1089358acc77821cd29ba99682747197;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc85c7d59e776101df5165d827c83446825374a4615463519;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86505ae890cfa013c84b5d1780720c7c756454d74c4046408;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h91a1b5e191f868709694bbd4ce6f31084483a9ed9a7c03677;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h64e25a243bd7c85c29346b278c587d444af1357d569afc2c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a2242b0296be73408d025a4c4407f75f7d74e07bde533b61;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h401c2459d462115ae1179351170d1fadc9867c556dbf133dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44d1c3eb6781cf5782d7c96c9a748703db95c18ace9ae753b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h555216060a5f330dd522a45fd25a127664efe84a6c32c32a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf546a6f9f2103f8d6338eb5b356c27e5112c74b53f2ca15f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94aa983261c518c82e13668cdcfd3cfd4adca722cf3ac7f77;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hefc0cfbb3e301c104ec35263fcfb9fdb0a46cef2dce48a5bc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h938dd0d0debda6a8d917b0daba1b2684b0af65e2b5db0df31;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7b32f527bf2980581a1574ee33bafff181f62cf73cae3b3f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h899c308ac3ac5fcf7fc403e7f8b3c145accc668a56c6b5b20;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52ad91553c72abf786871baa35c7c7048e92e9e50ff2e36fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1457aa5a0a862326593ac0b71416a5c592c84b020f37b8294;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87a7ac14273d51eed86ce3748b7a893f74f4c70caccfd9ab2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he1077ca7599a6633cb259a3661f914edf244adc574d933db0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8565eb61a7421f449fc1d109bc9dc80b3c0e0887f57f6e6e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ead3462d69f8b0f1478ce65f93bffb2732782995b4a16cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d32afacc4bc1b5c71a937ad5b2c296fee0daafa787088c44;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ec16a232bf7a2169ab5841712f77f4d0408fbe7cc49ace43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb967c9937e71ce39feb12f0df98a8569c447cbaa7cdf0a69c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h632d0e1392dd89a306cfbabf8438ec294e58431db06750d75;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3f4dd5498546c102af2022b5f0a770739f36d22dfb71fbc0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35571bcf0da3936456e2d815053be80e9d43c1c65fdfc3b17;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf23de514a19bf151382d303148d8ab51abaaed2b99909;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3dc5c296bf59e98290c988d707203f2450ff5e7631cc3e9e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcaf045256dd73e8d32cb7a051eaf3142ad1230fc3d83b6d11;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29829d9dd0efa62ecba68bf99b30ba0532d2622e9dee72472;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e6af331ac54a3ae283123e2f64024e0242e23284416df13b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc365f896550d5845046fd21883016d6be2d50cc3abc538a37;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd3d26f3f839f8f968dca341a1bca8281b5d304fce080e16e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59edabd2760c08ff06325a3ae104a5ca0255d73092d665058;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf61cf6a29ce75584c7c30b3cb4fef0366ee389daeacbb94d3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc7c3f11792c034bb804695735a8d1a68834002a66b17f7144;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5aae0c1722a18b0995f8005525207032015ff084b7b248672;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59bc72b06b5c2a1a905753b77b4d1c83f5e22e7e33f0961b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7744184a7a85487fe877892b8fa220f4201b7fa2b96ab9814;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2d05729fffeb34cd955f331083dc6048bf2bb5f117e82034;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e5fbc91c5bc0f02ba99c9e815a8074b808b7a9b6d48304a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ecbf1073dd1a32d442c7f13a1f568589e9a97dbb6eab034b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22dd62a6a32ba1591b171dc8c6388f160e78c1e46553907f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h907e05af04117048a912f1c2e1ad4695638054be45d906a37;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8866ed1cc86eaa527ad387bc328d07ee9ec49c46729f89bf2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96da03f58f8059a0b9d5db13a8745de2d19027430d367cb1c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a79bbf26bffb07daff29d9c63b96b91ce264581ab28e4d36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d1b15a0d11eb629cfe89aa369a61832114852d402b3fc408;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19867c410196364e8c7fc0e308b9c462f4f19a69bc81ebc76;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf834ec6e7692e54642d8e05a27f46043813354cd130f35138;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7928b5d72315922ec6c37dc8b0d2831b14a5bcc56af821912;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2a02cd05481534e479a40e1d421e2a9b5aa672b3742b26eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58633d5ea4c65c2292a7153b02a8300b481d095617bc8255;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdcb92bf58840f428cc4fbf3009c7425a1bd450de6a299ba00;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf098de525e6a953ba7be0f3a7b74fc7d77ca76162784222a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59dcf184353cf588f52db0ed976d76d902a4b824a445a7ddf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdfdb437718c3482df69301452888477ca51ae08b49bedf061;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d391072966afdf310ac35224db3ec20dcc423dd4886aa353;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1dc78603a21b21d65edf271792761281caab0f0c53cd98ccf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdfc2d86a2ce66f02b7394d6f0cba9ab7fb90316d8978f751;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb874142e5630e31c9456281ee740d15ecbf27a0141b4883e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h116960fdc2999d5a99eee557a65ee425b59036bf2836ae924;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8cf746b2762ccdefe53f76ce8b2880c011334b30d71527b84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc34acf904acaa4a2d9c690f63d24fe7632104676e632550a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he8c4cbb4d804aeffbfe3ec2c7d5dcca150246e5c711b0692;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8914849f0fc7b945e4cfcd95ce498151a27090fd6c4aa6682;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he95b27a0ebcd5eb8d77de506d679fcd90792adbd731d66a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e0db42147f56ed6433b32c4d8c7bfa5d16651b3efe3d1571;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had124edf230853c2d8562c9dc52fa0ec53008c48d20af6489;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h158008d07efde70dfc3311fa08bbcf7ece6a82ffb2e01caee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b0fe20b00b5443c209f7b4f381ada48279e8f9cf33d73418;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hccf467fc257c8715433333cdb4f395f8e15ceb2eebcb90b1b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf4e4bf8da5a2e3e599fa87645b222c3b03f9d6fae92346f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf47a2e77e1cc2b034b0d41d19984193312faaacf9d94c6186;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9cbfd88ed46bb498a94d3cb518d75fba174ecc0d26b03c34;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd84151700ecbfd49f75b5d022f01fd0c5b36ae970163af00;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b4fa3ac2218e6e3b558230adbad7154364316b89a2d17cee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h774451aa427635127a96ee057672f0870d7cfecc1a0b7fc02;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa2d6ca31d98f68c74cdc5eb76962c3aa836f820d67375e8b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7336bb2175b2a052de347d680eff9deaef33d2e06e722e081;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6e4bbc47f3757ed838244d9a3e2a2669a0c562e150354bd2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7f66721b9545c921d6b6756fb55ccf3751ce3ec75bf390fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h227077f69d141c01d8a0a1447dd1507e6512bc226ff8ece7c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b93e5b9840741482b5f7789867cc41ab2c2e9a4ea633774b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h293b1702a42b76e8454675c09e415a49a799bfe3703078392;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3f9fe7329b413e8862fdd0f2c1ca5fc8e365667be3cefe92;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha68ea8b349d0e73f694fb789fb805f9fb7ea882219951d53f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ce388d6b24dd1a63ea3d0de6dc9670857a19489b34ecc930;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2cb270fa627a051266593b90c9087e7ae2ebe5e3e760f645f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hafa6d08f1b85e994f49c14a41456259c20b596ba5a9f1e97d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5461c2cd164032c7cabe84cdc99cc675a49595dc1b0e8b372;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3a7b0d44874a626da9202faf97c7c02a7659839b048e0f1e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6cf1d2618e647d606067ca7c3b12ffc64ce9cb10fba39a5ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86ac85964ca69a5eb74dcaf16155e30e56c0f92729763f385;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b715d9f7a4d7c4d743e531dbcdc9d92413be2d06d0731d23;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d304d4317e409751bdda3cca47fc7ffb513602356967c08b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73d3845ddf5ee5bb4a050885a03c0a56a49c59d2b7973fd97;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb14c1e43b8c8807667978168b6a357a08355bb9b2a480ca77;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5e5c3b617efb78d76f10081c68c55be999c4b729805d72eb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a4e6dfd1d08a93e3647c829cba191d1ee7666273f0a9ae16;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4bf269b977ce319bd137bb9ba1bd768050a827b7419556cc6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h493cd333ba56f8deafe47918baa1b738e879751e67b6fc242;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h83185b1df13e1e7497efe822f47390ae29a22f8cc98254e23;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h201520d9633755c16673b1339975344adce0d0ab2470e3aa2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33e68430801308d970ad8c39929db1189ff14bd1a37958351;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hedf87b37cf21e2176eb03e98bd3ef1c217a70d65ff25bcc26;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb1798cf1c730f088f5b3b9f3933e0e0c4927200335af93401;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5625dfdc465029e6b44790dd6b6ea945f661f198d987f851;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9b66b308e7101426412d73176c00ee237bb4e0200ed4817a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdff21a8d78ebac2e8628f64c67d3569c72fd80e73fb046212;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a7b66d40fb5f214cb8f8b4d86ebd2c70bb56a73c38f3d2f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc87b31a75d2fefd502035a78b9ce7fc670cf8523051679263;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c1412fc67e326af8afba27b392f636b0b6b3397fd4a1f2a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87c0d961b2c15eb4edea8623659c4cf0c98c671abf62f6db4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h584e67f85634d1de1d14510043336afae34be0860776bea2e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2924d544ab8c40ecd3ab344f7b8f4e2c797a67c6c71279f0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38c43233c765a2ef66091f296d70d2611de275c0cc05a16e1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58ad07667ebcb8512c1eff5cd3cfcb87d2fb8c1f336c75726;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f6ba08976478e2e9dce8f197f4ff2da47275e8c6a0916225;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26ed639af450e65df17633146dd58bef27a310335ff253edc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he00470268a23f36b6475bf37ccfb44030e34bb609c8fd0915;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37584ddc7226d0fad666b728a11718e527e17bb5e1519d85a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72b9772d57b8f963615429acd187a68e2238c9d6be3537318;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h976abfd2e77c15d45709b1f6562816dca0965d9c9ed17b64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a56e61ae00b91356552ac323e87b1bd1d086ab57b2824f14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heac301d38fd483a18b9f68d4a532a8ff300198e2c1756f3f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce26711e0bf0ff877985a63db87b3859fac77f5d667c88ecc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9b9515a9cf24423cfbb511c901f7306cb60acb18153e5738;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17d67c394feec730687e1273715e229a6ac6522f0689453db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde5da484cb02759b902fedfcd510716ce5436a636c2afbcb0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h622182b20120b6f6e6cefa9c71ca3d4a1d3eb1b48fee1bfb9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h185b3ef15ff6cab8ec2d56ea1381014477cacfb296e5c5bc6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c9e95014b08f2be8f85a965e7225f8a0ea3dd912ab944991;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69e046038c727edb4e1046fe6b186380d22bb8510cf186165;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50cdae1fb329685a0eb59e7edfe89e7a94ea18a799823397e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22c335020a146be67e0cf7cb69eb9e6768bb4d49d22d8027d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6817144bcc4eb772789d75b32103a9ff8308cbc9ab2261c7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89114ccf1247dd506f7ea1e37b31c631b7945ab98e015c9b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd8136a33d755b285658459a21dd6b8cc6fac11ff5e05ff94;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h43cebbc479e0bc1ff747963afee6c4b5b64a8e677928e943e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f70553a1d0c1fc0dcc94d7238993416b7eaff634c103a27f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h817a707eeb060554265405139389b26a20d9fa6935df4fdfc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha63d6d22ad494b2c268fd6ee76bfc54a87ca356848d7e267d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h678fe26f7d394d26749f5acf3137267b37d7444f1a7f34340;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc18b8a0d1ede07f8de9edb4bb3d12677d1485c6b5cc312f09;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4793ff65d37a5886a89807a2724b28c958a89e483131aaab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2de13786494503282bc79e3156fe93265ed722a951928fb1f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha39710acc6b4a1fe233e6f2c10aad0b94dfd5c348349f291b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9cc988a0a47836e55ca8de99f31036150dba1e6bf1888f6e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc12a2ae2b827fe76a4d8b179ac2ff6a0ef491540f17ed93bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb21b4fd21e57807f5c43321fe1336723e6fbadac507ee77fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h218bd072e7e972a2c88b9309242bc281e4162baf99ee771d3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d01fa89f1fa6a684b538dc87cfcea97b2397d71278d8b919;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h831d1d4b5f218939f8b3f63df2363b655686dfa5850fa07e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd989ba63051216a7a5609f77d3b23af5161a26f1d1c94657;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27048fce2c528a0d095ea92feaa501ea44dedf10c2f818b2f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h277c94cb8e68824393013f8b98312c11e0571634837cf6da1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0d828ecc8cd80a6ac06da5f00368527b87e6450043f8388;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d8368571bb0019e3764443c7648149b0cca667d3e2b5fe60;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb68558b9cfb47800cd2696b0af2d9e73babc181900eaa43da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd92c4b0ab1629c002f127bc27b946147cf8a12cfc184a8ca;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc651c3247dd590a791c84fb289696b29ff8aed488503ba45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3644338aa26bf5f1b455b39f068dd3cd302950cba024fe578;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7dd7c5f5bab9a367d4c376c33e7f9f87f43c91d29dd91450b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h981f0eb1a0ef3c9b939bbfd7705c04a4fdde038d61bccb9ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h246400a44b6d18cf2f871093d08b44b00f7dd5182f822406b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h813385e4fc5d6907040f1a49180d1900b6b2ef43ac9d4acc2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0db196c98731ce236a3ccf3b5ee63e6c1f12013fc2ef87d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h267f793aa91f3102a0ff7ffbb62f910fae15680b1b94725d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h36664f515d8c571380d954580aa7d8d974999b0ac8468d6a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7e04e0583840d58496f6881c37f8ec09c3f4ce71490a2664;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3874fd94fa163d4ab15be09424b058bfeee8d1bef377d291;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab41ca249106aac6111c78c858a5836351396771528192637;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f741e49acff32dd05c6367f282128d848461d8467a5a57c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63d20d327c5ec00fc7accd80ec10e34e6c061fca6ae18f68b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b1bd8a339e3534160cd1026d4aa679ba3261e875d7e10e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfec23daa8388a3b0a4f4d39a8e9cf6854134b3410ce29bf67;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29eb4a72923c302c3b582f225c4474d920fc38349ea0eedd9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff6b74be2ba9ebbd4294f84ebf9f9d3bae08d08b546442760;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h909775ee5f1f0ea9ed9ad03e1a7d0967c9390864067a70597;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24f844052e1cb2d0d745d82561104ff16e0eaba79d7d64be9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11fd8300af3ef21ada25a116ec683b51e89798bcd1e3a5c6a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hedc7302937196719538911e5dad54a9965c6ff81add26dd99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h362327fb1c691c50c88fb4e4ee6d82e449313f1dde1ea76b9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd95ad3f52b7ac8e97c8e548b5e446a753a7ab31efafdc9a78;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2300e822e346b52fcf0a783189668b1b8591b8b18c1bb100c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3f54ee514ce364485768745436c4392ecc5981b3955f5b2c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h298ad08f52731eeb029789927df5981ac03dbe4767b7f2805;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce03530c48167d55891b45fcec28ba2225e39b7badd99ade2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2add2228a2656ebfcd950cc1ef4d4fe1ef06fb9bbc3a0c59d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6af1b61a1ea33c3df56856d0fb1a5f53db568bd912182b3c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52f3a7fc4956af3d7084a5173fb5040b1a4cb448cd6597e48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc076c66ca80b956e5931c6c2e987b940e3d04d32a257ab8d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h467be776426af989ce472ed14e3599f202867c4f226f11e38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a935e5c04da601d369335b7ff861de88411519396d12dbc4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he28172a1a418f2f349cb8f9f4cd76f9e760a66b5d6c1be72d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha241eb109866c0cb918edd1e849fc8b56149cdb6b1ddb1dd8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4586817f74fe5f9d2aefc1e5ae7b29003ae4e065ea5000f6b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77197b7ae6248da138022e0901988cbedc901086dbfadbdbf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc25b88c5a122bc58c255c9553f73edc4f102e7940f2b1a587;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha29ca784d6ce69c7d0fa21b04fe71cb8523493fcdd68efa17;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5400951b3e6ac0116112c21d400be86944c1cb43e53ba48ac;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h85cfbde80e8882ea1d14338b26aab759af72918873211aa3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd586188fec84b7d9c632df33fd6791710d7542f1da0462538;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h200c923cc72d978d30b5b01b816e4692e1e3a07b7d5b49f24;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ff884cdff701f6ae3a30fdece6efcddc3a5740a2239eceb9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he58cddd504759d3417eae9d12b55c6a7afb3e5cbc5a18cf92;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae54b805b80c807770b2917ddc28c754ea6d02eace1a358f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6dca10e38c171b0d85b19f71a00d706427a68159d510af32;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63c84548a800abdfaf33843d0d573baefb3131710d223c0c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h91cc4d2a33ca1d9900e49e4441cbe447a6a34a62b27b1cd65;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb272da8c6bea4ad09dce90ab2509b88c2f2f3fc3387c1f017;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7eec1817d8a08ac51497e0aaf7c02a07916fff3db58b0e0a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7dfe7866b5300a52ec3b34f510f3f5458933e62a26b4421c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20e89cd1bb75b5b3c5b6b10ebecadad926181860e63226504;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb1b7d09c62e9eb85178e16920c07973de67663890611b096;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ca637dea5c7f01be18241263a2fd532e701e48c0839d749d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b519a5ec63d31ac7da7ca428e8ebad3f8a053cd1e2a4857d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2ed1dd839509174c8b883fbb15b2fa371dfff6496a2b3daa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33b494a39a68b11d7769f73921084ec2f6ecca9432d844ad1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h399678a29a7082424b933003fcf4c9c79b6ceedc6fe534fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haae044e29a687d1fb22a00eff483f19e3f0336e9720ca6b6b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52eaddba020bbd663880556be1d00d427eecea71617d70fa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h754558da757cc1606cc3261ceae10db09d2f8284b1c131113;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda1b3befe85b2bd0060ca780e48bac09a14ee642292948e36;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5eafb131db6e77e5adb3cfef0868f5711767b97d3b01a0e23;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h558d6060d1f8636633021fa108e21e42316cedb95318a81fa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f1772ce1192342fa5abe9db4b23974fdbfa0e2b338d32b0f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0376fa3d27b229cd74040e33109efc5369f55ff31eb563d3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f52456a4b6bdf5ab99d0e431f0154e323b3a28c19dc0b4b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd39fd6a2de7d56341e69a3d58060544db506393818b2a6de0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hecc872a98c902a3de5840544dfbe513f6992fc5cf56b1d664;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba36d1f3e5c7a85ce26e43d7a129275e0efb8f1b53400e650;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h23b411b176b5f4d2a9178c3fc9cd86ec9894a90c586fc5a31;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha469ebfe2047ba06e2150188ec58cc933946217970771073a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd32dd34c146f74b4bb6943082b0fb1ceeb3fefcf482764a2b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b1a97652975cabade584dd8f4bd98ffd6c1deb0a6a601cbb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33625ad592aa2db9a6958a4d465373169f9231ed33609d78e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9806016dfda0ea4e756cf8f7beebcea3a6c2c86ac2a7f5287;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h43a4a24416a9c27e5470acebc43dcfa212b8b723373a4bd11;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb54bc33926e8678bd9a04fa84d9da99beae08e3fa85abcd3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h36265230a64cec3f898c962c3e0f475580415b212c34d4c0e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3dfe11004935101b13e2f2223132abdfb57eb2991ca44f89;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4ea272325b651a7baeb95f832e935475f664579b855886d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h252782c6b79b0395cbcc951e4c5fe6d4105f44533070f2771;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52083d7fc31b4ae91571c8e004687a02577faa0b840f5de80;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h759b958bd60428f5a1fa2b3d7f45fc366e492927c6d992abd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f5e52546db4ff12184bc4df5f2a198de4edd7c3381e73a0b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7691d168ddfdaaa8beb4335e361b664208f31e442c05a9aa4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee010d77cfc24022ff0aa7792f33292f29eb85e2ec55807d3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57bfe3543315786fff771529f659118e1d1b8dfe6669f4480;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc55ca099e2f1afb41f0c129bc25009cfc83abe5421b2ab72;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h204435a4e2e0f7e63524af4c3389c29e316399bdf83d28361;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e0f49ee22b41dea225d5aeeed0e030e8e0381ec69134f0a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13148fe7d40759eb47de6cf9b3896cf286c2253f5b78c474c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbfb8a55a3d0ef2594de8cb7ebe1b2c9eb41b140b1cf0022d6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f30ece07678e9ca68189fbbb1e3b4b9faa86d8c28e38e20f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34d6f83585b91475b00fcfaa3f169c4876bb06642dd85ed5c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8bf3c034083e2f8d7e899693de7a9d3a80f9488d15a90292;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27ad526d9dd89d3883ef219db377d0c5991c0d2e5f3dcd404;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfdb3f48d66e59b3861a180a727326491386d350b9efbf82c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7839e777e95ea1537804d8afa65357ee8b3c1cc1788c8619f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c08849180fbb86a3daa836020c84a9897606cd00e0980440;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1647a777e136ea51984f4137a4ed03eec398d814921b1eeda;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7bad00fd3e566939da9af5cc2847ecd846a79b3ba857c8de6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf26a17724ae593393b0449be368dea654b15c44ca7659307;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4986348c11a68f351433fc78d17863759ebaa859c3753ff8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6bf218791ae1b8833e64079a7047f1ffd3cb1336f1710d720;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88204db0c1ccfcdb132eb8e42b3fd600e4607e39202da5004;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h602895b2805f86c66af85e4dc3c06afcd2e51d894ee7e582d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb45cfbca92442d1cce17965d546ab0f16ed53716f029d0620;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3bc9fad13ee03d6f5c7e4aeca3ebd8cc79d9564839a9f430;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heeab119eef0a0a8ce9aa691c7e2c97a36018e912b2f4e5862;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41cf8da929050a340263edc312ea6ed3176e2fba27a43a702;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h512281767f5b061cb04a31a0b8d255a9ce1ce7665ad52281d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7fe5dfa6b39e4409ffe7898acb79832c3361d2831168bd19;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c37ebdd5a2aa9b82c5a8f4a380bbc732f7eb21a7c1785b1b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48a6b4b19b0ff18098b0086d299514add9119b39dfada5eb4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61e3a1fcd13969fd86e38aecbe1a7a8b23fc7bb05c2720f22;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec971bf368817febe5af952a016c85e625fa8c8830463c0cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9783e2287c2e8a61ca435b34a46f321709802a267f578f997;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf514be1348f01f8372d75c7f82090c60b1a71b3e6374d4ddd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb90f6121d23b33c11981f358f0e72290fdd4df98cf4a688a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3cdb365ee752909d56698f1f58ae331b51a8650283db47758;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb33f1ba38c0c0e9c0d9ea26ff97098985e581180bdfb0859f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6aa18f50edb2b4da2e1d30444e1270d813e35cbaecfd3f2a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf41b95714858666ca364321cf252e3992caf7221a14bfc3fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb20a25f384bb62a6ea3d81167c46f2f4bc42d1b6d5c4ed31f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95696b0cc3ca50a0112ed913723cd0d750a0739d805765fa9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he663682e7b2eb13aac3bd8a7e0043fcc6dae3f0da47786ecd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c33b2daeb63c86fb86f8bb2dd8a34b9b1deef9743d4aaa29;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ec6c7190d605114021157128da0141e73d33dad7f21a933b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8c0c2aa864cdc39990fabe5b1ad93c9a1b1d0c49f72bf57e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4a6624995041b6d31acc02d59a4476987c1cd8e7d71b62a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h842a5740b2644d08ce4f7e3f442ccd475649dc580520f80a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9632256b61aec29426c7910b75c9333a306b9a4b6a7bc3c86;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5daae81089c089f5cbcd45ecebd4980fe21d6fd2427031e1f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h284ac77c6ee8f79749cda0f27ea9740e32c49f2d4e075dc03;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf9125e9ceeac1743ce7d85124878b487d738fded9d42d0114;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65d902b94177f24773c76b129248b4c07191c15ce27b93be2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c47b85c2e1f6bba359ea2caf80aaab33636308b30c9d6c65;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2cda7ca20c9c021181314a110f40d49ddf9ddfe91004b4c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4315ffdeab4124be2c8c55c3b0c48d13171ab310ba6c58cb2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48cd5ede4a2b7293d268e2a8a7a001e535ce433e5109deb57;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a8b197ca86f9ab979f1c00a0f577c44fb2710df9fe98afc2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hadaad6c6b3a38c9b0bbe0292b441618123d3c89fe4ca3cf35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a338bb948587ce65065cb3b017f91f2ea3b0b17f776fa52c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f1acb9b2dbcfc64bff386b377dde941bf6b96708c61b45ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bbdbd90d343245b019429f25deb4f6e4bbe05b78dc50f599;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdce160df4f254a1175699d51eeecc51fa0de5f3b1b3315af3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3b020066b0fbaf04050c4d66b6ee2cc0fbd0d5e2e3bafc2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6d205662426ffd6e0c27f6ceedfb62034806e6fbd75d073;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b51235b2a6b829b70163be11179dd4286906de7fb0839532;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ef0469427389c28ca861a780b227cb5cf4bfe053af02ec1e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46751209b0e97128d471242a86f3a2fd236b44491cfc849b0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b46bdb90687daae8fe755206f4912d98bd6ff827d2ab2bf9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h507eab19f91947f1fa47673a38cacfa97110ea309ddd368e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf96b6c3cb034f0f85c58bbd679b84bfed8b98d0bb5ec2ed8a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b91b86d189cb0256b2bcba884d63c1fa601506396c359fb7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e6f031caa1cf084a3b9ba8ccf48b40490a0a338c5c3319d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h104305c10bb93d39890461f7ae7202bb20cb7ca8c7980b27c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9dd8dfd4e2a7f58e28599e81cecdee60de82d1c7df9302958;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69b9566b172d5324b398fc1c1daff41a5d4d5e0d959f313dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ff6e3f920260f74ad2e09a767028ecc42a549211973658e2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4356392f012f3c5fb54db2f797f67fcd27cfff9adba687d9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8739f376a7ae3fc3e37d54f87b96cf9bf9576bf8dab34ae76;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h863500cadac023640a4416312b1a15530a3611df161aa1c5a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0c415d932e955cf46e148834c3735b124c798ee002de169b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a0df4c4644dd82d4dc243e0e8364023c9668fc91470d2b57;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8b7a910d97ad247721140b88a02f57becbdf90a734340a53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h635ebf62bf468e9df4226b08458ed66602116722874ea3c2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b1f8321a8ee74dab3c34c3d3db516cb5160fda00a2dbfd62;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f97a22dd7629e7db8a59dfb51301e289579263d8f53f0b28;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h265acc36f4c9e4a85a5562d536b4bfabf9218bd14dd8f8053;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6da6a643a1b3ff98d6f7e98f9714fe8c1c25867bc3eeffc2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2bd3a22f96c423fc14e60e04288807457b94fd4ca0dc27c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc14dd7265e43b5e52cdb6dcf5287fe9aa44bf3896adbcd3e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d444d8d6f0ed3f0ed4ef32e192efe2558665c003874cc6d9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c17d31b354874266c57cf1712648b1f04a9702683ea92633;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8976c57d986c44f492cd671a2fcf3458599db0b233d19c07f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h341fb7a6d31648479acabb90133b1b5d89d7c9d31e850e75;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h905a20824d0e64777a9fe66949fe5a6f9e2eb45d0783e1828;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4c88a6b5385f9a28b4cd35734157f1190cc6c886a53ff097;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5f66c3a6ad28e9ddd853e572c78d4b4fd9076aad86e1caaa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c0a6e0f07a080044dae756e234fb605dd241c58eecfdabe8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hedf82fa7e8461dcc439b61bfa001685d7899039880a0dcbf8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0b682abb845591e602a6630d03b25be72fec0cfb3b5b0720;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9738451a9899ac0e03e9b671479b2e21bcec35a1089d6b245;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h898189d051dc9175d51a117c73351ee768a4d12140f95c16b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa497c27b0c1b179b52a953768ab8e079ea597f8aec399bee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5844c5f16357962c993299d9fdd53f2300f60925fbf4f37e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e1ee96dde014d08953a3223913f2abcb2e125439043b956f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha54d7a23b603aa5f927120eb299dd896995ff1eba78aa3612;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2be48bad0667e1d8e3e12947ccc30591e918de74df531465d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3571aca1bbf072799d513aa98127a86fe055e868b222d8257;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h172c6b848182bccc7a9d0e2e69d628820edd4ab1ef1793e8d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf60fc9a9eba888e94cf21ee133ac3d4d503e4fb8e6263ed48;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha75e34782573d6525421821c6d72f8744717cbb91ad58edbb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c0c7e1b026ae1e154d2c3d2dc0a2e9f25d0fbc11636fd581;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f5843613d190346c86edd9c4ad44cfff5c30b75c030a06a9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h645fc90c08bc30174bfcfe3499eca28b71b24b955fbc3d26e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcfe0ede92c097e618b1b72521583d142939bf38d0947f770;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26490b6a48ab80fc6475d1b6f93010f39d58592684cc0c4ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he403b677054831e6290015c9e6412dd456f32a50bd04b8ab1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f72ca6df1ec5dd973e27633d7354910c23ce88dbbf7cb2b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47e1b1ed494717f8b98c7516b6421bb7c5ef27ca3d06492f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2b2d862aed6475edf2f4f579b74178938a1c81db65af6ac0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h641e90e5c4c8d77288d6a0815d63c955d35dc55cbc10e86e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e8ae692041127519f98e388fcacc70ac9aa68c41fdeb08d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h726a49ec5e7826ce130daf0b365cdfe94e8fa32e1daa6ae32;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc2c75e97984507815e964a446ad12c8a0d636665ec888b397;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb79dac4124e29c2b40c38ec5d7eb52f55b23b8668284fc4d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9011a39fded86671225fda89daf356fca794f58b6166d4a2b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6794b08713df2884f1ae425a589765bdbd512ae9cdccdc9c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67064a1ec2fa2bf68a3b7da087b3867055e87843a5d6c6e91;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e91311e472eca573f647ec5db898a6e4a1dcae640286e808;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc387774218315f6648fc87723d566194a2156b188547eafc6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7cf747ae19216d6e51bf57f34a68fc03f8a7ffb7cd7f2d51c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1c2cfe0c830ae8a07ea44a2d378bce6264d0b460cca9d97d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3cd39db638608a4531b5abfaedd05298748a73b602960c823;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90205fd7c1e610987d861f9aa5352bf387bf4050240d4a08f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5921f263b58d5d1e29be03029977f7a52a69a6721739cff2a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb68873e698a3f259dfdfef5fabad31da76bb4472e5223b3ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc749840836b18fdfee8c92cf4d1d379c4b75ab8c97e31918;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33be5432a5bf117bbb631fcf5d02c8237c0f8aecb8e52e7c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb69577eb869e2ede193d12b4e4d40b6b9aa58807794452de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h577b8b6760349bebbe53f1e59d2aa5b7427c6d49461235236;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd41235df1331a5b33dd85e87f420d20365b360f4f0a9e43e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c512f91f2557a7a6379a38de7a4fd564aaea8035c11fb804;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f4073d1bc89a550166649678901fda0f4052bfc4ae988197;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5516aa5367838214699ae02bf5ad310ace1bff94b22624f71;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed902eb00fc025f7228343889a694971692464f2e8ad53a79;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h745619313ffd24fd2f3071e9f8f7f971411ac87dc75727d5c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c4bf1a8be21780c11feb83f3cad8bf47a4b405be818cde29;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce1ff4a96326ef4172ecb7ed289715674810df46e7f535a4e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h412e486261f8673339c398a113ae63e62c12e1c7e42b75627;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he50b90e05ca6840e23033c6c7fe8f8cc51cead8a0eb4b9bb2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8f085af842968ef0ee018340e31f2a1887370bb836a410ef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h251f37fa91d747175405b9b814973c32a83520fd2d41c154b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3efd20845783901e6eb9114478f940a0ee0ccd072aeead69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc3b9d21a84dd68ae411f4abf332c46832957611ad8f4e944;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfcb1018ae6a088b078460ecc2ba292ee2d085946115ae7283;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h299ea39b2d4251a1d25bcf3692be7b04dba0b6208312d6955;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h97c95b37ac47e888900fb14b2aca8782a3a8a673d15bb37a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h83ed3eb08dedf3b01aeca0d249df7add65c5b9bcb64fa29ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76623fc312f9ad6b706aa763f462ec1e4004bd209ea85f6f2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63f72d717fa72dcf9eeae9faafaff84cbf658955d3c3a3202;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0604eb7224c6224f6833afc1c6300b031fd7544406b078ce;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc2630cd1c01c4f7f0839baf72c5b9b409077d788a30009316;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20d1ad1773af06713f442409d9c0c477e8b2ea7d79877dfc6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21fe041de07918e4373b6bea05d6d6d52054155f2742b64ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9389fe7f84d1a03019784427f030cb79109cdee2a7b216c81;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71bab57d028574489157b11415952ab96bf97d9ae9ee877fe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc7d5e1c35913191e06c97b17096ced48644a9ff723fd89cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa77dfe8218b5601f209b4d8a2216797d0bad3caac3f4bd9a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h758ced86caef080b064be471b43b845e40c25ece28a82a425;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec60b8631a0f6078c854d318177cd62ee0a93ff47568e259f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9fa0d954407e272e327a29a08ac39221256affc2115f948b0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb208ef42f88c8eac55ea4a34175e83eebae88950730f3cdc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3fb2aac8fdb30793d0de00680e1df5bdd381a5c1481caa816;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e72c0f990fda46f037120087eca2f0ea74d3ecf22dbeb736;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a6c3481d0e86fc610a34c2acf220abdb3bac85699222d90a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd8547e78fb67282cb8a2f9b276b53d06218906136b450b7fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3aa6a4887cf2cab6696bca3745edea097d3dd6ff9bc2e9557;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e18e060f591e8a8924d887b71e3f1b7679a476ddcad976cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38714cd3c1fc61f94cec040023e1abf8f097fe76b9e5c9369;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e3d29fab3a494c9809207b1066999ec5c8d304e123243c9b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd68418c148de2c6ffdcb67c7f4083389cb18a8e92378863d8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75172cee75c3e534aa4960eab3e659b7b8c68ddf658b1fa94;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hacc5e47e91a7004c982643f2c5f4c1f62a910f139733d5f1a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21314e210f482e36deb68a108decd7ad77d5012180a43f806;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd54383d7c6b5ddd265984e8fd54beef7c3c5c59daf557860a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c1ae17c9b6fda54e5c9361fb667efb72a5cfbd58c290f87b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30306fdf8aa40107a7eea4b841979797abdf94a495bc7c246;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9feaa570ac371de0f2710f9b1163118a52628b481a4c66c32;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8a5a9832a88acf60fcb36b805464e792a57819515ba8080f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he35eaabe596ad9c14497039d567f3e0bc66fbed5799030eb0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd92c4487f0afd523a001b40a7eda7b967b3ec1eb2dff0fc7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a59a159f3e50dccdbc57164cb796cd127d9918cbe2b067b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h470a4925fb52ae935403875a3ca1cc4ec47a4d8b8aea3007f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4bbf519db301613b102e287ee889dddc3a337659c74661754;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd22c2ccc4775470eed53eb648c733d5290b24418b1309bdd1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d22147175c2210a6d82226ef1e170a118e8950e83b96f4aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7f8029edc2021e814bba0ef91efc0da29daa38cb91afe24d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96be9e47af9339fc40750a24af56fff58984946a77875aa14;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7407a736ed5d3520ea5656e3a807fe92388ced9c6aedb0e8a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fb30c512d69741022fb9524d540bf41cdbc70fad529e15e3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he8eb47b8b5ffa20326f9aacc92a722c0a614df636a7b23030;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e9287c743ced6d2e6cfa1a2cf27cf31577e7e1ffd7b16ed7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3ee1890a276269291d95f6f4caf582dadb19025517669fe9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h479a857fb9f54a7453325cff98cecd3cb561f58334c946916;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5211f2e59f1f4b606c2932e9f10c19ab4b08e5d2194487241;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a3629abe68be41b145d3516b209e8cfc54bafa88598f11bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb7383d3ff329d76512379cd1d0443bd8eb8aa83736d21689;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89738803591ac3ce7abcf32dbed58dd538cc4c304837638fd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5750e7c493639ff463f1d1b157aaeb7c2ee4bafe4946be9bf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h493b7b6e1ec31685f2c5ba0037dd381abb04729b68343581e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h305008b72e1da5fba23c905eee250d26b8ce64fe0e9a3951f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9853dbc4be17f7c66dc754dd235829995cc2533eefbe82c4a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h292d19fd3b54ae58b0c5a91f87fd93cbc7b15bc8d48023e2f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d4a13955b713ba155a32656583639d06db7311d335529108;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he384278e18ffbeff767c4f047fab8c3575a9cd41e0270e624;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb566d82288eebdd2f39ecdec3724ca33816264b7ca159b21d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha124b768ac3f63863884bebdd2e8b0c593ca820050dd8618e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h83a59d606e7b6a461d3151e129309c4f2c7c20685717aead8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77a2e5a1405fe440ca68f5476bcf9c03299473ae7d0b33d58;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha29455df5a1e6b838cce973e2c19a29da54a2d6ce393454ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7dbd82943842605a8c1fe5dbebbc252fa537f9c7cb67b8b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b0766b4c54effed58f855d73784b1a018fa4a9c1eab28337;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c4fabaf82655277ebd67491740941c88ad6228670026d69;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb270ec6543802a353c19bdf63b67be0bec072a634cb291645;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb19abe6e36209156456234186666924dfa1461c66921fc6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1662013f88e821fa2cf0e19fa23eac52e69277cbfc98a2890;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4d262c5309f3439df73881d221efa166be538cd5d2dc32cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'habeb4921de62584aa1ac9d608d31f5996a491821bceb243ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h55a3df2709642b8afa83023e4b46d3576c23af4be55962dc1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfec981bf063eebb8f6a8de7d783b317777fe6a8031587e14d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6bb510e3e5391a3318ee0e16fd83e6fca35bc1f699d660516;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2623f71f672dc036262f6fbf5e42fde5d3a6c8d7b9eb402b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b3359e74f2cf1bd26f664073ee273dd020337388f795d390;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13b2e7bee80547e6c8d268df1de3fbd89cd6546bdc4a279fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4266f0ad26118f0b42bb97017fe3c1f2808e9d2c5a0b6233f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd342c26922a5878ec7fbb59d2d3d99e20cb4355db6157e22;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6661d2d41c07afefe45b4cff9f84d3149ab5afbe0259489f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb21e1da8e70510f7bbd91bcac2191339f1450346195736c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb04586719f359891ea6b31856baf78f05e0ee6575e5247e89;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he263c6623d4eb92f36e64bc58720340f77c8456aec1d4c5b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5c890f52e3a64ac4c134a2403937636f645bbbbed9816b05;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7dcb0b2f5a920979784eb205b9dc403654b1efa5e88571460;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h561df538993c55db4dea50c4b8ccfcdaf1f1c2e6bdec7a401;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4d66efb33ea338fb294cde461720998b000961a3d1488c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h244ddf63195f4e54ce1d2834f7df4abb357953ac0aa4ea675;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3e802d2cc841160c33c98c0e73269a153b927939ef369466;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3380ddcf935f91de624d6e3d53233e84f6f0625448d02a291;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb279ffa89d134def3a497005a195c0fe463a665579881503a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e5bc24ce7ae1f643ba79d8bafc95c7b6c30e5fae22c7df37;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7dca8b45b6b6e982a72b574c0f9d3cd3c2751304265bb5258;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7e634f3a2c6ac7c85ed37706b8d8209de01812b775c392e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7f60a0b732017171b8b4dd338ba30900b25d573607ee93d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h751409a4e8e11e2517123a33af2c0313028ccfb96e184f2a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb69e1b50dbd6e8deae6757ca7f360a959ce483b4258c588a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f700e51a50a4bc0c0fd96e1a6f97bf8b408f5eb046b0f496;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha55c719b4f440a8ccf866ec7e7371f6d9388743859d5c1dba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ddcae1f19451dfb561364b911e44f7a7608827cbcaa45ebe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd17b823ffe04d7ef6f2522929398078a7c08fdf95d2bd116a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h467eee51672f5e1f4e3f970d6226ed7f59d587d7d016a8fed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab76098bce32f55260a38868f870487c722dec7cba8f1bfe2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc05decb3410e93de59e5b520cbfbe1a105453137569f26eec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h85a5e1b90f057e5123040de6297fe3f202aba8152841c5a7b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4cbc774c9db8e4c145c8e95f6558efbb2b280ba4a23fd5ef;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ef6f75b54bb593116e61a3eec3ec9f47c9097253d5ebe219;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb6672e6ce0d68f08c7b625a42cae573fd7abcf6869876461;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d83f512942e5130c749d3421509e81c971928d3073dc4805;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h417f2a9fcd4065cbd4746ce15a9b6864f6562c30821419f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54a9034f10926262cb34ff7949122dd9fb1981c562e9c18c7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11097413a455cfa2d44f5514d5412c11224d31b4f8be6fc52;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1f8bbaf7408f1828b9ec5afb568f934729531fa490dbb17e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b2524e672348bee7a9789e67f5e264fc3096a9637471aca3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h232b6d68774eb29027c4ba2bceef675a88e5827d0ee228eb3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86b5d812d6b4ca277233b64f2a945a9722dece408f107906c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd36b4985c947e5643efdc6de48ce2e298fc7bd2f472d06b8b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd450f6dae861e9f3c6b559d3eb5374f21622eb4c063f74c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hddab7886c8be0a5569a6a5f3178783c16fbb4dbac95fea0e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2835ee27339ca76d780dd2577185976083fa52de917a7bf0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8c3a062bc0e8ec839239209e93a3dca6b18877ac2f96a183;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1e39ed439ecca2bdcddf591b2d5fdc3f0291fb68eaffdb92;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f9f274c44de3379cd762b32811741a042a9c4924b95a4826;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h343c6483f1ef7f8382be40067c42e9b2a9f5fc5bf673493c7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbdabf9940983a6436c400cd168c46fb56bd0ac58fd10275e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8178499b1f59f321d217bb293f3954160c16e75fc5350658;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0f58f209275e7c93295f4f2caa103dfa3a859f614a6d6183;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb57d3f661edda3d2f34b29a5c0f6a2871f40695eb0401dcd2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9224936e0ac55363495fd1d6b52b27417ec9bf01ea1924a35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4ecb1cad733909c65e36913755f7ce402f5e72fade756eb7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ba2f9ef06b05fbf3eccd6f95b74081ccf7f5b1174e1b7a38;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff5d61d860f9c6bb50932774451b9cbb4f0699464842d2422;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc48affd5e34e51b775baf4f85edde6dc1713ad600fbc0320;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he24db82c814cb677742982bc858c27298c0dd01ad044ad053;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3c1ad037d7733fbca1b82efa4aa1728e6c8181e65bc10ee9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c205c4a9b03cf97a96a416f43558664d6d3cc4301daa4c2f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2500056aae27ba0bed9183e76b513f79dbad9ff9eb0153dc3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h43f9ab40693965fbf9ece1010b2ebec0d256f9ee84294b12b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa5125c72a9ffc3c53953873baaca24574bb1f5b3a14ad91d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e2319c60fe1d9db741ad7abfaa3aefa7ec1a956535237ccc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb90f6132e34ac70f2e0d583260245b6ea063642acbb925db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4319b51051e807166e85752a0ce845933665b3036e4cc0bbf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ff2cc19853afd049cbff4b9700bc1336b7ce701e1d30a585;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h394a3ad8398730b8b0ce404415e996778667ae46e3447400a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd41c28e041e84d1c280094cc9d1038ef3569b5e7916158d47;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha755602e05fb40ec81c918950e630086364e1e088729e88b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c2f27e40ca1d5faf04888a0da33f0e4f992cc540faad3877;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc15fb97beb9acc42720f33f8e1e0ed0fb752daee5c0d9775b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5bab61acac6bc56614a8f9ff11a0afabb6e14f8af474dbb0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h588e02356dce891311daa8bac158893763c7177f2e46bfc73;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd54cb78690a0305c4579e2b8bb146b0aaa5dcb56627ff91e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he24d529ff0411c9ff9e87362d3296cb8c9269cd1890bee7a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e87182826824777e6d163e7cbde27e9c701dca76bfa022b8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6b7808a503b58548b9cddc5350c8726397b31b6b3c072740;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c8c351e18e2dc0f03338806cad30193bf5da5c5815b9bd64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h345e7c3cfc98be55e590414a3cd6b54642b841bf02a34cf28;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7dc68d13efca64086d4c5f8393e0468300ad4c798ca09ca3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h512be7a60c8d002be6293bb5124c86e29b387aafed402daa4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h620da94cab4d934b31df9eac1b7f312b2c4f9a2ffb46f0459;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f2829f656aa804123751cd032a51fb76987f0e169ec14d4e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd8252bafd02fa91dd6b003097e9bde88b1db39cebc99bce40;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcfef131cf441c54cb529ac6f87dd525799ea471322f4bd913;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4fe82c960a772bba692ae2db9e93815244017c0cbdb737cb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63a50cf54e710338df07b74bac756ded5729a09665c382c79;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd09389ce31cd1e6441ef76ecca4e949416f28cfd3e6c5c19d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c2c98b164116160b78ee8460a028d8174a078a88823ab196;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f210ff737c005df861dd09556bb7aa8b4315c667cf8d512;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he78c6921b137007d730149c0e935075e57d020abd86f71111;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52c87494b6466c510ec998f8ecb36584ce3d1c2bb53635326;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he019b38e98c1b39f4e97b793fe43d14fa8078ca18e49f36aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ebbbe7b94d0d5afb842f7728ec57932fefabb662053e3e92;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h267fa07b9b523e9d1af13131e424abf1f27f4408faf3d156a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e78e790d4594260680dac756a8bd01136661ab65ac0ae14d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3487fcc1954bfef65654c44446daf561b39487a82a6636b3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a2c50105f858c405c8ba42fb3484be5f986a954f0125593;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7dafed20eb542825f49458104f2f77388173a40c568601420;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee7ef75614bcab18697127561054255dbc34a15f16403444;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e0ea7a72a29a84e9cc4118012611097fe3834a03c8f810c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb32725b36c3c838a53358461ee66a46721615d387b4c6161e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfdf6859a55dfb5b00548bdd3d0ffba55947fafc5924696ab8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89c18798beb809e4dc49a0fdc01e70a5ffb6f2ce1279ea304;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56e3b69d584d03aa40a38f17a10c723a11eb6e7848c03eaa4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34534f1ac6831a3dd8b194b2efe3de48569651eb64b3fc4ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1dff20c335f3e26cbb6d2095c4711c3b9b555d4adab681ce5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6564a63f64939a3fe151eabd945b5dbabc4aa1fe8e748244;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce3f921e0c051023795064106d1febe54d56695114e3c2db1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ff0de6b662e523087d2dcc1aa1e5a4285d735a5c79dc19f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb304e13dbe89a0ca2645eef04e1d0946d58552614583fea64;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a57990d5022721709dcca5dbb078cd45d0033c7fff810a34;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf32d63249b33d377d128b419a79b9a91dd2a54b54566e18e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha117d385835ee98e43b6faf0934349f62713bf03c994d369c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfee12fb49a49695036a939d41ca8ea7eed1187975334c5d16;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa495407c93e24387ad1d9fba83c0c3ff9ec06b7a20589379;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h375caec1be2ef16ad758acfbec9bbc04e26d9d0f5f166de1d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc008bdc86d212aa45f2eae4e40318ad9cc7759c26f97e519;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc64db2619b4a6accad854efa786a70f533fc9692a3653b95a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b1ab654014905bcd54a699ae10df9402454786957592448e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6365835021fea5aa356a9ae8bec00d34ba6d21ab47638a585;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b047251bb057c73e1f9458303e68c67a4d38f8acec816b53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e92f7c7e16858837446eecd8ab36e7ff3a20b4b670754706;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haccb25abce179fe24c6567e602dc88720fe13ac229c344c7d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee33109e5f9efd0aab8eb463badb1299c07801b6b5a6ca254;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he23c3527681d07bf1ebe611b8d98c98f5b051f38ee749c93e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h628fd0d1283011419cbe294b949c464646da0c7f9952bf3f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h397f9f7e1ca16b0ba3d727046980a8e520c3cee9b9da6dfd1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b1f9aff4fd1075c784da23dd3439c78b80db92a4b94a8d58;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28008a5491cbb39fe0f96c055a347c36b35bd0980a14f8914;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc255c4971a8549624bff3c175d0269b74f01f83992bcc675;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5a441b2de54ccec46fb9d0b84ac4cd8f78742018c0760c2b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c1b6e3c82213ac8b1777ac3b3507556e77e8c56ca6b2de;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h416a04cf50e6c860059947811c23650a89c99a94c525f103;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d543c834126fdeec8b71f518cbeddc571052774908505f4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6df1b6c2acaed3dd8d360aea5837992aeaa583965fd21178f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3af693cea6fae3a2ed1a06b1e7ee535b6bdd4af7b714e25fc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd5f797c556b6bc0405c199069336a30b9c910f03f5003e1f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e2d19fe4fb8053ad5a313a50d1b9fcc5397e1946ea404ba0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1cc0f963f44cd7173901ae95c2812cb717120210414586743;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13307ee4509107ea19ab58dcc4cbcaeae71423273244ae978;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h66f2ede2c6258da2045586ae2fd750cbd026d97045be2330c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8a118d824a464a5dc187529c5c65304630e07a90bc029702;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d23807b54d9c362f72eeb29b715db23a277a90136389973f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4b989861fbc5516facdffee04d739e3d0f6294e9b67ff01f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4de571b804f28b04bd5cdf10b542ca536fe489ec47b714e29;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3cff146c65f78801817ecb4bb68acfc98e8b323da95742ba2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb08e38058de8e1470bd71cba7339c144dd5b871ceb4b9aa2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3e85bfae53c184b889832f10b51b4eaca33fa4fa84175e71;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf884a103917ca232a82f8ca289be9addecc949dad9a9225d4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2422d4e8a84689d778b32a94e4990a3f2876191b513c2aa8d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h626b21bcbce65b1b6eef916810969d4bd788d59c792349db0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50d78dc3c415884f06e8ec94fa540eb90ddd68c6a9f8af076;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1cab83a6bb606043769146e041cbc086d8372bce51b621c3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6ecbdcf45a025bc8877767f5ea135f13caf83ed1a42995a2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h588fec74771d3c95f3d78f1b10a9043aa8c8b1373100ba394;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b6b5aeae0f17a9f9f222fb96e8deb1b3b46df9b395ce36e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h529d4276700985bf34f3065edd67ff1aafc8dda37daa5d3e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7513bee1a04aff6c36714326a901992bce2ad27a3d2d64a1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4bc9ad092b0f7e6a9298aa19757cb18626e7e2e679b7dd01f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcab0bb2ca5a44bbe34a025596180529dcbfd5205c3e0a9530;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb138cd37763c6701cb3801e2d88f0a540a0e02815f9f40c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec2d6610933b9dc8fb2e330b3dddeabb360964396e1b01e18;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3c965d87c0513afd06ff3b6c050792b3ba717467b5949ec3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f5433690823175a56825343a386465fe136d922cd903c1b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8866cf1ac718911a1c87f1f4e046b1a0ed36d0102f42ab146;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe4eb95c896b0ef8cd4dbc890d95905d1736a37c104f301a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3507b67ec29ada9370d0a5a7ab2dd2487b204d2dc77333a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f0da487666bec99a174ccd978584347564d0bf5e6c7c8326;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hebd4895fa62204839159a6e644b2a0e8a4c12cc54d7cf7229;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ddb174261f603000bf1e53448fbea05140aea3d8857449b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70d11c3705fe2b4ca3996936a2ac33c3428385540e5530105;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he02e6a3c32184bbdae28a8ae6141388d8b6559d16c1a48fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec408d736d144bb76552af8da72edbc624b596d29a7ab47e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3abc7091cb473378c14c321a55fb29d328509f08e66dd993c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7cbc32fe507bd08341846ccb0f3958ee07039218af8c9dbd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he281d60466a147b5b6aeb48feb2b3f0fe0c8ac54ed3156b3b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdfaeaff17cbbc36e49a60eca2c21cef9a0eafcc74278860b0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff96a30ed3a9b5017e45c19f46a44cb5df79e63a2a314b6fb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc88c9a6b8488c52933a4665b9382fb42abcfe123f2048c851;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc64e56b1113ba6e8f53a3d762f83102f3fca84719dc08fd1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e005c184c6b0e9619a0b97e5e70c992cf4e9c9e0f719dafe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60e42b9e9bb7ed4d1fb230621873004c68564455eb99c2d89;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c38506b28f8f82f8a723d240e2c80d43b73767fc5028f569;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e755b4bbca5ec1a334a20c07e71a87d6bcde0cdb70d45cc1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a1e078fff1ac72a5bf163ce1fcf440bc5fad1ea237f496da;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e33d92dc32b72b8e37a1a4bd70dff5ab8089ac71cd41f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he96399128e801001030c056fd4297d7af0a839691af79ff9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf027fa082ffa17305a83a675356bdf19d32039a69b479e05;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb844f9a184f50e574c07935179a94be8d515191bf758cf132;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7e2dcbebed9b1a819bc7b5ee7a01520efd4efdc813b2a14b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0f636916eedfac4330d937f842d0d90aa2cec0089de6b023;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h277ac72fa03a8e63458a25338966a9f9d83e545034c31430c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51c205e4e52adc16bae2a5abacd4a9685467a8cfe5c72b382;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c4f80d322b64adb40f57bd99919f53f892b7529f024472a5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10917e586b85853de19d0b1a15276b92f1284ce64e1099a57;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2df24ea8297fabb131ffcb9e121af887abed2cbbdf6959540;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab7dfcdcd22c30166d527fb5f132950d5b68fd00802cb2300;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35c1253addfafd915b4eb18bea2ce67d71ff9ad104d16132d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc161fc6a0890fdfbf145d3f410f4e290cbbeb237148f479a0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde4cb5e46311a879a69da5521ec861d76e074baed432836c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12e75c3f52faa2ba748c87a63e76c5d71809bc3cfbc10b721;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h488a2bf953aab85d6e206326c02ad3aca8ee046c6e047dbea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22c030e414f1cf669cbd2b02cd7d7aaeab9e5761444672517;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5ea2e45c316a9e01f1eb3244a86a1fbcdebeb2bd630cb2a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76d31c12fc889b4ecba45255893b98710c2934ceeb21f9c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b10914a04dc2e22760dd917a7caaa0c82c580608526aa744;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e2dba8427e83099da6c6876c1e109e4955e55ce310d79153;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb44441c2ca330eff6983fa619e5f3a939750f122bba2748e7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hadbfd1f2f54158d552a208b464522ff7258dea1a40bc5152c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6cde4c577c03360eef2dfe9f727fd5441c1d14010a85faebe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h757a5082e4bdcef5496888a9649c2d705d2d20abed0618490;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52302152dac66b986b42797154d880a32d15178ea91003fd2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1077fba8081f26d43f373e730db64bf9fa42756c71ab9e5d0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd95f16ed5b2f091ee8a34661117bf0d33522cdc09ed07973;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8fcf87186a2016f4d997bf9ac6b469e97ac4c77eddf05328;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ac6695e7f050b4c8fcbd037e1861430a8f427b223281cecb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c92ce7fde386a5790d691de5ef97cc0d7c42d17cd896b6aa;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h241c8124169efd74eef0038f77f7d1392604d8310c994aaa9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha4b8a4db9d356a8d272787d650c513a75ac6e676e91488389;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b54805ef0ed254d57504a80a0b9ec47b8dd6ec465e11b25b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce88ca05f7dcc5e15abcf6940c44c91ada33edbb1e233fa16;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd3b799fbc761f0f11495948d8616d97797c3ef290d181427;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4cd2ffad8d94252b2d6218b6cf44b40c032cb3bbc4449d45;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa2d436f1eccb7ad09efdd96182d455955e43d30efa1bfeda;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha747abb687a10c97afbc50d51cad83784d55919033a4ccef7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e0f8582672c175f3afa0e450bef13c8f25155972d2be189;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37ea6252bc1a0ad501511dbf1a5c5b010a513f9ec1ced39f5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hffbe900345edd6322af9a3ed6d4fb20584bbd1bc06e12cc09;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7754a5d30b20db68af6dc2676d5b3f6f5a4e8f1c86d8ac1f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10dcbbd6e9c45f1e9a3b4f5346bd9767a0ad933b247a47a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ef774c8776a41a458b9e2abd3d63ba61b424cd3e97f215b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6cb7269f66b5c009ad954fe4bc1346a42032f6d994e96546a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9623c132ec8c3628c299e62934516188034546714de024f5e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h331aca84e6265ac7ff442c92589a723b7836dc728fd236af3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68e51f2f9547b6a8dfdd6f6d8b005bb907b4b8bc4f7eebb82;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1bef82ac4050b5c066df7947cc20930f64800f92ce7207712;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h493ed38f5503d8948ccd55d30c91baf5cdfdcfe0218c09a43;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5a45cc8f769a8fdcdb286994b48644d0fe5d9e72a831a055;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61d6a31f544afbf6d85774721dd71892278e89d3ed3184ebf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h437d8f997d15b3bbc7b788e9781909c49a35685653133d7ee;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h219f4154674c0dbcbc3883dace8cb88d99b90b2dedb684b1b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2c7f01f358c2da7248e8ad7a20c1aeae090deb4990f8b1a8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h384d6953ebe7bf6d762c42e24371cebf74b38e631b1a01950;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9df2f8ac7f1747adb459bb273a0e2d716bbbd22cee4b5c759;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27d6c5038d70e20f8c0836a28ad1966efd7a5f1908edabca3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6b0cb61fc8b543c2d6b680d9a1933f7623125682e14b64b2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h385452644a227c62592ffebdba1faea061060b547ade95c18;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16b7128ea144e5ffcbdbfd0937a97a69cb2540ac781c1283b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1076399ba52e67e1d89c8862b2422ba6744b1e6134be3c19;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h444c15a2c86364c16e656098741e0d6cb407d2476845ea53a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6abc2a4236611ae9ab46a22f95600adf6f3c6af24b992ee5b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11739c5bce3a94c4a8c793ebee5d7525af6fdd329081e7ae4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7213eb7b53669f993df3d0d6aa9b351877641997fef696ff;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ceee0f36fc85aa805d1a4f7075d1723f1388d9b33609e107;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9bae7db41bde66c6bba85da06966455fd2927398f9a5dca07;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf107410ba65e666bbd6afb1c527d27e91b0ea28f303ab0101;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heebc6101e24bcb1b1d6e6e31070321da19d2f5d18402b3829;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd073362eb322591d8959552ad8776a633f9a93807b7dc16df;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h91ead2186cc1ded3df4e2c318f7d72ae55a6ea114050fdd84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d8233ee6249299154ad80220007bc633d1b32ece5de7f093;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1fd8aa637797f1bbfb5a70dcb0bb6270e89d44b19f0024153;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4c2786e99e935f65288bbb7b01ed03ac7f8e60fe5dfe84b5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b13eb029fbc3f991b29713122ab4def4df101a2cb5f4ffd4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69707680c9df903e36bc7635ded2d7ccea37b8d425465a5c6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heefe3f9c1bc14856668ffb957eed941664563b26bbdafabd5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4791faaf84ef63573bf1edb9dfecef259f8fcfb7c676c4d58;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19d69810e3d4b44f6df3ce856b15629053c2d83d826869114;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab398dc3b9a270b299cccae00de0e5cf36aeee24b8c993843;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a54583bd3be036f928265ce4e7e9d45ed76efea086f3cf97;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h291742f9767eb407f2d1ca14f74eef81ece63e242a81d9520;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hffe5a3656cd281d6ee55aebed6b599166da5248cadaa54373;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h372c0bfebadb765d7a6b7349c99e6859f5704fd2391195505;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9bdc9f8909772fb59cd6bd30f4ee8a05a1d1b9632a6ac998;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9e5621888b8c13c7531e080334c624afbf6b350b09957ed3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f9e9594e0c8107116fcdff1a1703552ad62697f4c61254f6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50bb25763fed3bb3a0f74ecd42caf783886637c0800d535cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ac654b257cf77dca5dabf9344e7ff5cbf2d9899022a9b308;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ad7f3d47ac62d67cfaac28153f26381a62ada49c33822510;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcdadc7beed4320545a131bd2f250c75783e09c070b5ebe0ad;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h822a6764eeb73b05489bc1b5458ab00cdbc8f3c65a8133698;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe9ef323645fad31720f29b5711b38cb4b3897cf2b8054242;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h442e92c6ce9b9423bdca04ae7f6526f5972fde0e1af29f5c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h127817baf7db91d263e79b37b22e681225ee89fd7ea90a6b6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa0e33d28377f4bfe62b5ecc0e4d763dbd978be071b83bef3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ca5e7661af592c02857ec302f796c70f3c0952258254e7e4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa0a82607734d4ed7fd81a66b055eba0497c5c53821c52d75;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6fa8525b2fd916553adf5600db7a32332f39d2df4063fea;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf63e398c3e15df75067e3989312de6b6a0dc1e31ec60e4120;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd497498c779c5a7403d1ad42e209829f6726792bb68d576a6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1866b03d7205a0af34020080cbb1e90612ff34e3cb8d9ab31;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc076fdb565cdd4a347e06e74991778e3d01a3ef80fb84dc07;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'headbf57be2dbce4375fdf1200f4f660c21a25b6a9e3a05dba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71c675f0389707ca85a433255ddd3386df05c013345d7039c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d5cc5d25e5fbce2a6c75be9e4e87fe9c9480f9b33dedeea5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32c7d0a7be8985877d8feb705cf26a9228316e16bb241766f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e45ec3ee3bf3f1fe117ed57653871892bf00fcb33be25ff5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had2fa8b1cb87fc03a65cb678f78a3ff185124d1757dcd2480;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ce03766856321f459e4e6b5294708482eeacc15fc840720b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10438b0ee96fb4d4a584acd02291056e0efca3d9a872e5b35;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe7b590ac87539a493b0fdb04a2544b409e2cb380b7088ed;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10c4e0dcbedbd7896cd8ebb7575f44a9e739c0b6087d39d4c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44916a054e6f205b3fda50c33201a2a7c9125273ad00231e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h516c9aabaefe3dbd9287e79a3be23e128051201e6f319e4d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90b3f5231c26e99b88775b155b1b597bbd30f69aafc709526;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5426c96025a82c2554a43e372cde84f327582b47e1ca5223e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9cb91ed55e186a85d0133130178a3e77ab5a921cb8f256d7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9e45cb4d21b9bdaae0feec5e51345250891b7a538a8e3dd2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd17632b1b8112a9a858b536283e6af20bf446351d40358578;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38aec67eba32fb0985d13313f14732a046b1ea8a8899b4779;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3deb1f0ada8eeefbf17547168be4a1ebcf71ba99301c796d2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha38a93b66877d1ba5a7484ae9dbe5084049c0ab66e88fffcb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf45279fab86b32a88e6d9a3b83a853670bfd076efb270f4e5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5039f9dc3515595e9a401f869af7893bb6917003eaae9e84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3da3baa2ff50fa6c3bf3cf919c684cca94fefcba2c47b78b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8972c0ba775efea2da594f5a99da81b9d90cbbd3b0d924409;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf62664298b6ab2ed6cfed576725f58ad429ce913c615a6b86;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48039535e1adf442abebd4746fac7cb76922d4817cac82e49;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbcf57d324e4484f6253ea3ab9791a4c0b5ee6cc660127ffb8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h379ac1a5ffbea6c1be53603cf83eb41c4185d91e7a310f8e6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc9e6a71676da25e4ee0bf7dc9820052b182f0d2d71274e7f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7fbcfb5205a7b0e758da32656f0991c5bad139429dfbf8530;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h291ede54869831f486a41b7a94262adbe6dabef364485b5db;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59f9b297043e32d86da54800c60f82bb7322e889aea7fcde2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41c5b8e00e11afa6cab4395f82f8556abfdfed16a6fa8230c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha13de41d7eb9ea32ecb38f3c5cf5856d178b3747f01b1e0ab;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc80c70603224e09f2630f36c7e02fa72e5361812b9250df76;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h622f68b8e13958583b28903b92aeb25ec64441e6222477290;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3baa98657b3ae0d96f17655651aa80ecd9ab3a0504fa305c4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c872bd4342fd52b10cf88dc32afb68d3079e91df9b0bf8e0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3b2e2c8e73a8bbe71642f070a14f61e7c202779471b9bcbe;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21e80d3ac538a1ef3be714f902f89b27203af0959ef8a3109;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3823816cff52d44f1ef6e860e553badeeaf67bce28a7b384;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e383290c8a9523a54f223c49d44592526cb4f99b510189cd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0f8cd312e070ba1d711b174fa450db195bf82cc03b4c56d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he001444ea24ee24fc1707fa5ade85edf7f6feb93da88cee5c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h237cc71e71a0764bf0d5c2b0ad8e9722773a2a7f3525e53c9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb95a3b38722f7b5ef1cbbfd0a970b2bca292ab29e5900dfb9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9dcb789e7b3fba23e5721d2ded45ad8b8b243a44d536096e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a069bf61c3df2e441153e073c9f5f86766944847faf7c40f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha00bdcda5d9b39b0cd2ae820784e4e9401a7ed81bb5ceab24;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34b3bcdca6c2310765e36a2816e66fe02f0e49ff045e7545;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ba583c38c9d5126d32855a1baf008dadbb2be1ef61915ea7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb263458b5ef6419fdd9ae1d519bb8db313e66b2022fac941;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he334e481fa1cf89b11497cd2173a91d802bd4e6cdf1d89b84;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5952cd321ccf506fc375000bd4885c6603462b095b2a43c5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8145560bab21c9048f010116b2d9c08739227ba862462241c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf25d5c66496648b6a05af9694c73912216f8c102b61d799f8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc39dfc0457fdf7251da1519734c52da6e26c46dfdc7be8a15;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd89ae1446b721a36ab92f3361ac4dbc2620bc6bc77cfce59c;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcba51d4f9950e909dda9e76c5547ed08b2aa747e46b6cabb7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6eaf1795d1a9f126cb1232e989ad91b191ef4b570fabdc27;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5e0cc233061f2ac8693a890a68721d7af29201dbb9d78a53;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40344d6895076d83c03b7c7c2907e8b79eaa5ba00fb7e311a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c9f23132844ac23d881bdc26fd50b1723dd603a12d2484e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4050964864fe2249c54d0b5911d333c0d3f8502bd6385e94;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c266a9b33722e4b8f53e08a9b93466f8637c7ba2940e83b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77506b06979ee20d6743ca110f25a00dbc6393a997b101659;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6397b47bc33ca5aed7a25e7975346227514149abddf19896f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3625a3c928f72b77d11f61bb537a6db9b25da6d80b84e0ada;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a280ac4c200b529d7fd933842f3e19d054934c11b9e25409;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89b4766172c3423a73b3da1f1ea7afb58cbfed1b6c05d11ba;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf96197857ea05c85fb1d4724579629bbf56fef0c37e4d1a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41b331654432713a8f0b29b471ff03446442c4828fecec329;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52c84dcdc439ca0b5541675ddb459de3518d644b68171d2cf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60f26bcf3fd9811988f6bef2cd9059e5257a9587da13405dd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h91e5f27c1dcbb316c894480a1d736f51b9c080b372be4524e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he869e31181c774e59d71def0eb572770df19b683fc296fa49;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf3517e1c090a03f615da24e83464d15f7cc3d3fc8895857;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc3d8c537d9784bb09c6e87937695cf464fd792cf1f535695;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63d1b0228631c6ea3d35455dda223633b9599f70409bf8c6b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2276887bf2977566ada9125d05b4a95b85dbf05e27e3fa9e8;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9709e0cc030305b07cc3b7585d05c25f60ffc77d708ac96c1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha72e182a2fd9bb60d2210833b0257ae2f96488370276cee32;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h165d6193f2d4dd715acfa2dd969501228d6a2e3b3538b6beb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf03873066e88d92112762dc7f00804330dfdf4cc2c68935f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7098cbcfc2a15674d7579ad6e8d92f621a179693046532d54;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h462fd2ebdbea4760460bf5d2bf432407f0a354a6e8e04a982;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2e2b5cc1ae6a01c5d7ae5939ea4a953fb14f5d20e2921928;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h725a6f5a2ca9dfe766ad7cc07b53ca793026c91fe722ed1f1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78f0e35d324fef6930c1b8e53c718394f63d2b5626b66d4b7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95653d3ca902355d6c3360c947937b72fff9edb8980b66da9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc892596609be66490455c5a762b89c17b960de22d9f85be5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf5f1dc361a33d2d7afe37ed6079359f77dabf1dab8f93d0a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0e157921b63cea314a4d1e58bfa6c34cad926b5c1a94ed65;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90453f639fd97c158e66257f65afe24b0dc805934041442a3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6ee0cf2afde4f26f9e9dde89ba82efd4e6d39028c9feb12f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21152cfcdc361387c734e27bf2f9e1a437ee2bad6419912b4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd51c293267421887e4736b888744c30643842c40e71b8b62;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c62d086124edb562f1e5d86a958c949647801f4e1be67c50;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3324e1f2454234482c798c55bfd641e40025fb35dc4699bdd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce1303530829e00643d9a17f69a1f7691cca4ce9fada44a74;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93d2983f283b9b1af7a1cd12fe2416794578fc537c90a77cc;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h902b9a0f99f9f9387cdf2d9880ce5c3be35ae1c47900314bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b49adf50eda54ec0355c417d3fe67133197006dcbb5e7dd5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5878075502eb072989589d6fdc5dec55187781b013305fb1f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h838eeacf185d5d430365029bb577469f2c8cde05f4ac0a0ec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf045c85a9493b3df01683ba03dc3a2d376c356ab9d6fc371d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5271235cc982607c7adc6f503ca46e96d8ba32b65836b091;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h235eddb2e4dc107d5ddd2af3925cbd7344b5f4c90dcfcb400;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbbcb3a64cc5246701c0b85ed3927d34528466f8b8f5d5556b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e6a41188187fbb1a7e93d925828b70c735260fa0ea0055d1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29c1d9129ee8097d4537f7986f1da75d98fc02e42f7dd389e;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h688333925add26852af220c98dbfa738104f71e9f28e60a7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46616948d4cae5e0e96439a7fd158f0b97da46a4550cf6224;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h394780c0f0405054052e3450df99c80a388465e05b7fbb9bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8d1227b74483da0a85d08c112ec34911523c68bc9867b4ec;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e3b2e44ec6b89a9155814b90a63f32348dcbe2c5704ccde9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h836e601db6581224d529c55998b0d2f6098a33ffb64014b71;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45a6e036b20bddc958571dab3cea8aecbb1f78d0cbb46fbfd;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h55489d008770e81448c8f04a7a3e80df88eb3fcfbb41e3ad5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10d2d769894d373fabb4dac196bac1e4434d8065cf71128a4;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d3503e19e3e74afeabcdc5dc94ac7e20bcff6439db4e08bb;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1c2016dbdadaf6a6e558f95be2570eb5f63efa81475ff023;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1969ea800c406287531ec64958c85c3b0fff4cb4c56aea8ae;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had746477110a994a00c6a795e886329c583263841168e8be2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6feafcc509439db4d0c813dbabdabf1a5b319615067c9dd52;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2bd8501dd3c0b17e77e9d3fd6bc66c0ff208e5e0633752755;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf1c8efda4831a4773c727e850cc00c482f3bb3c26853ca2d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2e75aaf70f4b340258e10126338a9d8edd6a5fb7080f351b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he208070b71e6c3dcd228f36a13e78a75de190da51760c6d9f;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9537469672f41df2ff6b57878bd0af92f45cbce3994604291;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57908f2563d471ab8b03a3838d2cedfdb1601f7f5d2f9aa95;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c0f80c6cb4cd27ca0f61f921e6b5091099d17fc597f44a99;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff64463d3c0a3340a50bde615f05d4e2debd70a09eea0034d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8b790d1bf19614bb7151552e28bde61726527ffaabc06d59;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbfdf30cf5275cb18487659b23c0d062a1ae23dff4a7d25b56;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h36bbd5728ba8dcc4959c7a6b111100d0ac5493a0a5b4223d5;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ae89463a0ff60080c486d9cde6f739f3a3946f828b75a188;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21023fe6b1c4dc0e6dcf227fd581cc324974da0dbc35e7285;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0991acaedf099624d1983888f2555543a7e9be9f1476ec8a;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a885d4bf91abea37e45f164b983a3a547310ea10bf9bfb82;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b62ee85c36b724727e18350050b2ec0b8f815e9a98660ccf;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3c8275aca83e6eecbc8fac41e480caca76be3d0204281476;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77eea9b259952bab28588d1ff9491011a152b9718dcf96648;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8529626364b39ae7c618356bb80aacb2fade3986d641dbfd2;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e7f32d583f82620719abe55d7ec4a33ad8b41b11f4266019;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ad204bc12d11c873303e90758c44f8884e2b0841a32317d9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd78113efea8779c0211d7d3a3e659585b3b35c432b19be3d;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had4d387afd7001de519482e0c82b41f0af6f232b27d31c80b;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7348a090eaf88b0b0b2a308ae9191df6e64782d6223b71b1;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h789c59107dcf2b028a3b1aec67b1703cb8b6f3b0761b9ff97;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0281fb120d03851461abfb064efb0401f34f326fcbb1322;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51dda602cab23ca91e90fb4855e21cb28d81cb396d70b8294;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6c2141833e33c1075e755081af3a96c4833ef657db6b8341;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9bb738e75685b67a78cc76a4d9cff7bfdffaed06dc2c85e9;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9897a4ec7a069fd6dc272b605b87965e33f2b7903a2182046;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb4c5cbe735313f8be857203dd33bd087403136e0052b89c0;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf928ba20942de8cdda94156b9688e2d049ee9425929645f7;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38e6363d2e6f45d0410fa2938d7795011394e6d696584eac6;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c8a41ecd34985ea4b9d323403def4aa1f002be2cc29e54d3;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d8b1c5eaae0adc2e476c0a2c9622f41f690ab93e7794aa04;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94ffc410dab59cf8a356ac8e458d6ce9caac0e16888dc4a95;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f526bbf51ef378fbf5ffb1a22e1a357bc7d304e0bf64db62;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49a35c01b8fe0145a9d80083bf26b7a87c17cd578ece55059;
        #1
        {src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4e9d52b1597d0e2a5d8cde20f1ea62d171c2958f4fc9cf25;
        #1
        $finish();
    end
endmodule
