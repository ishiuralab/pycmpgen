module testbench();
    reg [15:0] src0;
    reg [15:0] src1;
    reg [15:0] src2;
    reg [15:0] src3;
    reg [15:0] src4;
    reg [15:0] src5;
    reg [15:0] src6;
    reg [15:0] src7;
    reg [15:0] src8;
    reg [15:0] src9;
    reg [15:0] src10;
    reg [15:0] src11;
    reg [15:0] src12;
    reg [15:0] src13;
    reg [15:0] src14;
    reg [15:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [19:0] srcsum;
    wire [19:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1267685dc41e051b6ec28c9a92c4cc16206e20fa42e39c1f12357e00e709044;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ab9d9387d62e41d1c50ac1c61238c06199e36b2f1953f6bd22ba351e42b431a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h367e3d5055e5e0c65153bda569a1cd795294bcb1a9f9d1b3ff3a550a514d7110;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60860639b76af67e6578e3165480744395a161b1d522275f4139906965f45812;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hada663eeb8d3e14fcb34afe6556b6b003f86ac3fe4ad6a8bbe3b066f32586bf1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hba3f4b58c94c8aab8056f67db02e39a22dd94eaba42aad3926d574c41212f419;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9bcdea33d1c6f9578bc03aacf9acf9d3d3b09b850f2fca26167850ac0d3ab953;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3784b5a3b19b2fa2987b51c636843a12e97364331dfd44289730b57c1c682140;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf2b51e6888ffca95704b18f756bb1972572335e4d8c10c10e580fa26aaa548f8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a53bbcecddc40b4e99ce07b487b02baefd6ae3357c0a114d132d4aecd8d7a58;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac85395f2bea17f1e85ad71371ebbc43d3e7dc414998413bd93c739a7032de66;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hefb015eae38a60dae68120c5e6e93e16ac7c4f8a58bd072c6a4212ccd8a8c482;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6903ba82093e0f6b690cc58b06a4493fe88bbce38d0a9ee957aed0602eb710bf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd8b8a6d121029db2fa2e0705c64bbee5600e8061b9aa9c6a5a900d88e61b78f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd4c04bff7fe3cbd9016bbe6222ce8ee920d08ee186717bab0476b30ff1b8f337;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc71d8389a0976f72fb1d7e427efe9118d8ad1e3ae0b4b8dfcea710cdc8a7c2f2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d69e06e659f769690d6f381dceb0a6b9cf2ec30d15bad799ab2745393ed6c03;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he3e4c877b53f030cb841597bf61aef1c74f9f8f30beb0b6705fc60a21c6cae66;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h13a9d18786258bc987aba0b4372053170fde5b064e62c53163eb45020c36dd6e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7c53b62785885965d692fb9b6f9b3cc782a9e5237f3b2817dee1edade18e4ff1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h498b8b3e657ac5989210cfbd7820a05e29a6e5aa87dc3b3b529f2fd5eee7db32;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4774c10eb0f4c6e08b827c55d90275be8c64f57bc6fcfeaa99ccaedc21cdac3a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f987e57df467b9856f95212004bd07b5a8902e5b78db64575970220b3d26fbb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h82f071a01e3be2bc64053725ca3be52eb7f50138fee311527ce93ced92e3f780;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd160cba82e718c643d7cc7cb2f55de03443b60debbbf0fca83ca05e9c864237;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ffc29139f651dcd2ce65c050af22ad28583a3ec347593ef81bd4ca32dcf802e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h523ff4494fc195e2cb945e324e3832ba3e08c495578213d9dd443a785b64c3ad;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ee676780e027c26a3516b42d65918a8ba4d30bc5df1bea632797d52e928368a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h175cc8b0411bce6e3979b3f996edf5d690da140eea66cef2a6dd0a28b0eab0bc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7e50133c0fef4e61d0b42d16119633c23c90ad06c7c511b98151c06f399d0e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he8ec2ba3cbe0c6bc78e7496c0069f5cbd43f051d73a50d01948c687b39811f9b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4467893b2fa80c1d646f0cdb14262a4ffe5a73ce036394e715e7fecd789bbe10;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h68c685f6dbd1da63111e9f7754852831bcd6ca760f85b0fe1801e50eb30dec3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9510b0233659b2e7738db1a1a2d1d28d5a5139852ebc310ad07a0ff2656170ba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89d6f62f86ccf893dfd8bdbf6b244802ee7f1dde190ea6a073c9a67aa27e8093;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h65b536323649bbbd6b8ac23874ddf560b8cf3e44d85c5fb3169ba372f1c63201;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcfc11360b6f5e655315ba26b2be27acd13126f97177d29693ce1c85e00f98b41;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb0fd92d0ba63b07b68f0d66c202c11417ee284937059cc1fe098e90ffeb0257;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2500473b242c264fdfd52813673660da4573ef5435a364dd9d2c345c7b07f920;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f4cb02553ca43627af83985bedb17d87b4238045ea8e28a53d3fbf459703d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0196df21faa54d8b8f81d5fa2f9355b8b8f141853089047695e0a6c90467e17;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc0c18f614737eba9db96de1f2791c9bb9458508eaa73822caec2c6f36b45542;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9b7265fcb7cb15da297e018aa4e68f19a3f90cceebc8b0ab82ae846ce14afe51;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6ceeb9116ee578c287b5e3c8d68eb9a5940df02632977319f49a43fdd9340a56;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h97290ea4c5e9a986ea17c54ace13f976813edb52da4037cc4de8e34a0a6c59dc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h158fcc986ebc1ee7b636392b5ea718118423f3e3ea79276cf841d0e84d18611;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee6ba4f44a2926d96cc21058797e63b808722f29a1a1a0a188e49a5651df5251;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6af31c86e0d6dec08be52e9985e1a1e26e3a1ce9aa3be8a390db3351614d350d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf4d8f77ea943031f453b52e1121ed7bdb221c0a5581761002bc024a008d63fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h828b337bd1dcb7042b34167cc5263fb46d613f5ca4de4f274a1b5b4480a0432e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h210abbae6875e554fca61865d76d16fbbf9814a970c7345eb2ae98283b1aa1b8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h87b6b3032db59de45ff56febbd7ae1937e59f30708b45e8337198bd00caaec48;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hafe86b7499ecd6c27828bd18a8dcdad2a6289c2f7118aa90b808a25cbdaa117f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h35cc2152abf16b144c0caba1ac236074acba249d2caa403a8d986d0e4588ea85;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hef4160dfe7fbca7839ae1fb67003626cee2fd67943f36cf10067473929152719;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he2e32eb9d260707ce2375e0caeb4318353dc676559b34babac9c4faef391bbdf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc697853a8c3fd6de0a94e26da67187f571fbe6f8c5d669a2274ac6ad51c606e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he1fa9b9c3dc2c7bcbb497dec285a0ba65618eb76f502a9446382ed1da8eb229a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a91d911086adb560b8629b8f7426e1a9300fdbd2b1eb5cc246fe7c2c9362677;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6fe7204d7a1bffcfee169f7f9671b7e1abb2bf45a4f9ea8481c8c9e9d181898;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha78a45b3cd1b2c80f546379f5c92ab65d4a4d92931c89fe72979ebbe39485ba9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h995bfee7bd32a01751b911687f1bb4ed25a2ae084c50377f5ef8a7fa68ac00b4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h575ae22b5dfd5bbb80315dea34a33ca60234cf1a2eb8100a79173de5f05b240f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2aec7b53e787114f2d7c84c30389f92b5e0d0ec6fc837f628209a7de35e27fff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e5e084161b47b173712f3ecefa970ae09182c2f61a0d6397bf81d70353e3445;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h536145506fb36b886b244af7c4558d0ef6c524a67701c887c6c588fb4fd18786;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f4f7c704f78c5fafd5ce7b041b127881853bc42f64bf8e5ccd13eec769d5a83;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd507d8e10c61dedf1b4612a4b386c2431d38e3b0f128c26ba7a2ed17ec6eae0d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7861a9953c20cf059296c091a5c64a9dc46075836dc3875237e9d395f29e81b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha3c087463fc89896adefeb1e475482c77921e2e02c7fb1d9ee2b611b0bf465d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8f14845a08303ded032b7888249f73acefd07876e2621302d32b0fc59d0db2dd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23817c2818361c64b4a9feef6debbe944f2e4cac841adb672332b252260b44a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcc2b21cd4436b6b039e554e0965809b8755a9aa13165d482ee2f0646f0be6290;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc710a34394ba4e2dd9b579b3ce6fa107402569b190266c4316cc2094a231d535;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a9adcdfb9a1d4445b4e4f9844a692237c82e813c45db5748bc58937ee4e28d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36b13933fb34f32b4748a7076a842022cc092dedb7db5a36c0b2c08f2547a864;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd3942f59b30f73834b8c08e03616e677abf64d892d9962afb128fc7285f4e038;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62372e4f43ba15b76cb1f46d6a40918182eff69d4ec4ee479158fec6360221b6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd703a43346d4bbc7fb496b568fcedae2e4f1c2166c69ad868d3b19d94d1d929b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3d20e5b5b468d3b06428262e1ecb706ab9260a0ec05a0e7dc7dd2bea14ae7f50;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc0e3ba17b44abc47a477236cd67f06627c0af1143dff184540d689376a32639;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1335b7594f83769433b597f4a38943e083b158bde0a95d8e8b768f25f8c77e9f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8449e3348fe7558ad02a9cd1e75dbb7234b435e1a33febaa9cc46b2426f613ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h442695f2f10fdbb25eacc75afb0f68e6601fa4d3df43169d1f034cf59c8be238;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5190d60d1825d555c1453d92fbf271d6ab98afdff266665ceb44f48ae892983;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2bdd41623a0e68c16592af7b5316117796fbdfe349b0ac141909ae55b3e3a791;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha5e112771a7eb9f49b01c1288d7adfd53285c3fbdd313b8f2fe9a585ccb6202d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h67ceb1c9d24f0fdce219918ceda8a52391885007b7f6c62ee5ec5347ff7b4640;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he0b765d9ad93923697ece60c11e53fe3c149c53ceef109c8cef801d0a7d59f1c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf72794cade900d8839743460502c57a82956e86927dfb2a612566c921596b442;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdc289ef8e85c6253b24ed81e1581fcab1b3f8b8ce8f46406088f70ef3075bce1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ea07604ffb5812835a325f34778ea3f92a9e2e4fc31cc51ae1d37ca99e2e0fe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb339bd51065f791b9efda7ccbf43e872ffc434e1dbf0135c7a0cc6b7072eb949;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf19995f1ef1462ccb36457f073748dd6ef8c17c692a4ced4cf544110fa5edf81;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a68e6317917de6df2f98fd1b331c4747c9900a562e8c65bcefb6da41603d485;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d204752b4f6fb6ab3c05f1115d14a254ebc223ca161b5306acce7b891d41e76;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf55952fe7c6ab1b1696ed5d583508763e56859d636d26aa0380b0e47ca0e610f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h939a0390e44616d9630259f63dda9e9af722e05362143055e6c4f102ab51bcc9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h446e3a23f8c34696a73429076bf3c508a67403460f23f7ee3f54dfaf14dbf02;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ff49da6270cc2f36f431c2188f1b18459289f9042e9e92825e0716a3d8a09fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b2780ea4b68fefbd35c0d3c4c59703aee09cccc149f90ff77ac941d3ab4cab3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h25d8a4ae4297a9282b80b6088d704e4b2a225c32efcdbf2209cff42d1999ee2e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e952ebae0f5cd36a10f2422ced504f2aac59cc39d9ff727b30b3754861d33b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb72d18786da50f2167dc2cba185b94b20d8e1cd565ec6e843cf104a644502ca5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcc037c8c45c8adb0501512196639da2da7b016b270f47b4ece19f5349a600bb3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha4d98cfdf541298acc675bba6679f855829199908a6fedc2622a42faf7b97b6b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha89b883e5248220073968e8e06fc1417762de188f9eade45b89b93a949a24601;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb21ff0d113511ee31343d3d5864e825d0874b8e221c1fcee2cc8d373bd33b29b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4185db22c6fdd59913e0631830ced42be38abd267753e9075fae8b68a2547e13;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd946704165a43eee7a8ddecee3e9bc14ba2c9de9223f7d6ba7f65dcdd15f3360;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha8f9a7fc49d4e3252a6e85407e7ce250009d3ab463d9def17f0e31e76935ef6e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h64bf8a7698785bbcbc162242494adb6e54f3a6dc6ec8ea7a89ce40aa9814fc57;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6da0f138721e8ac8d3902d912d0ffe6d5325f57d86d144c52b39d2d3f45898e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec39bb1fb0704b25a139964e6d5334f4c4d5d526d5d3fd3fb623dd1b8487b9f8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcce01ec20ea803c796f329b867bd630aa2fc0484166bc292f705225b2788e511;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd4f81f8b52d533165b4a71b30d5e9a8c01d50d6fc634ceb081c8f4398e59af7d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8c001c3375b1bf970df7a36d67ad6f8683a9abb38600c835b09061a90ac2b34f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc00155e40e247139e617294728110dd4639f4deb3075e9cf42bf9b7945c801dd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he01d0b1c2c78742c6f0d886ee5402a36ea913f12720736e42c6cb400b98af57a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc6df82458c83983805b229679b9c7ade3323cd967a7500625256a9db1ab805ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hacf184ec3638ee653766baef921e4d6f94a31c2ff0e298c4028f4356e9db0cb2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17f24e719b6bdcdee3d9e8fad3067e19310895d775bcfef912df415b90f0bbbd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbff0535507f2e4862691532b9a891ad6146df0d799fd6213266d3dfbbc9f89bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb15d25402c04eea12ada36895b18c07a7adadaa79d9e449432bea754768ba7f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb1fd1a3464e22dfc97907d0869c5a93799022fa3dfdae498f02eda4defcf19b3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7618925ec0d5b20b3657d1ef95c6d1b2e8caee9ca56a4a7b93be2d8658da3091;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ce114c2d4b13619c85bc89aea59b294c544b07271cc9b01dfffbe77eb98203a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h793de0da5334c92eb2a8c85adbdd1c84cee2c0d8247c9e8bf87ccca65de44419;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd9359e3b6782d7a1990601982e1f59447572b7606727f0bba79999cb19725101;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7c6a8d7958887127e1feac42b3564757e3b58bda5635732e60e9ea0fb8f4aa37;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf48a84aa43f3b8588396e9c81fca592526674819514d56fa6c8226143a08978;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2712a924c44de488c0edd7fef6ef4956e5c3ab617e7ea26da1c17605ff151e63;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc72a52d71eaba7033c1b6ede99d98253a827654ce56274d5aaae627917d1b3c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h444f4b9b19d5217cf0bbe74ae43af6db37d260c607eba120f934dcc06621ba74;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb9d9344190ab7404b93ae667981a65260dfb123d95b0cc14055667b8281ed997;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hedc2e40540c107cca61844847d6ac1889c3d1ddb51745d5b7a4feabbde98e3df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf858e4f638c54c4489ef58c2666865033b2a9825b1c16a81dcf8f19bf96353a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha001214a54d55be3c61bf52020218cc807468a2720dbdc915b163ded1e9843dc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e5e09e65f91af5bf6881d0a23e84b636128dac033dc0051a23b67723e0beebc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h856f0a7d7621d94651a791dfad9e6322d34d2cfe548e60e567180f898a769300;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7824455d881c2386713bca8c6c78e04937ddb7f346f8921a46c68975a14608aa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h526c05a16f73146211dbd4d5c04f1289cede069ef78f4b58b46050a1bc105d48;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h663ad9fa628cfc1fd3bf38c8187885f93f836168cca2c2ea5d7f9be7c14da8f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'habba6959368bd1695068ea0e10c044632f6c55ef2671874511dd68e922333aa1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7430d365fae73816a3f4e8da204f644ebb71c0edb2470cb9521fbe1bba4a111f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb192cd21da71769a5aa40016fcfa589714df90cbc46508e345424d647ef3a24d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7683ea17e5728ea46d992d56c3be017877dc4393762f5616eff50a39d4d08c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5ae402048377554c65153c550f8261dc21ba8df2216fa4f8fcb4595d9adbefe1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hff71d5514e5df9ac26c16f776bfc585937004ef20a3c2df4f94c8e7a747144b0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h61d0a23ee31b62cc7627d1a2a4601f7d56948a0a852a01c5fb5779c5c36e0f09;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h755cbf5402d35e31efabafefa50ba44b3bc25d1d4165ac536aa45ce5f657d4e4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6dfb1e626d2b56b040d8316ecd75585775f279c7d878f975a2b5cac0af3bd35a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he345205306ded2f396ad3dd78f42c030c1db809cda89ec648ad6a4ebe5989555;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8f673bd0b034e0b676d22c552e17daffc7929b3c059316df690703e1bdd458c0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h90fc531348cf262990d4d86dcee9c46c2088cf55a11e4d08bddd7e007a96009d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb9a714d1f1492ee6a2741c48fc70d38b9d3e793284499188fe756a554d275b41;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h129e9cc6dcbe3b42721bce5e7b9dbe65dacfee8b29d2ef313b277b2de0ecaaaa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha5e8c1ed37ddd795e84db1358e0c32a98f8488544375889741aa3e69191aba5d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h94be4474f08aeaf899e300a1dabd9245b903dd62418be5fd01acc299f29fe6a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6835945173ce68b041b533d767de29020200329e17d180672b11ebf1eeace8e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcb569f05c17de1d9a4abcc9cc30bf4a00bdc35e17ffc599a9a038ccc826ce48e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h192cef6347d8de0faecd2231d49262024b6548ac65e67af973bf30b22cc2e977;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he9d68ca00688c4bd2f365bf73281231a29809810138810d9896006fad367e24e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he808099cb61111516f3d0249103ad64b33b8b6b4a5bcbce20f0cdaa12017ce5d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heab64d031964f412554799b26f5ddbfd62db69e2988038d8f5b2e446a8cf2a80;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8deca1ebcb9a19c93dc14a0de76048776234132b1c90ee86c8b4cf45636857d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h788912d824876cd6f418d6c89d86dbd331162dd209498c4eb091175d6465c162;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf48e790490295ebcf2406c351f9c7e1c3b9cdd7f0f490112064a48b0eaafffe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5605331d6077bb58bd3118514690aebd40342461d6edad337748ef81d043ad1d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'habcf636358f44ecae4cf72cdb5b7aadd6f56cc5d566795480ad1801f313b4daa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h66879c2fe5c8f57acc4144a74418a19e52c5929977ca781d943803ed519fcdcb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haacd7cf04c816e52cb50addf1bf751bf74d4e0040689021f6a40524fd80cfe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heae0d5b0eb4d6b5d5ff3f28b246bef6e7853e23f36be09ec917708dd3af3bdc4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h69f1cf2ebca2f1f26767389db34047b9086f3cf01b27236e51be875e17cf1a86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h95fc162830b0c49889182424c91e36acacafac8be2b12bb582eb6e31edacbd7a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8dc650f992be6760dccc4f5c78d0ae98d8a15cf30ed584ed6c4011df6b03959a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7857a0aead038a7b28b0f31a30b143903a80d0e38650b4c17919dd637dccf036;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf9ef562f199ad6f1f33c734f879aee8c07fa243f5adf498add02a8e13b7d9faa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9df1d54e36de567af93d5b6904263438daacce79e3b6ab9c13d0b4fa3cc4a42c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc907f889f83735d46e4c78907ee2a3bb0d4a212138e7453ac050d7e447618dd9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h334fe060fa07c06a45b6fdf8e9f94d5d3e7193aca50656378fa10e8af529e04c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce0838350327fa769e8d80d620fb7924a101b4804bb3db886f53a9fd89821450;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h87c4a0450e8da8e92ddacc8f77b1fe09dad7e466153cda419c45ebef9d28cc4f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5159b9a6583f39b328ae632d5a557eb361f65b940caa904c8c565c1b009e7f0b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h63d6c220444ddacbba98ba0140078ed442238e4045ed2c7263b1b3cd44c17693;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36050414b63f8c5887220d39ab983715c05907de5810963405f8ec2f9707d80e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc29c4836cd5fba43daf7c74a2a664da1acc677b9ebd06e26e5d6c98cddfadcb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23963d5fef92613b2bfc89438e96b173a08730292050e1fd55d3e90290021fe6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he31031ebabdb189eddfcde3e6436c42033fb3e75033b4a9a761a34ab07891008;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a9c9335e1e74439fb56d030d13e220b49deeb53acdd7fc8739558c515ff6868;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41ade0b71c31d913ea6675c1422bb260a1c2829da5c12611dbf11d4ccfee85e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9865db36c68e72bacfee1dc2cf966941f83ff4cbc4f699e63712ece40e67c289;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha861bfcc180dc7e36a2d430b16b312970efbee06f151c0d99bcbb5a817d1e824;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h170aecc0a103840602c7c0e316ee17f6757470583ef2896e2ba94730307df011;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h87225a49278b22c4739c20415ea3d118446e4eec85409e731b7589b9e775190b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h334483473c52210f7290c22871f269da0b95156eeac277f166537735fe164b1d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha63633c494584b27218adfc41a5dd1f668d33108c3d6d7ba7f0fbc90f2494685;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8c156402b3545268aa6ddf9d505bf530808a40e7c137068fe93765a4a4935dfe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77d210bb6478f72d477fe72f649e9fee732dceb1e849758f03d8e18a9937b151;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h564b9f3c95620623973acf6a70f33d4e16bbf51b9f10d7e690e8eea5dedb0150;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3a4290cc4885d3793be1f3d4fc6215d3693e8c38c76058483e48b6de9d202208;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5ffd436023936e83a43698c700cfc6cc1608dedf08df4b30a55f271ccdc761fe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h668b71e0c458a5745097d0c3ddc4f85efd950ce10dedb103dbdd95dd276e4eb1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h326c1f084a5caf9a76e2e2ebb6c1543f6dedb394c1092d71f567315e0c02db47;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h730956ea5397d170b55afcf592f327ceca1e5146e485fa6dae9f71bf94e34932;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2311e246913360d16eb0b783bc56b9e44dc3b6ac92344c2eee04363802989b6f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd919cbbebe0e523f7fc80dd4ac47b4cbf4194f9ae97865d0a1a5f6a1d8ae0144;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h337c3e2f7514da2d53e6ac8bfd0d44a37944af6a628b7da0ef94f7e60de515ee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc29142e532e4b07d8589bad77b72ec5f4a80118fb4885e113a95da9977bf9dba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he32d6546836f08cfba141b0a11483e68deac03396bb26d336a7f858cc017ade6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62a1f61f6c3ce09c59d20828ebe434be7eb8e7c2e9eefca08f396b6c51f07c49;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60d9b11ce282c8a8ed58eee4134ff184c602d00417d269f8746ee5272610571e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h94b144e6caba84b758af9316fca8c67d68965104c8ca5e2fc82ff09dd85d62cf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92f5350ae3ebba19bdab97367fe80f697cfe596e8511f2252466c00759e524e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he78f958ee67eb8dcb94795dfc14e49cbaa6c9c2f573d2b862b24a1fbac50816a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h704c7b30076448e79f5bfaddd660b5aa6094629d59699b3c83ebbe5d34b7fea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h86b0192a37bf28f9df881953022f784446f876e036d089e1de3f51b82bf2c773;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h65a7ba625f02d1595a7bf8f96bcdc8e5db8e5f1de7a792eec15e47813d95a798;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2439501e287da0c165f3738bdbc29cb16f620ca7fd7a9d534f8407c180488356;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha3b682fdd3cd1ec505849cc0c0789ba9c48e9a6fdaa64dbb6d23a7d5f11dd54d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h31a8bb47e8b063e5055cddac6d9f852fbf77865e820715d5a924d3ca957331cb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h80007287a0ccfb61b764b402e7f1a7b0466ed32efc523d41ce41d945ff41c8f9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83f6bb7f77c119abe062fb586de881b2709ddbb198f0c10fb11a7e311831b4a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc27a50ccb0bb646e05a904b68ba6667eefed084ac7b388646e7dff637d977f9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc749ec9b7d7a7685454114a045e23c546e23312237e4dd1c52fa53b286ebe695;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc4450662920dcc53fb5a36d6dddd7ca8fcbccab1837e26b311f33e6e8432158a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4569c8a905aad5eb5ce324fcd5e071a71fb5b5524ace46587788e625a67f8341;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7a4061d622a35312252fc56e8beabd0c8707c49794d5586178be7cff240ffd3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6eff70f4f9f083fd0b7c5a3ecd379a2ea6aa66d529bb5dcd4c5d7811016f9306;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h15aa43c4832e3106697ec3514a7dabdccc6bad92b9067ec8a89dbbb7a3cb1df7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc506535ee2a12acd43458d24155c035d905d8d7c1f88d45c3330c1c24d2122ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4b0478e646f66ff340e6ea4175a84640bcb2f9c8ea7bb5dcbff3b004ba4af099;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h12c5cb533c78293fec5d612e6512d764a6e40a438be46fc3c6b4a417b054ed2f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6d6f5fc2a4ea56ced74e38f81d73ce642d83058d2f138c49abb86640a1ce6bc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b080cd617a85422c3fb65d74df49781df6dc7900bdf6ab38cf65036c4a2f5b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7c718e55bcb4016e294dd44c764933c609297053f24bde4d441c61d999dc044;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41455e2342ceea4c54ab0a563ff38626138a22d558b3c20314abd7bc12b4fee3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h88bb593127797fb18e1be962e4258462623f778f52ceaba2ce53421ce0a69f48;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haad0de08b92739b2fe5f78950eddb5d2afce28c34a4136c03d1075504a322699;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6f519c9341a72e35a83dbc34da8a9369f6322d351c5bf60e04ad98f3f8c445ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha2556fc2684388bbae4673b61b1e2fffcaf99eada53014f9b2c96c258c8954ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h896226ebbb1d9ed46562a33dfe4318a2947e2e966cf32a921e056cdaa45e865b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3435021380edd7ea13ab35bd2a16d026dfad388e4690b6e80bf39d027f9e4d32;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62429adde9adba97210945476b1a6942d1acb73100bdfb9bcf2edfa982d16dc0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h16040aa1ba8a7df8be0d98c7200837e641b5f3d0fce957b491d5ba4dc1c3ca2f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e4e029b00b5729a4d6e7ab228b99d58416b6ff47e054c84a44776df8a0738a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h693958b93b7baad3a5bbacb726484ba6168b60cda8e76f6bdb26c5d3e78a0e8e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e0c493dc975bc1c63fc48a5feac99bec42e23050e9d2e3a91f54848628552f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9dbb1d0e1b4c641814647e183b7dc5557f73168ae361284ff8a0f35598ba2bef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5cfece3f525e91b5552bbd405f08d6d56d58de0b0afaf9c07c1aad5432119229;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h67b6fc53738569ddc7f9de8018866283c5cb2f89b41acafacaf0093b245a04df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'habe5a50c08ecdf3effb7752fd9d6ac094e9f2bef61dc0f4d42fc0d8e2b7f7e62;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he947f36157e929a97b3e490d8d34c768a6e474975a3bf6497f9cdb49acaeb80b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98b1378aed2e76ac66bccc21fd650136b0e225761c2f3d9f182ef6beb21c9b86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9840cabc57b1b94c30f351550e2634969be0aea20ecee60243de96e6e2de501e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h878f87e1b94cd0a1a3853400eccc4e242fc141a4fa5ed81d0964ae4412549779;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ae7e754e1e4a075544dbc15b8a9b67512ebd4adc9ea9692c2493f1e4641f1f8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha23981824bf7dc9334167e13447a54534a0239b247dc94b1be6d034138bcf3db;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h219ba0bd8bde53a098dc3a82a328ff6f1a04dfb6df096426b7f2b0d41f454936;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40eedc5c589697eb6fa3d21335c71137700d1d14da3b6e3dfb854a2eaa09f75e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haeca43cec83b53f67b5549fef45616fd13949ef324187908fe62a6bdb7eea69a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7f3d970c7223b623a6bc4ff56af6e61683dd76be31162975a560c9a67a9f23b4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h54690e73cdb3c198101276cf2b12163ac0dfdac64b2f77beecfd85a1c680ab8b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he025c16d7ed4eaf5b1d1e5651cec30a5360959a1c5f39c89d8ce0b86ee81465;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf393452d39cb2a3d054fe71b11a2c466ef8d9530c253b66766a0acf8d881d1b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ede80e14005bf3eb85545a0347b44829c298fdc0b35985063d137bb38545b92;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac294f632421f3407d29b31074ab0ece077881d4d4b365de0a443b84982d0a8a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h534e685035c7572429df8642d2613c54bc93ce301d8a66dcc1ec6c41476dc8c7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd4a27eeab962c0a289e77add0b04d1df7ea840079eb04fcc212ec52e9e3094a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h682895518ab58176e80a096a2a403d0c5e1849d540ac43f609d41fad4dd73df4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha04b3011da0d8ef764dfcda27306918ac79e28497aba90c38d6fda55455e76d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h99f2db6f670d3bc5a5e59413ad46e5a469d0e6ecc488281e5115f4eaa5856deb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he47dc7a9407fdfdb6a1f184276aa02d01a771feb99415030adb77481f7589e03;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf5d4830e3ea47098715019eecbb1984712517505b35706b7cc183fcf5e1ab357;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9642f89e80fa2774b684c6dd3f3ab44feb2af52b6b7e80d99e3318f62e86098c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd317f70268e9e2ab0c4613a3cb83efc261716991cc05d7a18526e591e5700be0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h193b24176a50061cf521314e88989dd59104ae12dfe39b479a4ad0ddd3c90788;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h959bf185c2ae41a7627abb153519dd18810d3f5c839cd181cd11ffb89bd926b5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hedb5ea9b8c569566d50ac0a606a60bff9b76c4e1d38a90ce3447f35577524170;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92a07d89aaf66104b09480ef543be6565a918107f509006beaea798701545097;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h145679d5a83db43ec1e597f34793c7c5fdc276a785de135bd47c0e66950f1076;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52eba2d0156c0cdd1a7473b48d2cfdd27624fa0c6bd473cdd64d948d124eb691;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3c40bb077927a65d7b5e0131dbe355e0505d2f1bf317d9f371c33e945a78aebc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4b244cd1f69d3fdf78ed3e27cbf05e4fa696a5166dbfb4291f15af8f32bd57f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2e85980600a7ec96ad018eb58f582d87b6c321ead4243410b4d586de676ab7d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2edf3fb13f13ac22ddfb02a62157ed88f362c143d2325de8a6405e92fd1a0b53;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a099594641f4affd24a5b3d366f04999d7f169b0a56e4f2b43c2c824166a0f0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdec80afdd94fb34efb15ee0d179dd8dcc223bae26ba42d6998e1a15bd98faf51;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23e1a5d06354c2843757c0c1238e2bb1d72caa8a874aa326b02386d32d7d19f4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h48923f87d6356bc8732464c168500ad1cc0161626a2e1b5842738e25a0ce90d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6a7ee91fdc990dced2ce976ff78cdd11d6917a9bcecad52212da768a5b6ca6cf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he39b75c1594790a55a4ae4a4e3f60f08f84fd27b908860e2ee1235b07e1cccb9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'had0b1d129007a5d36edb4c19c83b08f337570acc37758f2918767e8f1b994543;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c9213c8176069375f6cae12fac911779c142b2e49f451150be2be4914198345;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h781270526fd8138ee85c1b8929c8a90831f288d06f2f5f8fe6d216714027e6b3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h75483a362fba8a8fddf04512ebb14123d00cc8a07f374b86269b03b00fd79d5a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93bc6945ba50db95ffec3ed7a7e0e02b879203380f21c25c1dfbb52c09830cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89032da09d3596aa0043162df60f5a370677b450a11a17a391fa3902ff93f93e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9485fe8095d1f09ac72b07a17854e825b1ad850b1a49742cce18030636f5f2e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf89e95c289005f22ba3a9133bf3ba724aadcea268764fc9073ffba8bc7ebc138;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h27efa588b4a04a0559f30f205319298c86dc74684ebec0c1b28a22481af6087d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf95e284c302e483807151d35f91ec01d4f35c4fa75d8c9d3013c75752a8378d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7bb507ebe67dfafc17db264f2d7feda04e3028a4ac23c0e888f51edbc3a183f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbe60bf5926abe6f20c360dd87cc331ed09a9c6cd726fd56b3b08491a3796d646;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc6b8e63abbc409e8d397110f4695df7c095b7d8aeb98fa8dcc19502fd73a4451;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h44307f9ccef34e7b632884a34dcbab853ffe29794fe2c376ff054a0f91a1bc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2ba361dcee491ba175871436dacead1864374aa08551abb658521e6a15b172c7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b95535b67b72adc59ac8feb36722c0aed37b33705a5df6d1b7dc8dc1d33cabf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc1736f6521006c64f70e263f093037b2f7f50f5c266322f4e05949ab270ca5bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea7eda667f2a51a58627ab908a460f1a066df2c82a00c273319c22000e7dc77c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he0e9872e606c6eb5393e126d91486b877ff3ad4419dc7b7055e7c3d303930963;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdecfc0961ecb612a4a6b3f614b430d827a42df77d0ba108ff3ef2bbbad8637e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1054c37ce380bead7dcdb3c95916d12f1e7ff1f4bed1a8bff9bf08b61b1228a0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h14e011b33618dbe5cd0c4cf1afa18977f0637ad01015824b70c640beedf02805;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hddc7415d40d2dc9d8cbf159f34e22cecba670ff5ae63f9ab9077f267b056c9e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33901d132820ee28a3311160e0ec950a0c0e7b6fb9bd461889eb78d0da9d1d51;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4a54e089a1b7a4d08e5aceac11c5682fc6d3eac66004807be23d5b3aaa0a3752;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8474efb5fe53fc7c0ab5dcebcf26783b1ef7a5a0a561a0c9b7c0ce24d01ed5ee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9d31d308d8b6c3641d8099fec8df6924e70ee0c0d6d73ea9bd17ce9db763b661;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h25735fe5393d328f6dff1bca550e76f6d3cf5964a8ed53b4f97e1f280add65fd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbb33075ffa4d563145c9ddc1a3389c4741dc2af4a43cb930b3d66e6c6a679037;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f6ae735da3c8db0b2ae9dc7d756f68907069771cea4bcdcb769f47c6d201a41;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc39139f1095e84b5e14533e92f53783d8d80d577658a8da6d60e173a7b1f6bf3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h45681c4d943e1783ed04b67b8c5b4526d0b6cb5cc24639a391b4b4f09670cb79;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b7ad36bc81747e6a3bd141461b61dc8c2f8a012884fdaa7e85659a909834d3d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd3a7cfa17435140605d2e32623a10ac0310b6750f63fa5fbec58ee778e21d8b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3402290ed3d03aefd6605b5d5cac6ecf7d4ac3332d0d05b3e0d4a9efaae98540;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h130f6fad90b96f09309494330edcbf4c1e9c95db6a63053affc63a6c91a5b266;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h47bf2dbf05f6c708981189e5116a266f9f3896930831af7ce173087831b4e7a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd20a6ff99c6c95573e80b343bacdcb15ca1583a2ef8590792c6c22b45703133e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf5e470d95e18774599223433a0c2ae74fd733c2ae7dd69b9144e42e498573a8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h60701579337a9e5f95260cdb2202559461e0bfe31ad1e96be1a913000dbec281;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h73299f69542963fba4479e38f8cd2859baa1cf7fc384881bf71e077016e2e871;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd61f90d0bf120d79697551048c8ffdee9c7004c773508ea4eba10e84dca4d862;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h473455955c620004011e42a06ddf5c9d0a96f5c709c32835385ee8ac5a1a1c19;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haff28f63035ec79fb2383edf226bc1a2ffc10b0d1be75f4c25baf45d0b53f89;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9830a6a12b7fa90716f51b31fc7706dd1d2e1c85f261e5924e59413cd293704;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8cad2ba596822d2c90f06a0d14ba4414d4223c336f00e3f13d65dc0f9db6c609;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbe6b3ac6ccad88b65e08cbeb0fdf98bcfd64f2e7ed13bab4abd35c140048fdd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1b900587a5d0452e4881fb49167b6034b0e119665de1b24c5e0134b3a2c3e0c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h63f13dcd9b67a6df75869de04f19c60362674f5d4ba71980f68a3a17214835c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0fa41bb9f03c52f0f0914d7b24dac7185480ed8f5a5ef9f499795b8d47fe157;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b78e16d7052f124c719d4c2f433f9357b425ae28f532bf35decfb5b919403a0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb3eee642147c868b44a469fa607d32bd3f7f345d1b726df4c92fe56ae936a736;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7cdb630f20f958a1ef5d7fd6d20313fa9f40d4217b01e54461870059c18e8307;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h65646e4053921aec91f992e201057f39a38695c6a65b938b7aa99200ce4a5e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9a49d988e66bc6d732b0c0e1de80d0b4abace47d3332b7cf16f01c785fd0f24b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hde01318670797a3fe8375e6334c941a88bd286b2bd2335dd2db10432cf90d5ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h393e7771defcb68e4f2e87449a671560a98fabd70dcbea49c310ae570cdd4ff0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab8fc8f1c99fdb5d551c0854933b2042c584b02c0dfa83904fd36aa7c1d3e79;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd2a26412ed065a77f3f5749b1646b5066ae9bc5117c6c6845e30269eef3ba717;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb88fb83c10caeabe64dfed022a0cbdcfe163af6a1cf69d580398402a9ccc395;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h86b9ec3925bf604730a9f4206aa4cb42f5a74970c537c6f0d1d8df0d085ebd3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hafa7de2fbef8b27676d00c3fc8748ac8d019cbe5d4d833b2f99c58eeffe9a6c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he6c32de436d6a651dcab623a94fc892e65e1a288ea51c2f984516c9dc29f0daf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9fbd041ba11335a0b81503bf4195a62e97df58d5bae7b5b431e7ec320e258940;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h26f870776ace35f1231c771bd8ac54835a70fe5419bf5cc3d0b431d31c6b245e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd28b442e6bc835d6221d9c2d19da43a0f990f267d3f6faf398f334af7d510980;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1d918551c2e55991f978a29813a29e288dce0c8da498d1936883deada5b5036a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf099f984f89e551b69b1697936479b15eb23f4182a6df232939852a75b99818;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ede0307763c487567817c67aebc49103fab8ae6e73bd76d175403ec5357a8a1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b00891f681515e600ae397a6ed3e3e6f1f97e7f47ec8b64da3b470f5179ca4e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5c109adf26b44a6bbed66276e228c1eefe93b2222f876e6b3aa8984fd0d7476;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h55ad317214b81c18a661ce6979851deec48b684edfbeb7dea09ba72ce3e503b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9286bacf1d24f7feecdae33f4873e9ec28102f9db1c6801c00da704ad91e276d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcc1503968fa77fe9a14ec8c355ad10501eeba2496b504e99dd45a5415fe7d361;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea323adebe1ff535ecaf396b229b40e3ec267e5a28a4b5b12cc3568021d4d9c6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83cc0f7621412c071353986e5924d123074128deff2c91c3ca7558dbf4f9e63;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h78af04ba51d32caca20c996aa72ad60379f701c65e9abdbcfc16d8afeafe9d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h43a78f4d49d29a78916391d3628b993b13c6d9fe5a4db3f276fd9d434d47606d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7ed0fa9cafca1b16cb936155425d221687303b0e7d2b33925083f62651425cac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he85514a3fff6c3f6b9462b8ac2392d0fb624c6c1100159671d08ada872f783a9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b32f75c3290a27343d773f47af2d38bf31c06b2821cebec5a9ad5f5cfe1639a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h580012a67bd2f52b5cf943bbd3b35141e6905d5a59c5176cba7c2d8045c2b4e6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hde46b381b5109a6ed3aaa46e5a0375193a17559fcf734e89d009a0c38c9191d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a57ab8012b7a292cc7e443da83ae6bc9200667638c1924a2d4475787b107fc8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf63ba29cb6ebe2bfa6f1a0285f5cb32812c27aef963578458a9667b23b470190;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb89cc8021d00a8241621622385c6ed82ddc6e43949d02bb1e9f0760d49e8cea6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd9471c99019b3ba889851cb13023a10470088d83a56b51b2571166a813aa1083;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h951969993ac0b263658643c5dcca2bca2a396bdda2d8a0f41a7f35d33bf67f40;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h995fb6033ce2d69f96a6f4a05a438372e6e082cec04569d06305995d30ef5f5e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h647a2ec0ab6bf0a2aa742c73ba1888bd4c152521074ad6fae2819ef31a61fb9a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40ebe921101e4be6dcb792d958e79eb2e55338548fcbdfcd1510b6e0dd02ba58;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9b3a654a5cff7b762bbae5699a85193ff69d53de56c7e0cfd5e2b62c22a4fc1f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2d56f5ba08ed9462f294d6ecc21895b1407cda780c50a876e9258b97fbff5b6c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4813718347284ecc026bd806cbab6567cfb78870f3954d298f5870c7e48c1580;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb8c4675d8e92220a5e424c5dc9b0e291328791a0e63bfdacc0d343cf8959e6d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h846d8330d49cd50fb2eabeafa0a39f318cd9c68cf8689782d9b5684d5dbe6edc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f3ffd7ca1dd681e252421f477f131a607414a12f802188f7281f268a4547c34;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd1307789730562ce97d0ed3a554931f0bd4fe38312d484b4c55a9195c068acc5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd28ee098d1299ad2825f089d760255804aaca6b940c2bc5a20c479a0c09b66cb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f445de946b454084efc037ec5da011152b49f41fc28c06b896abd7af3e06880;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd02cff0e0e6906b8e62c3bcca2212a43e5aa7816f7eee5f4e828391f51c0d42a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37449f382818a9e47d43b3c688764f25c70cc852ecaf4515458edf9ea5ed4486;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h146b310c70c0388b77819fd60a50d6e95bbcaf0365a3ca6f438b25863680b70;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5767aa5b46e162d8d003abdb571a5bd79ee3d9e1ece164c2b5c2604381dbd846;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4b4b69bb0cde3362f734748aa514b9eb327daad062d68c76dc46fff115a6f25e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7fcbe2ba7e69a408de19bea629a506287586ad3d03ca0429a6079aba128beee4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce1b0289757d4af1b471f88719c335647e66e4cd3042550a14a3a0fcbf9be80a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd4f0875da01c4462b82fff08cded9388413e99e0756787da24cc5809d75b141a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e4cf201ba9224360591020a0ef9010c96a3918b71c9c66327bec02bcfd79cee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2021e47a17048d3ec2039b6df0625fbeea63ac6121c5d728581ddca6abebef0d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9e2e857580b2306091ea5a65b55eabc7b1816b374fe38d92508ddddb9646ff61;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3d5f534638c4586cda38d60f9dde10d2425c9a55b468f65c7d69533880529834;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf8b603e12ab6e52da914dd0df1263a310ed07b0dbc4ec37545e2498dc2714878;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7db55882014a567193364db2d000e876ee697bfdab40f0a456cd4c209a0ce9e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a73c535783280ce1fb69ef46cc1fb6798b282a9c6e7f0cd66b45a89d2465f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h49fdc79081d780bac8a2a6d1ac8ad8bd005ee0b83984bae8341d30a04e15bf4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h444a04788bc5b030143b712da55784514a9e91408a3410b8cc03369a9555b65d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbba89394d515daa597184d1ac33581f2464482384a85cefc4b811703b803a014;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb4c8177475d146564eae33afe4517d1b00653e073974d8915c461bdc8b6e83ef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b1bf0a8a3d63a68c14fd2ff42d3a4278b61cd587bfcba477fd9ab7f739d0244;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h984f0c05d7d0efbe3bfa6bbcf2a4eb8863a586e2173faa243239bf76ac7f4450;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9ba97a16199e516e3d8eb1d5e2991b32f716493be7751b658dec0993dc296cf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd0561c860306d6d8db9e5f2413d205734524c2f248eec2cc4c7f4fa11299dc5c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d1c9d57f85408a7e5b13517f6ef1c34775cbd6f74d7a33edbb8c69a49d138c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he85b50588498c0894a608f57b8340d9622b3630a763958c5255e0e399cb995a4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h457bcb283531907d695f0287aeea0621b0c252f2a6182fa7aa76bd0865f2949a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h68e81e9103ac7004b9d8defbfae2abf289d4a62161a93a188effa0ce998ad9b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab02234dc1699e7b0dcee613e0904883135e1beb7116d27af846421595422d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9e92f0e9384a247e895ee5f8212664b4a99e168a2ac10468260094c92126b707;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd4aaa2431562521366de112c793d5e0c62c0dcc9b5dd3cedfb34b3f8ddfad672;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f782266b2d3779950860e327fcfce9f71d961b3c69f9cf3f140934011e9849b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdeaed1b09c7c962fa31418b9aa2c535b5a409d87c47c28f7d845f51038d8d5ff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6584c77b142caed46505c3954e25c6a4322ff0417d61dc37a34ea80a85c3479a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h211ff98022a82ec20997c2e725bce831a1f83247478bcc9bde72b7dcbe28fe30;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a954f0306c906b86e656eabcaa197aae054b1f3da0639695b6785773e4c55c0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hddaae9bbc7433214eead15892b35e902d4102cde52ea75bf72a3642c0a632ec9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b5f017660306be7cb88c33c98a226432f91e3b22f677e1011c5949dd76c4d5e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6cbb312f0b7e016e16d8e93b3f2e883b43924013f336d07e79d99610ee719f73;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha8cb0cb001b4bd346690cc292d72298e62fe82a6e1e823e3da169804e474fdcc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36658a459108e89fddec13ef85102faa2fe33a750dd78479dd38e402d825312e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h286930b643f9855fccbff95062930b0f57d066a75faea748aac94dfcec44c34c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8961276ad5701785f5bf14216d492899a881073fa3cf26b0983b0cecf54b1a53;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h95db6dd532e367dd867549a6ba7f72c1cd3d3644ccbddeefd777d1833743f322;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74135a79d2ac9c4483912dbb74ce0afc2aef4a347475b246d399dea02b944e82;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8e46e71e1e1ba6937b831e76e35b79297d96a6c2e4f1353e51cf58832e0c0bed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h499bf0b784b83315392bf1d38a76b70deb74b2c3a9cea05c3071906d63e432d8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h70ae8d986ca139107ebe1605728f2db5aaaf11a45b13daf5b3ffeed79354cd0f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb060357156476015639184d6cb4cdfd5289ce7cb64b8f09dc0110a8d04a362bb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd02f5254163f2bf7690a12927959b3a2ce5af729d8d71bdd1381a3e0b4d1b7ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9c5eb4eb33fdd488594bc81a0d15de358ba78110934630d8ab6cb23037dfe1df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h91c01c303b5b752a0a4627ce0d367637a36741336f316d8cb83cfa79f85690f8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3040f218130df25bd12ad7a8812e35cdb9210aceaad0bcdd09408fddbc82a4a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h43161a0a375a082a2f81b7edf40daab944c753f2e48f0a6579acbd3b27c2ffd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf139782196da44705995e1d24a44e2cb161af4a792fee9847ae71766fbcf04f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h92eb67c487c633761c7c49969d2631bac8dd34dac6e142f39054d26283756c99;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h61e4d8e2799cd30d3f502b5b5b697b7595b4ee9f6533976ba9b43da0ffd9e4d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb531b46734a00771a5c255445bbf42100fa89163cd20593cefe559a205fe5433;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h889cb542d5cc975ab0cefb476d7c90baee45e12b3ea42a3575928563d3798d5d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5741519574adcb6b1775fe309b089d61cdb3462e329626e48ee9ffe3cf619218;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haa0c58f58236d38267bd9e1b25ac5d8d47098f9d07b361b37b189ba7c7c73877;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5acb30a3afb94f540b97849cb751db1ffdd2b18c1298d055e4483c7514b8593b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h811ae200d4227d44e901d104f3b28d16ba38f7fa197123e9315f389f5fe4db30;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h311bec913e569e515616584803f8ca748dc38e6a2107dde06699b8e2c2ba3ef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h66dfd277ebbec2b031da5b9a482d94fe266a1418771020f879f2a07f6a48be5f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd83c688f726f111bf3f654c495a67695d820805c90bf81cc0274aa9d30470bcb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf650c0ed342895cc59474b5934ad44863ccf2a33cfd3a01b46c82aeeedede598;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb5700dc626706e80782b4fbff3ebab784b0f68ffe9deae1868731f00ec5fc61;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha0175aa60f3908ed38228bdbab1eb778b140662ffe3448c7e7fc8497b17ad67f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h88e2a28954d00fdff926fad3992c44a0db68e2b6f12118b40c4596317c32eab3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4900d77fd6fdf68718ac63c3417fc1c676605484ef901358024187030098c7de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72bdecf071027e140b2d19633b3077bd489bddb2ec8d42b526274f127b716d86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd4ca15b036d1f9aac694f96bcec773c4a20fdfa3e7457b8a4a754f62821e5b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h566906366a46f7a565276e0142f8ad3bb4312cd1e19f1a1e573c1d613c38ee9f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h324f2526bd7ffdeb08984c3079599c67013ff89769cec95bd87ba4d80235cc96;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf9d3206bc6a17fafd35c091fc3e57c8af8d1d89c72392c55a0fa20cf47082e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h106a75ab20ec2494d102259b7a38e895ba410e4a4aa441a13599789870e1f00c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h101b9d8c5134a3756429a953be84f47958c91e630c30582cf067205272898dbf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3fedd00d2be59e4d8ed301d7ae709a68e6a10e5bf17ada241952e4c89d1def36;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e4d3a1fccc9b0c83a5e01fbb04bca1cab74b971c3be6db5a272f46e3b0161d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd0b90795b3135c2b319c987a296e7f7f39f50ddb167e557131528c9e6a68363c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e58244bc28609c3ae32b75c81781cbf1fd855364f0935ba22e366c7a18a8b3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc1cece3afaaa919b4b75995276588c568e1d9e439c0f574800830ded965f6047;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h69d2bbd97c21125182cc7591f5c74208fa00a2bd7fb2d4dd351e69750418b7d5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h86ab46b993ea3b4a03a40929c8bd2a6027f7e02dfc89488ef87bbfda6a07025;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc9c5bb7f8bccfbb7e539da2e717dbe439f9c80214ecaf0bdfe0db9a75c3d686f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha9164add8d25a9cf817c2e744602dea993896401d09d20bfd9fd449c844fec6a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd85123474ed256966e04c27cf780da54d3856bff455c7e1529d155f874026713;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h16f6c887b0ffc1e8162814a0050c1588582d9481e8875f7448fd2f82023a2159;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b04330353592aa2f7c6bf8aa5ec8c4c272bc097dd646e003143bbd55f3f3113;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haae10dabab413b235a6c0907e5d1b2bc41924b61581e303e26a1fbd38001e4df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he4d97e5da3670a3a4fed37c7a2363b068625e8af6b22d0288caf0f5b11ba3f93;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4cd0f6a96432b10b422e0739998391ea78082436f35490bf1b342829a0c79943;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h73fbb539f9c61923e42cd7931ba224a0260373e5a01988e1fa51fdfe945b22a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h38e63f9f81897d46e0539234346d33b29b8f393616868eefa8ef9e3db846191e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4fc6fb74adafb25de172fde967e1bc9e72cb9abbcfb72dd0068b858c51822e34;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc6ed5936f47efc17fdb1db88b7b2a8e9f95323dfbd12d1ace4a850a255927031;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8fb5b7a91889ecbd3c6d8cb980db3b4e58eee38cff330660fd2e4501822d457b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d2450273f0d2b434b1695b2e0f3eb54e853d89129e0dbc9678c9205cfc6c6c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h49d2c1ed8ee42b36f5c1a39b7eebb5851b285b43703f095ddf6b1028af7ac0be;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h882787712f73be5bb8f030312e95a3b4a2ddb2b011f68dff8848c745fff33a8d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9cb94e9290537124e998bc42da903a3459662c2028fe1f96fa650cfeefc31396;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h43aeec9d2ec091b1cc1e0f12cb45d2b842605be4a88a4d747a8ae6eae65f88f6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62e332b71226dcca95ebf6fef0ce6aa07232f5626a2d40b645f5df1882ac1c88;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5d52ff8084f4b4b4c23175fffb58fcedd28c508e038068ff326c5f368787ebe2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6ac5e62195ad99e1b92ecd63422abe6e9ff5c87ff5647f8ab973c65f32f89cc9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac006615c29f9058b867f4ab7cc45b2db78410270132bd6160f83c98b7196906;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd136e17e945d56e880fddab516f00f846fca1e175e549765f194554d9fc3084f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1951ca5642cdf57ec4de1107c53d3f54cc7c963bb901e96e1e2b65e41443e3ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h725288e7b286b9e5593a2b73c0be4a5af789442ac1b9896ef301a1eff43bd0f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd2059e969974fb4dcc75469f0eaf8f7c414c1c2e25b3ed063aee34f449c601bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37a023469189e94b4ae472164086768db533a5190f0e35073ecd59b8f1371747;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h789fe55ef5460219226ff7c4fa5683bdf15d9de1b1a1b8ad7957817c2dd062d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4edce18cdd5c9d1720da39584b18f57448af17c5be0d07e15119dacd0bceaab3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h365f1d2b37a54b6826daac5e9b43ecde92a057255b6e43338f91637e16e5766b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h561ebaaec535a942cf443b48367f70ab4d7d1ef7e836ce4c9b84985341e8c491;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd8fdb3d12c855eeea6c8c814fd54dfe01705b4411a60a5050b114cce053ba68;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h21cf2664fd6780446832ae481d27e04bb87d5071293cbbd251a8ebd36f66a443;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd83794b07071869b612c47febd9384691b5471c9a8f6216882b98183849247e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1d004fcdf18da8a9f6979ec886f7bdff269a31d31c60e79e36917442cd2625f4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h204ee0429a82fe37d4ddf69aa7159bc9f35ec477a6ddeaa7f96198ec947cece4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb78919155476e165cb6bb05bc191f8e2c47607c32a43b4ef5a3ac0b0373d725;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4502a5691c4af6677ef047a2f43da72dee03355389e099e34f420089c679c73d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2e5acf9f69cb3400a6307674b7c98303937a5fbc1c5e9c8e82e47944d24d6698;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdfca55d04349f644ca2db3173a48ef433dd6ad821dd9b4e540bc60efecc383e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf1efe4feeed6438897728aad5abe9722ee16ae66997184bc190dd3394ea5222;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf1fbc9bb99d83dabbf41fca449ccd8e1bf475f3f9f569c6d916e4f4a7a9edfdb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d4cc19d65cd5840bdf973cc7bccae10315deeab3bade4cea48aa0edd16d1d34;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h81b4c402273a5984456dfd233030684872bff8698b17e25578fe9825ec09047a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h35c84216ab3ffd7cdaa742310fb1370e5d33f6a812e5a6229f707d177662cc9e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc7dfc3c444e5c0b0b20093fea200c5ef5c82f94c092313ec1bb765286ddbda9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ea1101592edf572025507e12e1459c88e021a6ec5a03a382b7e168c2f1ca404;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h786b31d54e16a058f8972fa81e881450506c9fd163a220cf536e1cc3465ccdfa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb69c56916ebc551a5d7c5b6bd92861955122dd18d10c43bcb496492414c3fe09;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1cd54ec55ce1068fb7fc0ac8dec78c5fe391ec64ae4e5241f12eee95ff432a2f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3fe04b097af482ae9194131a6b6ad021dd66b1613a860f97dff1a6681d479319;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h73fec33f8f8ba015b98b0d5777d145c2d28702b870605dc21dcead0c9614daf9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he42c6738d75f25c6a3c49fa63e62bc6b7e7e729ef61bfc5882b23722f2954762;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b5ea5c70daddb2d77b26220361f6d88fc9894c4dc2acfbf285dde3a2cebcf8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5a3a410cc50ccc7d7a8532422022f3e2311230548644cd3f4772e5026cf669a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he401c40eb21ae8b88b799c57c914a1245b8034852df6537fff9b0791cf428333;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haacd4abb8d51e5f1b48aa3a5fec7aafce37559c59959b0790a807e23524ffffd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hec83385b355e329d1413991962ac65c938fce1dee5d37f7514792e3d10cf089d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc61bb94db9dd7dcface5ef0ca8791ff14f5c1d042d4e27397a916a94199d1654;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb37a401bb098137786629a258fd7911360dff723e5914267eee4fa43c458c3f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2141e2ac1bfa98c025418105586b8f2dbb6545f60ac8895dc7957cd6bdc03e68;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha417abde46e9af9dc0f3ebf603e6848b659a90828826658fa85f4e5dd38ce351;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h844ff959687787d2731bfba8b0df0230a4d77ff84786aef8c7b0ff23e12bba74;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab0e62b46dda6c45579e78dad6a8e29d33a06f0079be50625e7b07785d9e398c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c4ea2e2e9e638c3b621721d3d2565cfd531f20a450fe74883124ff21c46fc18;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2ffab040d9848c3559b8dd83e2ac5d87df8964df0697b0515a7766c5f99dc5b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h10ef78293a568e435e5ca6b27e5bd63651570a5ab1d0b89787f322aaae8f4c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h575b5ba8c9b044dc467f6fe7917491357cd84a8c4ac35e436763860eca610191;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb70edcd49edea0d8e80252ba1c5123395d4ddc5505c97ce216a37295d418a7f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6fe41e234764e9996c4a63b53562d9442236113652f59d2644744e8f8f546318;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb1ebd40ae2f54986c41fe7d8749439c3e6229540d9ada336508a0e0c70005e6f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdcc99688ac0c0c639b70bf437c1e9fac5c030ad2c984dcf2022eca75eaef4507;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb45965fcc1f12241816f76b316c4ad64919b062684ea245b0b421bfebdad5193;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3126859211c9bde193d7571995c79542b5627c52d448a8e67041d23a128e9b13;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1fc2f276505cfc65fd126cca4bb4d4770ddc10fa86e8a5945c48089759e522eb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h55809b8ebd5d5d2c6df03b8c64da4fa033668532fe8e653da0b760f0410346f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h63608577a53b3ee5329107b3b8dbb4582608e0a9107c12a4d5508f4a658b40b2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7aaa0fc0ed552486ab56ed128b89eb5c9d8578c2678d375237363996f1341e12;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd539466f200a0115bb9adb316d9f44c5e404c0c1c89cacd22daaa1afc3d615f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h564baf39b8c210b9c60231767c1241387714ab488fd806952a77a8e723f65121;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h88302f741651f2f9662e844ca3152ffd5094c4f686126ec3fcdd50d43191945d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9429733e9d63c8962f1cd5bda32d3246764885ff0dd9b28f8673b221c898fee0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1e219ef1db3a52f8841bdec8a46326bb25b1133f608d701455dad55e20803fbe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee546ca91c92395346883b27dc24dde2a2c008e2d4ed4f606ddda018503c14df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7e092a9f27e7f1801903aeb6e73ff4838a9a7a46679fc774ab48216f529dfe5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b7faa3b6d25920d6ab4da11067d4dc41d54cba910be82b418bd8edbcde841c9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3221a36035f1880090b4e4be0a95cfd4e843a09236884e24b32636def4168943;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9af174ece5b30ffd6842289a270eeb1b213b6c1f07554c45a5ae878182d9a4f9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1567e08739afdf03551bad533c6c476100a7b4cd5739645bc562bba1541ab90d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3348515516a565eada48e411f817e3d7bc7e5e3bf3209a12a54ffac55d653e85;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3ab3d4319c459a71b214a79f2481419f3ecc2977ccdf46c9f2944c5f9776afdf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e1f1cb2051966ea89a2931669da727eb131cbc2c59a4ba1511d4a79bd0bda13;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcc612c449ece60c6f4722ce315dc7358fb62da011e05f82b4800ba9960a69d14;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b8ee8dabf335648cba922761e611a7bacecfc2df599ef1167ea6f1f79c101e4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6bbc0a87be209147afc42ff68252d8b6a5499755e955d7f0df4ead10aecaaa34;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6cb4036f0b8094503b647649df456a339ea4ad23061b2b934e93dd85c4d8a9a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf7d963a2c048964922476e79f335ce1d8e08d40079a6f7e0e47adedd009c8ef0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4e989b3620f5cf961602f48e0fd31265f0ddc32f3bf5ae5ec420b3323dd88110;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h86b631b86428d04dcdd49427817824556ec3950e32c63996547e670b55b95ec5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hef4f50d3b27d7614aee628994c4873a559679c9852147f93c62dcea78d450671;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he13b31e8d9955a29d99c755f043c65885cf733dfc596e16fa0fee5fa06f9ed3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb385088d9ea82c7cec038471cfc1ea4de0573d59cf8caf649d91717a3f6918fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc6f4c340bd044ccd4b91c96911a44452d88a476dce903559ac6ab2a69586f128;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd89247b5cc98770029752a24b24005bfc16ffd09d854aeb2480ea6c0689dde2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8b8171d4df245fcf24a75ca1c180ab54ba2cb330e90ee1912cb7c62f910d3433;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4400bcfd98146ea0a44e4c9fc5bbcfde9f937b69d7f191b4ede90882ea42142e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc37a7e7a795d076e5afc9184fcfe1c43506b02782cbe52034c6186a5b8e12e80;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8cf76588e93e6e70c738772cd4acec4f872fe5b06f87badab6c7a7b766e7b223;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heeafbddd9296fee526e5e0ffe6aae8c56ba00a4f457af74824e7ba22e3b16721;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd654198beeb529bf21b6927d4778a715ae317d02077d59711b639fd3f6a4594;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb400b289ec4c2f9b3236e9cc25176843a72633380098dbc15a344376ee95ca5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc5c91b89dd92158b66675013f12b2b95b318b7052d458ffe276f564b135a4922;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h86a3444a7100c512583294da2be1ca95e2ce1f531872eb984aceb923ce03ca90;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf10a4ee25f803be58b284a78e661e71f1052a3277c4f1c3fe1f1ed60d22715f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d3680b8023c941dabd3f6d0807092180f8656708b1b5be270cc918507fa4fbe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd4042f22eec35b5dddd195e2f849e48c3b2f69bd6b730afea90938268cca6d70;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc83a2018c2eedfc2bd9bae543400d34d241f2c86e16d52462d5f59eabd972588;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5429313988be8b92254bf9fe1570cb030087361c9266b21ea7ac31e201b288b6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9910bc1995f0bccd3e87eb16a753ea619fe63f597b1f048f9faad6c2af72f558;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b339d157de7ccfe3efd86871dda02ceef245f29cb07b7ed1a1014fe5dd9bd3e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36a1865a6f5b3d10c165169a96ac5fb9f78f61e69c7168f431433090585c0555;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd5342a614c1977debd51b701342513a8da205a4f3cfeef575ddab223ffc4afe4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfcb4168f0da87255fbd60eb7c60a99f1fe1eb150790424ba774d5cf3f70c1317;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93298821811fa79631be3b3c65de3977fb895a4e5f9d2b6cbb308a6ba5c32de4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h229c9569d98b5d6b2f47b270bbcf6d2362d6969108030a75a0d5fcf3079f5f1c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h142b43b00a7cbd9f154dd76d70d2a3e37fda5b651b876a837a8e9d79e6902e18;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37a4c54a9744c91492c412dce26e0a8421f2145f265c2d939da0ce014d93c1b8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he935b2e6372215a68b13efbb8e50b4a17c77f06fa2f29fe588d3fc29960ded3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h26eecd5509a4af0cc2c5e34bbde796cad79c4d3b5347bc454f52e5f1c3d594d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h87051f076e739770565afb748aa0824d8d996c74a07ccf956a657a22d644e6cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h96d9c024290586a63f771c24dbbbeb261ec1256753a06e4659b3b50965f53edc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc4685ea550164695e6458f381b61ad3797d5184ec65b01210e0705aedc453d1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h200e4d442c333c71feda69e70d439ba82d4f9762d778a818bfc6b495d0edb3d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36a91216b70606873220a536944ce3ad4ea2b717c3310535e31741ae0327228e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac6f369925b10eff1b056455c97c814311176cf7939aafde402e220db14dfce3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h49a1b33aedff3c1f0d78d41510dbe9863ea6e761f843f0b6f16050722f0181d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h66971ec03dfb69af39f2550a0abdf94be870ae5652392ec419430ef37114086c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33014e6ba2793b22af5041eba94e393c5cf5834f362ef7fc855ee88a836e5d5b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6ffce97aff9a8ba00f6453b1968e96df555a0e089f04f528795c243d554dbeba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9d24df9df933c8174802948f7377e99ca4d6b9d7773e45895e51fa031352124c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5939b21f122d10fc7023f17de6dd7a179985f402241b9fdf9e6bd2f8d8751a4b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e5f1601e0251cee20ebd2b9737fcf6f09e039eaf6a022d2d7a220481e7ab7b0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb6ea3116aee5c25f8a9017306c2a876c432881546e859c970fd3f323cc783307;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h84a9438b1a0fe1f6da16552782e10a8711e41983e0ca88b3ef7e26225e1103d8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a7441fc8978bdaf596c81848210557d3aeb62b6fd387315db482e39a2ce3fdf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2acaaac67061822654bd1ef3216b2eff2470aea0affbda297d7e17c39f35e263;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6c32918339f2ee9d51a41d49cf6f36725102ee58df9169b4d3cf8f3bd7ba0f90;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbf0aa2efc9c0ac54be8ad55872afc60725f83eb14b01586072841fba80ce02cc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h71c2696530f49c4ecb4c6db9ad0ced2c0247991f1414ab8ac4433df402d6b7bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf9084a2523c74a76d06de2fc8ccf6e8d451d4ab6b9233ff0cd387ac70f912dcc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9dd52b5a1153a0fc91f3e1b9e75c41086f6834464019cff74e06346cd7703e79;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h49b2c226bcdaa751acbe20213ba259ff692b9d3ae7e9fea2e6ec08677b482e18;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h694784bed7a19f064ea88db68ce1312fc8ca1732068a12c151148c7e5f6b2a5a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb1181db7ec1887fa29de591be875ab366ed2667db748c46bfd2ebe11f76b3e46;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b8adf60d511da321f9e54022cf1f0712caf4d45ce45808782e1d5978d9f3f54;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcebcd5684b2d3c6bba3310ab0ba2e3e6ac775972d0af6d9cfb959cec2d7afa6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h129c7cf6253bb4cc4e289df8e380279b1a0f467b143cee8bc40a3a3cb945d7b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd4d7b433b8f574de9a06bb9bde059c845cc80243c3c1700ed6c0979b834dff3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33799c07e3745f10374374d5762ba02edb360b1c5154cebd286a982f863a0766;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h53c0669f781d3397d9ef2589596c8f257c4a742ecfc47a52524972f729bce532;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h91bb253fb65348a03b54e74814295d402ee23d4d4bcc66f1de07c2c803962cb1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcbce5d9884afab32a305df079304ab20972d0d33dce239f3dffa772f2f5abcc3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h91e63616cc796bf2aebfcebf22bc3dc394f0bce5bec1e874f4c24f20c41f3175;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8d23bd3b30e8b153ad47bc23135059b3aa0fc1dc43f29c9d1af078d49a995465;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf55c9ccaa588626364182ee6078dcec5d72b14392462fbccdda218b5f7365971;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4594cd1318682e522a6d6da0c4f584d424537e1d3a7bac8a70f6e1db704fabb0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2bfe5ed7c63e6e215169ac19b12296a6ecfd4beed3f95760b82c20dbe0bd4b66;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h91f9d42d1c0d1ea0efc1c7a3eab41ae900f77d02407f02dd5293a39ea77f39b6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h40cae5be95785afdbc385d9d90fcecc3f0293d6a096b2faeb10a0e2793f25dc1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6f8e1d2af1cc0ae69535003e258dbc17f795e5b534a07df7f5e292d185e5931f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h88090713e778f1e17dc3e3e0be14f6e582ecf13ca74a4dc28c97297166aabefd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h35c36b59437c468cbde5bc5b95d876254791f046ec8b93749f9fbac473538b09;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h54f2875766564e8fede79ab57a33281f4233d5696a00292d6ad9761dcde811ad;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b796d0074b4ff5aca36bd419a98a524c5e22217c9571a6e8e37305e81cfd177;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcb5160c3ebc27c0c9957df4af9f08fcc06ed0b8c628bf9b8225f65ae81aaf611;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3e2e681735d31f48d122e1c91845f212df67bdb68dd50fa89ce02f875f767e11;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haa4bf3c8df5fcba0eea08792fdc97ceaffd5dd41e0ea56ff85829326b4742b1d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h13b8b64be2e854b9c34d35f55db20629fd2dbc9ec749dee089e52ee34c0f3f9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbbc1054953cb60918cfbb0dee82f3d80492415cad296d2a588c0ca53204cb481;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdaae8dc606f5960a56d078b6296d347e99ec97201a969f6ca994bb32bf9a2404;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74338da15a053a7da590f6a2b77fcbc66bf164d9ea81cce81fda8a84fbd4ee86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h20e41c7f2e17a7b16b5f1edad1b3e14ae8698d1216ddabfe2705644f45c398a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h73c74b28daca806189c67c9b909f03f3964abc93face8993fbd6589cf2d56561;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcab52422e18cac7514e00a1e7b027a7e8d799e526255124a24209ea5fae0aed;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h562bc4faf1603d8ac43fc69974f331e7c46880c8e053839029a01bcd4430f7a9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h10fd32fa1da96087be391fadfb2ecd4690d3f03a4affc5c7dbd733b4b2506142;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf1d04b749544a7e4d657aba9d527ff386c568daf530818f4d25f0138b6add062;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb39504be24ad32147951d59ca028af42f3a7bfdff3fd2181719a6cc9ea8aedee;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf5d93c2e51cc9ec89e6c2542c3b5feedfe9082f2a4fdd085bfb9f24c9304ba33;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e07f45b6ec8ea395b2982f50db270d8835025ca6cc251ec5525e9cd33767b42;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h634db9461aa8d60a2326605c43ee1fe03556fabd6175f70ce7742d7f265a0c53;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h98bdeef91e405e85ea2c249bfffc960f56c80833eedee881ec3b03240cb328f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h19c65f4cf4a6a950b0fb9314b0629f76f8fd24a47c3586bdec5ed0ce0aee6f47;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h62779eb225b19a41161d285905fca839b6d5d8a121897cf849ecc1228c8e1dea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e16cbd2b7f9678278d601f9688a50f2384a6b096a7ec66bd0a2f07430161560;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb7b55ba7c4e512b3901443268e742d198ea1ffe0b0e8d74835ab10b4c4d07a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2d3e91a5b9b5174c210aaa8d3645c6ee3a9096414a84c3d73b74c411cf3aa3b9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7ed642c49edf5302e392b02f8a997c2bf2d7c57372984ccd3c807220b7c08007;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h88638aa4fde4d95b58c00f9e86c08d91e476c9d96920c227039d6c95370ad332;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h10da829d0c79b325b6a5e10be9967fffd7bdd8ef5b93c78b3c2a158c28914168;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f4234e68aacdcb416e37a23714e330b63d385af00a6e4dc26e8c4b344df1705;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hea89b31abe5c2ae513470788f7298b8d38f859a523b67600ea788b2489e49d2e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h78dbcd650bdd7eb1bdef215ceb59cc934af265cdf76dc2c198ed2c65fefae41c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2b03e2287ed673da6aa04cbeda9cfc466f7266a722c4cbd4d8b63e66a419bd06;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h25822be6049009ca9a21efaf2e7e0d2933c46792fad7833d3e0954d80c34418e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h585ca1df3f03572648ff3e135a72f88ed15bf2cecf2270552a145edf42333f91;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h297d2de7f7bef0e8891546a5ba4729e82c130046f2720bead8efe7d9a1672f3e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4fb73f4e5324c7a066dad3aca505fc5264168d787d64bca2c2b4f72b441396a6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he1aabc7087891536a5961e9fe3108cdbbc2ddb4663e260fe9d5535cd2818a4e3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h778c25a0091ecdfd5571f36da83f6624f264f0d480da0b0f91bef8787b3ac6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb4aa2f520c6bafaa506d656ebc2e64020f2801714fc426790143c30ad5fec2a5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc34db3b77e5c0b40de2efc0f7eb8ca881003e68f2e73d6ec64de18e0b90266d4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a61f58da1f214f739153faa71c821febbf5a155f852e99d3f2ac0c5a2799f8b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf0b5f6a6b8346389c222f9f79952aca0e19d817421a41d980f7d2772099c5d68;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5ebde98e911b9edd2c15f6960ed870bc5c60474a2089e37d825affe053d63a53;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h297e8afbbf7a5e9c78038e92132a61a83c1c1a148f3fea37099b37e42927bfd3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h59463f88346b619c362f73ae6673e45f2467b13ced6b14a2aeb2198c601eba08;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8a57c97ff21cde03de68f9b1f5dc4679c3a96a25b4c6d0dcae563ec347087abc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd3adf28b6caa9617edc81ef4a33fce2bab45aabfaa336c9507022c589ec516c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5324b4cfb0e4cf6878f7bfca770a403f756e3d518bf38a83ffd5eebebb509045;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd2c29eb8c283925afa61a3639d29f2a0b9fb2b45d77a7724b97f5176045749df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1b99c6db3bea99f73b91f3cfbd3ea5cb0441b676598a45ad3b4b28b2e6981e57;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf742a9730e41c7aac04f526c80dc08ec04ae292bd3d299cacc621a5153d404b6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haad0555175ab6c6e96d5e6c5f9d35338516539753d87211668c56adaf8d6c4c2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h31364bc181ac5487d8df9164e7727c0b9f317de2647d748f0d4c773e7bbfb832;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hddf1378797502b36a0bd99dbdb782637ca4a37f39422990497279768f4b2bbc7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h933d8af3f122af4afc893faa68750c4633d4534bc3b71a8ca4b6010b437d853f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd6c32e3305e524e1324e82cdbf7da133ade0a2f2d42afc30b7aba6e64596c3a8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5b3d157063711867b14cc15ce90df729a3f01759b624a1022ba7f845f9bb3da7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h39d4d502c66630b8dc3e4c15e18cd85e61d03d48374bac1a7b54d08425c555e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd81f9f68457074471e3b1ff08cf2b864c103860c8cf37f3b581cf6fd0fd1da4f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he1b8ead1c3f9401465ff816263f6dee040a62120537f740b344e013153b6679c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc8f465de9cb2fc08cc6f086eabcfa5aa06061c259adb1d3a8a38d5a034ee47ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h56d6433144d58ad935a0ec43caade7578ca77267960877812a9d48269d3b385a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h536f15f67c9894466881b118339efff23d6e86e29cd4e651bf16c1d6d2df55ac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha3e0bc8aa8da671f4debe5e1f3a6cf49933e46a19f94100e4715d7a08010f31d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1fb3ff59ff9e572827ab07294a76e5b42185b685409bca100cc94dcf20588700;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb496de9b15418860a5891614373639e89fca29b9c2726e88de941550eed6113;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h73292cd2e0905382ff7d6294ccb94a9e88e23b500a1d8f5753d7ddb4ee0188b2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haa7f2113f4f7cff068aefc106a92aff150885d1daaab29f234d5ed8ab683aaea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89826b6cba48ca92707da99b3ff392ef7fa67b43233228590d2b219448b99e4a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f06e844215c5da00054308f467954c52f7ff0748841ed2076aa88b81ecb3589;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4c6be6b004ab65033931109310c2e2622e68212ecb05851baa4aa3085199a739;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4702383cb6bb1010f4d633d87e36def549feab1c819486854608f05cc3199059;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha15088309ac206f683d68f79e9052f511cbad0db27d0069f798c29cb26695fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h171cac5b60d13962eda648fddb5d13ce0dfdba48cd8dd0233bcdcca8d3031c9b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7291d8d2793a9715223079f26492d621e9dd8ade489f35107b5864bb01225ff0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h80938a6e8a90137a31aba40932d16d3016824816f0417ed0c1778d113a7a9e31;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf43bbfb5dbbfc692efd35237a28d8d3d90d2775be4e4c40e34ca41ed26d4ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h56d406f6012f20d8557903fb9686ea14967829fc14627b155cc26ccccb1a423;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h455cefd80252ca09d2fe24869309658a9ffab0b468d55f893377a3aed71bbd42;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc3cdae64788e70dcd7f92966e87fb1acf80f103821d3ed9632e18c5592d5c94;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hae42f1656d4f891dda0e541780150f99b591fa7d837c05c3eddc2ec8b4c6364e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf6daca3fd4b6588328eb14be9d1d9e8558be1f99bc6afa10dd1cf0f15cf033c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ff8f01e39893e77e4d189b2bdbf54a7672fd7e3180f7865dc790a10005447a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h48318989bcd4bf27275c7506fcb3ed3d2fb853aa79e005a7772ecc14a36724fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9212c85222e393e7a9e708f399bfbc061ea2f44cef7526cb21d8677680476984;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee52447f00a06609ffc15aa26532efc90cc66b2e761c7157ff371daf1cd3a2f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h623f948b82bed78d3c6bd0b00f23bba1cf893e34de69d0fa5e3dd09f3e5943be;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha50dc26e10c042bdd31e24d1ed973c392f271828704d66516739b903d8ac1675;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4245b31b12b6972a00ac43e8214c61bc6c868b87611483c5d2d5cc46ce740883;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h21179c34a98b971d9ecef73e6e6c9acdd6715e202c5d16feacb8cdb41d8aeaf1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc3729c6b25de71a93a45c19c0de5c90d22438aded9b8711a175e21208f7c521f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb46bde99a338828be32986bab70a565dbdf63dbafc4e8c1df19cd84a7ef3ee8a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha87294736f08e52171d793ca21cf771ae4771afc3ad43b81930fbaf6db26463;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1741214c73d17ddd64c095cfe547608eed4337b1c8c09a7e1a3f4ecf0bdb0076;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc5dc45334d7c4f19e8dd9749e6417cddf9044767ca74009453cbd49c81651dcb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd9eeefc251aae1b5ede58e75b5aabcdcf497591e605ce35e61f141b16ec2a57;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33df7e731da7e741dd0a1d1843121d1f1136495c54b011c5d61df32f73498fd3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h73d891f54e60470ef5b3307770827780ec7044236ed90df879fc5ec485a2013f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7e35c51be7a33346f9428951de50748733014c33cbe9d11cdf9ded85586ed9f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5e44c589defc5b9fd7fc708cc48ad8ac00f4a5ef1bd9f70cee35ad62b2bfa5e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he45bfce1a804d692dbe7ed0576f8c8708dac690e2c25c08eff8e156dc616dd2b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a352f26650adbd81ec320446b69c29120996a52a564fb6a71e223008129456e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h16cfca82126b4ca7a830f82889e1e8210dbea6b7807d0592dcc36f1f2c9d514c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'had580cb0a1a4563cbe3ffaf84bfa84e4ba2b9bf3cb2d7841ff5dcaed1d57066c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc44f97d6f6234203073c91d4ec47c933f7e7d55b5330c3d6efe0837f43334ddf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb1d8fb35ef95c1fc85583336603cbde05fbd28527aa1ea9a7340eee3005764dd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h526693211728f79aecfb2b764b4372f98c46fa6026554a52ecdd929a2358eeef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb423358bb3e5bf1fa1d86054e9d7f3948577dde222fb5926e0749ee38eb60433;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4882b36784a59de5ee3d8d54c5398cbed3ca8e05e83bf106a7dbc8a62433b186;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbda291abb512fe480dd54c4d5d28f7df7abee51ea021877acb6b0096364c5105;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h78f43cdb35ac005c38efd7ca73bff51fc79c30876363ee6ef6387fa01663a15;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h184ca28a83d4ecc9a925dc511aca460fa73cc3a14966d7c45c04456008b62326;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3f8b5924a77ba91e3fcf7a5db3024987afddb16eded73904823498cb793c8558;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7563d587840b0254fcda43162409c8557c5dcbfd0dad23b64851e9e5153e108f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2f6c016aef64494a880ed8ff419406f6d95648ffdc9de45ef3ec069970581db2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h402b3a2d0352f03cc2d00fc73261b597cc5d17b645885d1f178c4e09724613f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41c3c648ec64951e9b4e62bee0f0c0717495fd25ea32329a82e3ede8d0a4103f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h634ce3425523c60e22b20375f50e07f8d8041f4b24f2e423aeeb5315caf5f546;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd44dd8ed7add85f83d52bf7dbea4c803fd4147e864b652587d1ca527ffc1188;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcc17e9a77e1a75deb6f77a597aa18af19c63e4dd7437570e1479c6a11ff2e7ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd70298675596acf7de3f43d1fd6dbf61f51e0e4f4feb93b152d6ec5e07fc4bb7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h314e55bfc791f169519b32a6aac0f6f56e36b10f36f4a3cf66fd122d619197a8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf4b5fc773f5a0cb3d515b3666fa0f6299d860848ddd8d636135d1e6772a47d36;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd8d2182c246c98ece34b04b02dedc23622752ce2bdc48715704e10b0a2ffbc83;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha35e8304a2fb878ba20aa040a4c9c368dfe06f590bf61939896eafa149925e47;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h240805fd1a2867aa7d43c60442a9240083c4751da407945b54de6c83ce403a72;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36667538cf2b838329d5e0b52f15f3c31695f2c40a1aa4acfa8b497c606e8587;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc3603292462f5c6e802861d4c066d8805900112fdb8dd9f9634ed4e9a9e92479;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8acce3c8a7e90496c99a31dde230c518d6902f3fd5002ebb2a2f0cfbee806491;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha35d45fc7edb0efc2471ed4fac08815f5bb01aca180713738b0930b5b5b22677;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2bfabdc811df8d72ffeb8a10de2c9bdbe17c44548aa121f7b7b191091eaab9bf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h905ecf2e11164fe8c12815bc2645bf5ed77f1956b99a6b98b2af3fadde11092f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb58b7f10ec537c101ebbd72b824fa37d054859478ce626cc4704c72ea16a58e5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbbdbc7b3ecc20356456b68b18a5d12b39609aef4884053ef7b63b4b0062698a8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2fbaac5b295889ef7b63ae36f70e3406dae333ff57db425b8f955b19b584ebe5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc86530a9c4690537a7db37caa9cd61f1eca4f1cbbf4026dbd94a8e34935c7cd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he82b45a416b10fbb695132cf72ad9beea971092f23f93d54f0a249066784577d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c94a4e0d3fc645078cb05bb97a651d6693dd4ffb33b026e3908878af1ef8a4e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e803dcf065a07ee3c9e959e7977fd8f3ba8029a3288df14af966b48720f8635;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h57f685c2ababa934d97a0f473d37877ec271b513374365711381da9089071dc3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a8e493bb4600697c548afc76e01722352f97dce1ef8f946b979267d89bd0cc3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha026dea8f19a1c830397e5605257da730b41893c00f816dea58c440d154f3120;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf47a583ba0d41d07a61712488d39d2527d0ee17047776c97601cf313a8a7ffc3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he7e2150779b80958dd9aff4c628b4fab4ea8c9ba72de5cf8a0e4efd947749c5f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce14ac8f1538d5a6afb98fae4288c5f12deed4dd4237ea18e67623c49fb53f07;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h93c2222e6ad27b7fcf7279c26b1856156d393ec7b66cb52c56b0f966f0e20ef7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17ba48cf58e9deb5a395d44afe399a6de1c2acbb465a0250c0bda4c142740bfb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b5ba843a2504c033db8b7c0b3bdd4bd535b21f82e22c983dab3fd93ea4f14d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h561747d21042fc54739939d6dc330de3aa0afdd157967dd35a8ca926614c562d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he9f6242164813e26cc7fae03748908922210fdbed1bec4adcb3ab53c905ad9c4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72ea158abbc62ba54e51377dee76bca9b0ea4769f254dcc94d59a131a13037ab;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haca4e687cacdf575b6cc659c235f70f087daf2409ee5012197a321d15112abc2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28d2f62c141cac897ef9d734d80c2470d1b5a307d231e4bc4a545bead589e50c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he3927483a4f26bba9ace2a28b4215631fa874fd400a16b6f5d279d7f279e203e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce10b76ae35b940a0bf7b30bcbd5c96d138d68544a8513ed941c7e68f847b458;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h64cc7369305de45bec2b1a5230bbe7d2a7010352f8afceb351a4415c6ceaf988;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9774bc7872aed6ae6d2808b80cd931814c9ca126c01f4982480e8ebfa4dfa49e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha5087774a705a4df5c725d991c27dd0ee0575f2a598dcc4b999386af29e1efe2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h61027f5bb6e62a81090c764739ddcd16de2f6a24ac3222e44c4fdf01fd5c1091;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc8702b8d746b7bbc2fc75d8782affb1ece98f6531c4afcf67d782d4ba5d1df6d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdd785eaa76618166b15b9bc15825722193c209afa17674620d23206ce4bf26f2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4a6b670dd37f0d9068547c2fb37cee0697fed4d3a61274f856de9ac7dde02235;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcd03085cd31df65e57e4bcbc9f9b4a53017f8c6dd1c97109c0e1ba9dc03bbfe7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb51aa97a69abc4387d7062301be619a9a28b4c8d00585be69ce1e9958ae03b71;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h32b0ba059fd543221a92e1d50916e334e5b17b59ea6b519f72e2273dff55009f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf8af93278c83233148095052fc76fd9e774814d371c62f6cd9aedf46be8caf51;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72ed5c9262878ceec2ae22f83b86a816bbfe61d69e5f3c5a6937a74b2fc292d2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf2f1b1ea1fdfdc7749d534cedc6a1eebf690ca4b0cf92648db462b85ad3d11c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h494f683fafe09106dc8fbf8ee8924d549c53975b19cd13f234b00e4f9c01be8e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he406978b723e9a2b8fc4d5f27fe8511693deeb7f0d674d74cc098dfbba53a1d0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1078fe2b25959858bb3eabfe4561ffb19d431c48c451415b609c92a40a6bb260;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9b8cca356bc4fd40fbca0d7c2da96f549ba136be9a08a4b80f1088f512af6c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcf6cfce6da13d0a5c654342e2abb6f6ec5939f0dc95f4717b786d4bfa48be1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbcc234864a934fd3e9c58f4ce787b845bea05af64fa37e5c7b379a86645b3084;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf62f33b35b94955a99b7aba194f0a42cf2790c362fe792ffecd7583b6acb96a6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h65075e8f2f71c2a6049d06b976ceed768433e4ef93f9b30f66bf0f192099527b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h94113cac28fd6d99e2b62ae913888f8209c32239b509d6e7d6199ee1ea6b30e5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbd7e4f889603b0208c31f04202a025a6bdaeb87eac87ceb2e50459aa0356a644;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h55c0762c4430299f262d5be134aacec29c076467847ac4ffe81863624dfcbb09;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa7c7ca36dbcd204c5719152f521ba625056e9ef95a5a65bdf5c95612b33cf75;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3da171d92e8bdb80f4d89b856cb57454666aca7764819a88f967ddcacf10e6f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc6069a0e45d4a90ff503ce282df10156824d8665d6b55f8747d3e91e30967f6e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha955c4a33c9c81d5624aaae49f74b73fa842ea4bed728f4afe68ed4e01fb4be8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h25618513087153a3e1cac816e3d4abe1198eab93c87b4143e3d4e7a2aa3059be;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7fb1ef0a745ece1e35b0302a783ffaccbd2a2d965709d790382903a2c7740275;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf2c38408d682ea75d1bf9a329362d3ff0ce73ff1fa5b60d0e6f9699f19def0bf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd16b65e748c297c53ee78db4ed1281eeddd1e3cf30664111776bae4de8a4b918;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8131ca06c61f74c705e21425803521454aecca5a9c429fd3b7514526ede7adbb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h946535182bd4275e223d872724f7bb3cea771a68eef54d9648a8d55e1967840b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2dcf374e07d6e2bbc5a0fe85ac01e38f5c55ca98149da72824012dd98dd33795;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9802c500b052237e672d116cd3dd493ddbb65e6d7499125597827f3367c1f080;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2dfac1fdb0fb11b70f8bafcc043927699be6939f9b23f2ebcca02f0595c562df;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hce81e4ca3509cbab1eab7f0357de4f809ad21efb9b22c3cece6c8ea168676e13;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3bdd8783eab233be1e31f58945d9d99498b91673a7b1d1508ed9a23d3f42538d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h13053a9643f5c5b8687e1c925aaeb43fa6b299eb95ae5e320130a6041c8f6bd1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb89b617cc8937efae562e74adb7af04d2b3949f13a22692b78fd0d31b2a7be55;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he6cfb5d3a658f0d1e0c254a3c498f078b3775d49e5f66a4419c287dc567ce2f8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h97d23e07e44d018c2575a464781309dc4eeafbef7142ef6ce20aa4665ebcd344;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd83eaf79cc7d6b197a1ece6118b4ffdd00dd90edbba00fd0609686c9fd99fd30;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4306bc31101615174e28e9cd44504b10cafd451db4587b685003548e3e8ce55b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h24dc6c4b5fc20594f5aef94139f4dea19969fa96088efb97170b3790e23d4e76;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he8debb99d000c02b5dbc22a834a1c484e5763afb95afb4c19e37f53d753a270d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9fdc46d04967d24ccead65588c6c82aaa1486ad40ca4db94f4f35924b0e75f1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h810d3e5a8bced06ca5d3da3c3be10846c62fdcc05ae3bc8721c9a6f9882b5ede;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89989a6042c46f7c3b0cbd8eede0f853ed661afac1da433680ab6814f2a358f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4ca9824d32915febc23a4a380c5cf454d6faf79ed43d89b7fb2bdbc2f587651d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he5d42b6c76164a88ee3e74599a1e76fa062c33c123fbda5efebaaeb4c6b35d87;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83031314fb7e2e60b4b77d8be0357f9b5b1c23e0a0888c8d4f12b216204bd197;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h88fae356a116b1446f19f93fd310210e13e4261b2d878998d762067d5b373aa9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc1dee3510967535e02ddffeeb95b8237892e29c90e2f41c4db3fd8555c579b3c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7cf1469235a1a63a4c66ad0bf03175964c2695ae08b5ddba401436c307716d4a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f74cfd5278d11c60c107fac078e998c1d74997cb748369da2ab349c6de04249;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb21b8032a877101953e500de0876f7fc43da927fa82364b8473429275d03660c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haf50031d74a51046941b407f85250555eafc011ddc436256d896fe3ecbeebef;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4c8949a2aa6c933cbca5afc8e68ade4ae5b684525f36ada492aebe696f4e130a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha6d4349119378835b57876cfcbbacf1273a6537a59cee95af6ffb3e928ce40fd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h718840815a8d6ccaf2d1cfd9bd244b3b3a5c0da518918fce30f46c9131487318;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h22a683398218251d290afdf91b35c7bace28d59484652390bc15ea4b077e94e2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1017e223a15d95a7675a18037539a73b561de46f14e4899ba239a60476ea4032;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he99249df3d1f9cbdeffdcb9b88536f1d73ea242e6adacbcd89f85e85d3b6cb60;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd7c50675b9d0c9f7ce6b8bc63b3131df3f50a3a419664d94cb64628f19f1fc29;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hca6bdb75be54197419d7530ff6a0b8463ccbd032692b291425a150ebd15883a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5311cac9cd9260a1e1315d0638a3026c0b7ba4c1248f87e65d36e73ab2e074f7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd572112ee19dbb243c0d85626252f8a25e0be754ff36ce444627cd4fa035bdfe;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8876ec5beb87c132aa58e0328d596881f9cd8e41e7be43526e597b6e0dcad608;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3dde14bfb3d1c95809b65b72e5682ff8cfeabe0ab3a4ddba5344d582a0e2f67;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h295c597c404c5592a36315954125251936dc843cf21a4863c44ebb2eb844066;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h324162d0ca1ba2560e50665fb967432c88a7dbd111ec2346e6a9afbfc96b67fa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c7cd891ec27eb66202d84e23e3e906c93e4388407c355a247e08ab057fda236;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b3a090f5b4d7cc7ff53aa932143c0ef57b24dfaa12031195e4376d5a20c91c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2a0aaaaf5f415b3110a8c504c3a2ce97a05866a0ed795e0ced058dac9c347d24;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6bbfc8012ccff6bca5018c7319400932c92054950ca675073bfeb88ed036dde6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b3ba8c5f48bc2f3c2692cb913e8f65398422b1e245e13b47513b13dfcc78c07;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h568b807a4083dde97a52e9f25c0f8e2bae046e714a05c6c986253facc6037273;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h182f5c86b43979ee22898e0367df5c3dcbf8f5f4f00a6115e21cbe43e9a4f898;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77436c378c6d65b69ba939bc858fd22a0e1be7f927bb5b2a886c6493594e3487;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he81ad630cbc8a7914d75b2de7ecd8573ca952babe3736b14b81159124250d354;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7ca74f01c626048fcec6f556ccacf13c075bb8dcfb1c401f4d5b8e3f36fc05d3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd4b554f8d251045b1d6e32d7898cab0d3a67100a8672cc2ed22f6745cc436d1b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9907f9c0011de799877e9dd1c3121015c25d90b87edea865565ef476818f4b77;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee91b3c5f5f21ec0768d45f5e233176e4ea491737f43a6be13093783c14a5f9a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h31798f4da97f971733ade6e47c40af6fb04e1b8449653e83831363502170e803;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac0b49ff4c961aa378aac4d1f8c6d03b5fed85e3c12c83c4bf06ae9a94b316d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6e503bf49a826b606bda53d33fbc95c41d844f497a9309caff3ebe7628905153;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfb48f43e3f896ac68197c9ff3f5610c61f2cdac12f4961367a880a65f22c990f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1ab7636a31e8549755390e3519131813c2c9c6653394693e3905719f0c5d3c5c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5ed6826f559d9dcf82576c8aed5e60102d781196a64c13c4105e5768b89c964d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7ec819e5a8194175df05689bc210d1e6604787831552a8807a072340c8999617;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h69eb5e3bc27729ebf009929664dfd32d39815b4f5c038e464018468541e98e08;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h74ed743a94f41eaa1f78f75fd7b3583c765b3ea6759a7922f954ce147c7cb7f5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfa3a919632e6ba9bfe97ec47a65e957f2d013aec8f466a94f69c4eff4c5cb7c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6be5f84a85748af9a1570650c85b79895b7543e2823a9b2c2b2efc0ee651d36;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ce6c1e3c32cf8754de1eb9394abee43612865ae246467db5bcacf2426a4186e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h61990f197b0b066fe31117f11c661347eecba7c58a2654ef2d9496a1510f85a6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h32980fef9b5ca31fc7f4d4e265ecc5333d0bb1515b17dafe6034f32584763403;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9e304a2d5848a2bef599e2bce53053eacc4d9d46b6897e3a5be50cfbbcd876fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf310b2c5986b778ccd9c3fcd49552dff633bd05c23c131487ec6e74382d9af11;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9c0b8322e61982ea0130f154f5cde7eea139c0ca70d90dd349c9ed537ecfc181;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf327890945cbf32de5bbd413c590ff8a60ad0429a36ec17eff45cbca1ec94a14;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h829159953c0e0f7bbe9e239c7ebb9d0bfe33e16646d3d44db7645980374b30ba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8adb1b6f7d11d71e88ca09132d222c4e42f9acbfbe1a9d5ceb006de17d3303ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3d99a490ddb9bc732a984f6fc4b29f78593e0ebfe513219c1abda5a7d74c43e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hda7eced6742cb7c12f9c1464054648ee6e1dfdebd52fb2a3afde90661922cd34;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc3f59c73c07deb29d12df95f78aa8e68e59540451c708315c65d02bcbfb3854a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7fe76751a5bc634a1fcb1e3154eeb28f1d984c8c9efa997c91b600bd59fc0c47;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h24bb1b4b16d68820b9ba1bcc202d3e14a73564b7cb83dac709cec0ff6ffde031;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8c4bbc7bc83f83817bbcd9c122551b4b4b2d3b7ab11c92b96fab84016af92fd9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5f05b74e444c8ba3153564d5728764c34ab5e8c3a44a48668a79f247a75ec99c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf22b5f91c3439a1d4b306a8bec9f4fd9a89d30dc5547f0f37eae0cb33e9be324;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha2b8c8d8c8a81d42ee35e81edd15768f51e4fffa455515f72489f4257d2017e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37ccbb029980fa1017b64b9d67e6fb67fb81807cf9ffe3ff2d9bf257a404efa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'had2fcff57ea0e63cc20a51a9711394fed2a8e23391ec6db59bff8db91e554485;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2580b21770df220d6950e47d09f89d91243e53ba25d606b3171f21123b5b052f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7e2042d16940341221ee8a17e460e42a67703154c32b7ce783e0567da5434cdb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h37b975ff5d503bb5f95479abbc7993615177934d81e970ece4d70925af3d847f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h33b2fb14d7ef48e2f1899246eb7ae5d438c0ce216823a21b64fd768b3771a3f8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h41c97356c4de8e020324a59e746d089e6d248dba8e4649a3194042e1fbc715f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h83a2723eb9205236e53262194a2b71f399ed6ee6333f98745a4c43362ca36c7a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8ef6dcad71150421b033e3d284b3d78947e4ebb2d138536867a4451685e9d85d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3b8036f87dc8f23b86d1ce49c4e412f361e59c24df2f97f56825b0adda584232;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfbb7c1007b2061274920af358ccd49ffa60df92990114ab2a2d121e019d167de;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'had670b86f854d7016e9e38d19e286af93f83e1df593b21cf8b28467927d29299;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb0a0a9b687e434b7811fb12cad23b02eb34a4bb6326e16a8bad02776420b63f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'haeb4abac6b60162569520ca636c302def995fcd87f4c90801c49394993710cdf;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h75b57726796427f0170aaf65428a26205a8019ab4661244a9a91ab3be2b563e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c4e6923529010056d994f8d277884b54bdb1d5c7d608128b9749701a6e91834;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbcb069a99f72a153ec64aa3881a4e36483e7ef5bb89ae5ea31c7138dad077760;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h154e0243574b2b004dc76ba0bbc7ce9b0217a10bdd93ff87c32b0d59b40d27f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h70495832ec30935e4d6fb2d8381c54b31462872a8179c363b430ed47bc7358c1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha760e8b7a2556aa4674e61716908f7e7fe198171b22d6397ed003e52fe62bf21;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcaed8ac51edc8399edeb9b76ad60d0a4d75b7e87ff630ddf613bf7fc52a703aa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd4131231fb993d35053a3bd23c890f299fb037309368a8877abdc55a876ceaca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hac9eee1c58131ff001b566ebedb7d9f63ea3b0baac52da6dd2350f09ecdcae58;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha718648c2cc1ae8cd5ec0f6a025ea00c5b28ec293ffb7d9197984c81d32d15aa;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h89d490ae89bdc17fc541057e74a07241f259582d61957a6cc4b9ddd3696e2d88;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4d68fbb661cc02bcffac5affdf30c2bb90d2e5efcdcdc0f83ae0ad40f254a39c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdab7aa6fc999a3dd74589640e9f96be32c1459753d888582725eaf414792db93;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h36b11edc4321fa7b28c2c4614e6036465320374ca38e9b1959b461225e19aa4e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7d290e366d2b69a692104621d3546e0f093c8f37d415960d380c4680b06fff85;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28c163813ebbc9803b13c1ce6268775d9217e562bcd835ca1951054f4eda07e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h23ae2e8cc7a649755dc37d5822f9cff144d53fb1eaf8100e8fd4245aab88b535;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcc7f020e6879c3db16c2083b7c77d4359a4b97d341e66f22dbb7f2d3ca4dfc85;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hbc4c730c9c0d2a2a4866c287e166c9e48e6401135d876bb2b6953983cd1e5329;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha62b198161edde38833b2dac8ccb5cff1f9c12f0ad80e94d9d7145e29fdef2bc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h615d36224968ad4f758d43b0681892bc902ee50f1341ed2edef8c3a2f0ac18be;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4cf1e0699719f2c5373ea601f907662c6fb6ff9198e4e24d9e01524ea725928;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h166103f5d1f7ff11449d0a198722b50aae4743fc5fe17dad25610b263572aa16;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2300b2e52440671622b1bde475de00725370b8f998bee85a4b137d366cc39eb2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h161d18b60556a692c1587c96da52522d540c12a14e726e811e686986ebb79783;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdfb55302086246a379e7ca9302f46ed8b7b5a6f0ed1c95dd19db7f8d3facb39d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb6d6ecf06c3ad156b523e123687d3d9081ca29dcbb043c1cf10b8e551de8d94f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hccfc83296ab16bab05d84b2b31a082fe5b6a32a822cf0cb5a933e470cf97dd1c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c67a261483e95868991ade9e4b087e937eae9b9361a6f8488e3ef19aedf2787;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h752ab8c02624d3670601a8e23ca22143042014abb98640b5b734324d7e2ee592;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb9c89d354fc3f55ee61b9c12d4861cf5dcd3d37047295946fc124bac4434cdb5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab11e1718c057f7f7fe6f1821c7d8f71d0c188289154b77422c22cd819729014;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hab7695e3a9260a5da5c3a22da478057d3622c018f0400b414227f589083ea18d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2c2b887b5bad3b9a2a786ecb9fbfb015851071ea4404fc78788853e5ccc63938;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4755d3768445ce1a34f03208da3903477036e12f2a5c19732a53044a026f789b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h4f6ce395eb0a1ef083ca58602f4163e5bb5e1d468f1fc5f9eb7a35e5c3b73035;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9a54fee32cafef9b4676c1dd83c6df4706cef757f971c3977821c6f0e2254694;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hf437d78393829e1c316b6b98468cb6177fbc687cdfa6afe71ef869c3d16c5d9d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h9747ff77602a6613ba93513b49774fcfb1a5681eb5581349554cff5f84254769;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb5729c5b6ffed34debc492757dd669c35048e0b918d7bdbfa6b4a8586ab005b6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h94cb77b73c29a405f0bbcb68defb5782a0dda9baed55ed47d0b1323f169d8a6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'heb85305f123df7a08e3306bb17335d3d261741cde5be6376a93ed01af0f7a7b8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h6b63cb96aebe4e078517683bea628d296af1066aaf4b4e1be1fe7e113c06e00f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h887e677ccfde9c581471a04721b2e64fc9b3609f0c37c4ad2cb9534ff43e3c93;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h236deb915cd47115001c8f97917c28de26c6436eedf87da61f9ea9c136615404;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb92db7ba7f1745999deb7a067575e2309ea62e3dedfd57ba6903dd163ae3dec9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hd47b1c7b83f273ba8d0918d3a1e5ef9e47eb1783df6b051cedb86b47a3317b46;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5bf36ab2bcacf206279455451dc0794722b066ea6d93011d3ad9c1ad31cbd691;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1c2f802e7f615eafc5afb7f9a2d19935c60d608d4e0380f51983d31054b4a34f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h11c419066c50aff597a9fae4cec5cdebcd1789cdca75bac9386968a0f8e53096;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h17c3927981fe9f071bb00c73e3f41ce77339a1777a4fca1e668c9ff362a7caac;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he8bfa6b8d4258afeb320b87e5aeee2deb326e02e247224c24eb8102d375ff82f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7a9f542b19b7f3d7619aec6809cf639c9061cb15ea34f9542e3348a310728730;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1a977aa1fca964c45d6fe10ab973207010a84ad9d924e70c9d81746a8609f304;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'ha924efda9c8f7dc2c9bcfb184b3bbe489a0cf5759dbf081d8b7efdab19894be8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he6e25335628eb308f611c2c74b53632221cfa7be33d7675a99dca45c9add4621;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb002344f9baf5aaf597d27a748e2398973a5dbd6e022f6f6b19fb1b387c3d902;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h3404fbf4dbdd57254ad0e574b11d9c6c3bb69ab44732f5a1bd82652862e7a260;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h32575654d589dd38153673ecc1bf8bf3ffa6420728be95c8c9904cd73ce54a71;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdbc9061b53333d8d15e7b902e41596dc7e6dd36d443e58e0d1c6a356cc58d296;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h2dbb392e7b92080e59165981eae37cf7600f7d5f54b8d8c79b3e8f7e302148e1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8c0a37e229a3d456ff8c3d899837629970657a6c0721de95f678733287dd228a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h47c2c73777acb755703988875f6f338e7345b4d02b58a2268df68e901b9efb54;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hee37f1d5ad1b7ab4e328da7d581dcb704d033c0c292bd2892a5ee71104540970;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h360956e00860f35a32fdcdd61deb5daf437bac5a5a5ae3a6bcb59b9c83af5ea4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h61e13283ad074de04ae045abef93e413e6d45318e13e2c7042b22909cd45248e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h69132932b6fc4158114e9150611d9fc8e73055919ec3cb4333d43e30cc5d6879;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he576d0ccfd408c8f1e9ef6a7ec0935343664accf3efeb15d4c2c32d45913e282;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8023115fac1a62d3e5a127f46fd962be33c47f8d84e7d464fcb40e7861454c7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h82f8a8420e4c0928507aecfce9a990a1b079b15a40303599a5d9b20f9ea3af7f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h8438021c4f4fd7e0758bd26119c8521ed5e838e5d5fce7124039131072e18a90;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he55f8ca8aa13901c0bf50b665efe6632f56b15ec293e63e47c4c995d03cdf7fd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h5625887aafa3e4bbcea6797f5f98ebb7e0838e4ecc3b100bf690be66970e750;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h1aabe1873002252ec574d19d0b8dabca43e095a71ac027893c525f9a3abe709;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfc4b88bb49b18a40ab08c037293812061b19a67d2e6c32ded57a465acfc0e832;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hb7e9eb93ff40410fa305c0bb8b1a1a402262e87f31bcfc6879ccfc14dfe48105;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcfc5e8e352b97fe9826ae0a1dbaf81450a1c6b3207e379bc97caa981c92e1cf4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'he93e64c0a69adcbc1a542e689f3c5cc3ac8724286e9623f555924ff828d5554e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hc5e1d7962a727a39b79e4ba09fc0cca0ebe21e84d6c38f775640123fe49af3bd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hcbde2a52bb75c372e0e26ce5e7f04c4968f58569e71f2f74558199897a02a1ea;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h77120363b38f4df69cc5d6030fc78805acce4b9d61a3a93f935eb74705c0267f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h28fb1a72b6de4d1b772346584d1cf7036cddb42099f3c99a982f017d37d51755;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h483264e9d7f75ba7b0eb7bd10091813e08185015473a731cfbf22015694c3b84;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hffa4cf957bc4b232765881a0bcd2681ef9775cfbb5cc02ff3d942615bb4e14e7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h35b9fee01376eb5685cd40faf8ea190ff87a7fa0216615de81b028b97a8a502c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h72dc930adc3d3c6b9b691c990495ca0923c0309b621b11f2a0efcb6f62b49404;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h52d6d8b416e3272c9fa773f69648473db3c2cd86826d6a50d6c9dd0f19a8da6d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb34d72237154cf32be2eea0e7868b0513a8af2bdff22c5d22315f10bbec4d93;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h7b8f99aee04c209a6172381590d7b1c4b4b34183f35931c6502089c8c6786a50;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'h12881cbfd33bddaf2a2893e5ba17a4953a340a2b10abfd971fc0f5aafdf34dd9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hdb9d6b27e758449c38a3ca2e0d3add7dbf206dc6d33d7318e67355b1e74e02ad;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 256'hfd63adf106127e0112c57605ccd2d82cac5a6ea97743665b3fe36f455ac68cc3;
        #1
        $finish();
    end
endmodule
