module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [22:0] src24;
    reg [21:0] src25;
    reg [20:0] src26;
    reg [19:0] src27;
    reg [18:0] src28;
    reg [17:0] src29;
    reg [16:0] src30;
    reg [15:0] src31;
    reg [14:0] src32;
    reg [13:0] src33;
    reg [12:0] src34;
    reg [11:0] src35;
    reg [10:0] src36;
    reg [9:0] src37;
    reg [8:0] src38;
    reg [7:0] src39;
    reg [6:0] src40;
    reg [5:0] src41;
    reg [4:0] src42;
    reg [3:0] src43;
    reg [2:0] src44;
    reg [1:0] src45;
    reg [0:0] src46;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [47:0] srcsum;
    wire [47:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3])<<43) + ((src44[0] + src44[1] + src44[2])<<44) + ((src45[0] + src45[1])<<45) + ((src46[0])<<46);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2c0c8a3dd32ccf6994b473879dce227ada425cf83dddc95731052588028724df3d15dff36abbdb698b20c2f80e8013dee650a9991e73fe20ef0fa0c4ffe9d8137950ce64af3fdb9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h371c5dc539fdac63926c0ed96859a25332977de4420c52b8674f41947858a433f49b3a1aef5ba4b6c14a33fae1c3d2ee619d72a0d32e313b91d4e5ad15b045d5283bb022963c162f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b424b776d6962993e3f33d0afe70a4a9963756080c6ce6894b8b6ebaeb69b899d991d5f8b5536e0fbcc808a1607edb5b83ff3da66f19dbcf5a84a1f58899ea078092cbfa213b646;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e56468ad1a96dbe5c329aefc195aa1e4131052dcd1a60a07c51a9d544b22eeea43dac4aaaf01bde740770246eca625e4dcf3face7bb9beb6c97a71da9a6e7cac6baba09adfbb74a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h84357d606b43523be67989725bf2cce2f0e7c1fa1f6cd2282a7317a67626cf7d0cc06ab8998a2d26e676f9ec97a1a685915f22e3137bfd466094356f8f9bfbcd96d0d0d063e3ab76;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbafe80b4e07b3682f1863c10c126ba3a239e371066e400803782220f4101bf5218a5fdfcbb2d089d922bf1d7486bbdcb201c2294c51afe87e0dc92832cf7cedd4ea6af1a213fef52;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe51801ce5644ada92a1731048ace6ca4c104ee569b032ccf9643c9496b45857e12e6440b44e480b46b1766b61f8bfb66a903483810aa7906499897a5a44da617662b482ee93a768;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4735a77d79cc6c5397e05db6f537a6b661f87bce80223151467da11d73d05987948405d8267d4afb4662c86a9e1d1610f6aaac558e99aac28be5508d22422457a4b8c6dcbc4e3323;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf5095ac7cc502bf8a874679a6350065ac268864f18ee6356611f7959d27c1611af67520787931a098252948d02d37f392c4e7f9819b38a71cc8711deb8a3136bc1d3fcc7ca8194b7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4fbf680ce5eae316da2399660d1eb086c3d94cd7bd6a3cd63862f805e887fda42e450d276d14a57ffae6f76c203fadf5f045fd3d1ccd11d830b4c2e511c25951248d0cb0cbec8f66;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae0c2a41af443985b8e2a35831ba338ec1f51335b95ce7c622162ff0f4ddec200a36e2b22ea91ca8acb2fed0d99cf5c17466bdc97f00b2789c39e19a53a8fab0b67870b778988fa8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf8427a3df84ff0dbf25ed8af4ae13103b1061be8d212f3a71324edcf60d78b6fa3a2abd5541b02b9f73c24e04cd8694746739b9881e488a80c451923e864dff0a6df796cd36f0cd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed5fbb3041df0d9570ad4d37eb34cacea79ea8715310ba79129e98fa58238bda7452c99cdffed61ab914847e2c7ee4d43fbbe00ddb727b014d8edab4a6395a2c09f195159df751da;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcbc136a08c50e880e5980a8bb1fbaed9a80436f2bb9fdfc521e20b71f1bdd46120d2261c35990b7f1698fc174439eaf2d8dd9164e4eed524ed238f7c1fe8a74a98e360971d90f65;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe822a494d00ddefa2fb8aef8f9c4298fc4b802aa1dd2b1f4d5766b282ca9a63c7097cd9f9e4c867a30d2a4179ca7d645835923c452384cd7cdf11be35269207f14dd4aafa18d77c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6613b9e6b5b062e870882b2efe2dc5dd12b132fb44973212226cba9879b9684cd6069e27d67aea96ae0f872d88de748515323d38e7a7c60bb8343a7e99cc6e75dabe8b71dca8c9c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba9346da88f4c3080748a53019e72063b977e68dcc3c58e15b3b700ea40d191ceab811d7ad795fcb5c7ef6db0ca47d5295b66211a01d0881bb72f09398a5f97b65901647c49a85ed;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e75d6c44aa58af5155f325a8fe519737a78182401546e68165d0c446ab2701726515108b7e7e15e50b2f9fd86fb653799056f78b8609d080d0b001b147d713a76ac2e1f66d14708;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4465f7e206a15a90e4754ea023eadc5a5884bcee742b3ade287988df9898c92fa949deb512067652f5cd12de8af3c2b19310aab5d0bceb1f5a0490f4f0b6b4d3895d924c8a715f37;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb01dbfd8c7cf7a89f9b537f89f1961b0293fc6612ad396cf77ccc0c0390a042f5662be4d303516f8d525a30ee5c937b687c769eab4d44f860a6da2dfefc51a112bacd7a98e9567e8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a2d112ea553d22177a5bbbda75d779f42d5a7e8ccd1e10233d4704fb98ca34528a2751bc2f18f378093dfaf71d16cfa8ab446ce2625690a1e539dcd3f090942d2bd6b2805dfafb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0dbd9e5657ea1a1859dfe8f199125a526478cb9667692b020a2448e8168814ab63e3914e28a5e48736b684506d4a102fdd0e0dad977a21f4953af89286744ba538fd6b09b6d3b26;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc24ab51d8554b125bc2ab3c39a4f25ce6d6292b4440a547caf10a8804762b317f595e79deee3b6662e77140e85fc13fb3517cdfccaf341e789a0fe4ff3b345d8704211a498b1a1c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h33f2606a253aacd6f06d1c3bfdbaab57745f17e5063e73031a9ec6ede15a3825bac307125955260f627b8a77c5607e0b50a4fe7b9a7ee9723b8c8c59d1574c3830f104c60c357645;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54b5ac2e91b7acb1ac4cb75dd8d6db0e0b1e787f3fb134cdfd18a3dffdea94efe01e86f2727b99b2ae4298f2a00ec3d2a0cf2611f7e3c5f48fc9a8a453c7fd4782286bd30c297bc5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd74ce4a513b0bd0e5d190fae7c127de68bd91395db16e447e7653e5e61841e27dc3fc5339f1013581d748eafed295b34cfd3fc5f94339297e46555d7a45e96164292455cd47fe29;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2bd75882599b8a5ea708fd0fc7c6dec3a1c7b24ebb3777b04c7b3b3fb4165091f7b0a12cdf9c15d0ff08651f31839aa74e8c5f8e8d16ff7fe473c5d29fc59d1dfa9a87b2eb1e11e5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c650514b04874a38e5a49add1bab8673a0af044328cfe8e7cc8de8294b1f4ef4900125c35e910d8558ed919a36fe6b895332b8bae556db6fe93365d89e15cbf40eb49698620f50a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf80539b6aafad797d8e4707329ab10915afd4e569927560c1022eb45637b29d7298353b39d3a130228de874c3d5fcd0d64e2df72499794dd50557bd5013a0221d0d0deefe37c4b1c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h459e7c5ce32ecee08afc06945f3a94fc114c2fe16b7c9c7a2824b4bed6c06031a7673e4349dcb30925c2d57f3c71a4f822030611f91f1785baa7d218db244e787d88c0e502b551f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb99fde8aef56cab0d1942afba05e1271d94380ad31dbc665801cf1fdfbbdbd0fd72f75e67d3f2cf095423c9be3e8e3441f05ff58d9c4151ffd90a7d1764bc52d895727ea2214a707;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h41fb142c33c9dc8a420cf286c7ac4f1a922a691ff0d078a67c92cd7c0355d3a68fda0f8bb093691e0c4b04b50cc75f7f3eae42c88f868e61476e1c26e572132a15317d10b678913b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd41252c9813c3cef980fea0876b8876378030e8b9ca261b04ffc6cd38fb28020461f28119d3a83d1924b57f6577f704f2c7d2f444b6db3c97ae555edb9d8b0131556e83282f1d7d6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haecf946e9f3352bf754bac5533f73afbfdc5bfb4693d4bee4b24c0b0f37124bdb32e3fce174d5b6e57ebb7175046c1944525a37e10c7f66adf87d77caff27d3d994497945cb2c528;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76e283a02187b8b28fe5785f9834b6e52a9cb246ab4617da2d651e9c5aed9f402cc8746e7a8c7bec1df8c2dd20589a6fe508b6ced1e7874cf4ad863d439636be5e24a0f249ced784;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heede6a2591d24d5cc8120db335b45be7a1adaa0f2b09c3bd8f67d89859f6fa0fc099ae6e7a0231a004274ddd45f54c46df7824d8c5f2815062c8035c2639f16b4f392c1adb795a44;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb8aba5b855666b5fe2e252dcca26ab2f26e4fb9655193bcf5d111268458dc97012ec0ef3c0a3c097a6c78f8a5f13ef61f9c79428108a6f7ca24a222a1180e5f369857a81fa12434a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40b39dccad891014af458f373cda0e534696ed7eb0fed40e660c948359755c0b8129690552a1822764a3c6724b1c32c4a9183f7607f4e83679f58d0e83edc0595833bc6f063089a6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h292f51f39d4b3b34f5828740cd1d8b22b6b45ce69967ae7a952d9753492b715733ded0594b71def1fdc0a547cb60dba472c6f808aa03d300e229eb0c015240c70fd61c26d1bdaccb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h244722ab008da122d7aebc605b8b0d706495dfd2098f716fca0a700aa74b87f1bb26d58dce5f1cb4b25206c1e130e297d8679de965839fb958d44082a0a6f32d029e2548f94ccbdf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6f4e2808c4241c344d093ce3e46fb54471652467cf10f3361a1ed66d741e13a9df2478dc574e71170eb3f646aa8e131c78e9bdd33ca7485e07a4dcfa2931c97e95f37fc919aa7c5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habf81974cef0fab95ebe66d00928add9b455415f8cd17c49aca591e71cd4612a860ba071940d03a298e528a9c3941da1dad8580a50249ad564e651d54c0f631ca6afe82665aa1d51;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e3db5cbb642899d7b4c12365990a401847a5760f3f48e2bc3d25e3be781cf0cfb67e9f0d253b411b3cbe639f5e55f8accc8f72eb9dac1e97b050875cae5c1dbc444d76e811e0581;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf757ad724197543474d69d7eb65ba628333364542163450974b0eeeb1cc456e2295db91e140064c9cec400d28d5d7d3d12875f45809df357e92777b29035b8971f980836c039d4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c84cda56ffa2be692d1c5814db7e6194c77be43af0fef8684414bf3ad0e29a4835ccfcd127e1567f5344fb15a3659a94ce3fd7e412a9e83a62064747b62fe080122ef4f4772a046;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff84517eba756b2deb3c030fd0e232a78d84cd52e831f36e02c27c3e7c64ca972885821c650141a04f30556d3ab6e8ba777b1c2dc915e1437645a03a42bfc5be9443e7a741ee0138;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd83b80364f7ab83366694c82298a4bbb64d9b198977b5736f5d1fde7547c8f1d93c3757250bf236a62e2228537af967db5b53019272092ffc6e75593e3510a05d8164a2fa23b7bae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a0d7d62a6b9537e6c918c5061d71eaee01fef94ed8412f296aba821a199ffdd161793927907bceaf5e5555db075a4796fcbb9051fd7815a1b774dd21469d6a870b12cdd118abbf2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he8be0d07a3629515369e7d5c82b050964765b347be15b84f4e00dfafe0680a1338859416761a3b36fcde12226ac0eb0f3715a1ab37d4d2fec81173ae4c0a5a05096116b948c65b78;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54ba716e117d9de7e4df88c4f3447b8e8bccfce1f7d0cb7492e888dfe60c9dfe06743f6a89b410c4ed307de7360b687b7fc4fb647165e6b70b4fe8def01d143389c9270906d10667;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdbb403aa46c43b9efeec31a490d8383b53e259a7e85545bd185144362631d7ca2c688b9cd510c787f9902d22ebdf25479e55c004714a5ebd37f546ccfa5411e7e819141cbd54e4f6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1aec474902e821a0fe8d422e1c9291d815cae7e32085428ce53d4f95774a5bba96ba4aac4b61e5d2ab8d89b3da9ca1fda165965cebed35ac3140fadfb5920e6d1b9b4bc47795d2fb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf290cfee02c8a1bd8611f93e9522d4affed40f0c5c3ee542531d7e99c57ac5c8c28ab3df5656c7077b5281b25cb0c50fb2773401a48622e65ae7d8ecc002b01b200fc5886fc5810e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd0681cee036cd358a7195234ac9275f48e9d0a50122cce6d288a54559f4c908fa0e71ae077063fe9be0df6be10bc6e36e9a416a425f9284f60349402e2b27d41eadce0218b92e78d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba774b2037d0563d709f2e168de99184c409d192c4b1a701659947bc6019fdc60f6fc90eddf224b31d3efb9c564ae766a1d3a6c6da39de65e8bf5ec59e6a63ebb29b2a525e1bdeca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83766cf72514263255d2970a8acfed05f7de6c829b8cd19888f8e37b6b2b06228b1761e2915e2ae0add0141d8dbac412848577967e9065129bbf113810d9c5c10e3d0073c2c2e010;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h258d4e95f9ede2b714ef0de4fea7e678ad4cdb8d5fd04baa1fe4af2d280215453e71c131258609d4ba15eabddecc104f7527124c6048096edec23381cc13e5ed4544fec90f71607e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5151b302ff29d9a518587ed2274ab1bcf4cbee8c72280bd5df1e4b1e87cd1b640f8109116cd07214cbe221504f6767b7ede08d23804621a29f97080f79bfabc27697d5e07809d64;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf999ba962c163002d09ed3eac2d69e482dae83c90618e1b4393b6c351050a80a1e0a55b1547291d6935f1aa23b7d87766171564625598adad45548d365b145d289de6d7b130abb27;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf84372ff24a656cbdc19db671a041f2f8e28f0ff62bb470fd7152ba84df1b9bc618156101f7f9a088f9256275452b1122f34e7fc4b634f2a77311827572b1723eaef089bf9690acc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8fed5c77191d2b29f75878d68215f0371601c0f62728b839d10c11a1be5323593c7660d28557150f2a2b67824974e3a90325e8dd5c90335e32fd674ec3bb5dffea7d5b8903e2e8c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba4e6d1668537e0d3d80a8f05ae9e6ed2afd557f0b89d8e2063bd3ad878a155f200a9e2cc01fd4ef1c4177c8f827f0805c45072e907f7fbfa92f67f39514e3179510665e261d2b1f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9999465d1427b348f8e1b8daa152d390d12ced29b67952d3eb1d2b608bde14a700b3d0e04894d19265351959f13ee98fa37c7f4ab9f481561f5a420420e9fac5acfca337bced2105;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71028475b5b3be6f5bd790d7189bfadde19845163119cee6678633fea5878bc993cafe59cf4af01c6d419e583af6e23ec24a9fd4894c5539692e599fb5c53f181450df47f758ed8b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14fa887caaf3ba892fe0fec25c449d9dcba0066559a25216a66f0534c89f66507da877ecb2492a160397afc607d8287f6c265f425f5d744e3e2cb2a7c8eef31e541934ffe7e1cf11;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7ef06857b10253adb82e43e218c847b0f599cdd4c7087c40e26e93a7ccea5d6f4ffce483855aedb53460b270fe3bc6edac816cbf1f9583f871fac375ab3d566874e2f74e03165dd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5baaea9f69b1b39c68feb050f333d9e34e6294b8de46ba22ba2450181abae238cdbca007c4c47f209e8e2be848b355664c188bfdc5e4cb2212d93ecca0ebb589fb132d7f30d60ae9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf79937478afa8141af0fb7bc4077e2d858a8c1598029aa363f08c7eebeba09415e6d74e1862f5b31f09322534fbfdae2cffff325b088a5a725298b0b05f7013c5508e58618b2f18f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5c1e658a4c290553d8cab98118405169a73b3e1e5a5d8b3edec6ac538d486a1e2a0243d7b2fedc1c77c9867a0acc5ce03ba78acd7f06fbfb82de00f128e49318941d3e1d522aaa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h277536d727461454a202e4361c871d7476fe0b2006520e653dc1b8d2071cd3043602cd83480a3ed29d3e13dd9f869475faaa996e8f1cb357edaeabaf57851b08ca45a6be38b83e33;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca75926560784682fce2d872a57b4676278783028980ea25ac159579c55f7e770faedcfc27ad9c61843fd69f8a55afc431a91d256164f7b6a041bfa70527ceefd3c8a575eed2e35b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b9e9c4ee6ebe3cf052063574a1b1e9f753328cef03a0442969a7346c4ceae408f80078d88bcd09021ce31d22c95cce8e64f360ad1ee00a3a9c6d2e2af970c65fdc43cd2e7fe3d58;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70a8069699b8d860d256741f0f3f7be7735315655f2717b3be6a9620c45db32fa8d71462c222dc090c8024e47ec5f51d5e41e3a89bee19ff47c9985c3a2904cfd9f895acd5d94d62;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ebbed80e0ae3b7e3208604335bb04b9efb49ed0314ca21f893e764a6466d299731f677730d6626dbe13faaceb367af07f8449c0e02755b9b5bb5f1c47b808867ca8a0e753799b13;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d3abbaec214517229476c1c636336d09dfb39798cdf8e2466d3981d017a6bc8dfcde425ac92d8c8b77e46bb587bba4ce191c095eeb15e8f7e39bb5950526420c487668e4f704b80;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc187fe200ef6622fe1d3fb64c02716ac11eb0a8c16d92e8d32c347f560e7cb7d350437dc1f3038450ba56aa8b38fe97325ff9817baf4f7739aa92ef174798e13da91e48a7de01364;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c4dad4105a41646b04746fa77fad54caac0601c46b515e8a1d4cc706b0625c910d513e3890e91dcbab56607eecad911322b8f54bffbe378a4f6e76ccb88100396fdcea2f82a5dbb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b0ed11fdf8e9a715a98a429d19505827ef8fb3ffa84e2db2ea5abbcf1f3400ca7f501a1e237c474be22c8c120f400da540c463292c5a67f7775484848ca4a1c07bf9777b1ef1f58;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h12a3adb8f2338b92a8715c489ad26641e5d80b018101a775c22b341564e7850ad27f07cc5fcafbfa8b8d5ffe482c4fd60ab199fd360c03603def36b740ae7d847fe34d2edefb3307;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b245fc7dad38cc3966799074f4c004e69f4389bd76ceca5bb9aa20cadda354de6639ec9ee6f3cb2411826aaa85cacb04a688237586532dd43800a63090ffca5b15e96b2c91d2d4c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c5f81c2d19e910089d9f971a7614fa27fb7487d565e9b91cfee1fbcecd1a5dbcc51a907ab43132266cae9ce0d56781392eae7fe83ba6ede4ff79d527e0f5e433ff8bc196f7de39;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h75547b963aa2c65c3bfaf43c645184f6e0c5529d1e9519015b1b30b956d44ddba33d36ac9e2d37303d4144fa843ec664c73ea68e9f2af7b4cbb0a534cdc7f50fd4bc62a06b133db6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35297de518ce6a3e64e598499d75178bbae2a472ae2f79839b922877ed5ca88de9a6dc567d53526bee987b7ef36105f713b6dd4bd6c24f068bc78b20ed566d9bbad66f66811ff0f1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h238fe3cb28289a08dc0f8952710da0a3c85de6ed9e195b40570e5df3efdd2adb735485c1e321fa587b49698eebfb16f45a1c043b2cc69859e1e30ed071401763d6cd1f45f0215b85;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83950fe936382dcdce1237c5e38327fb16005fadc832a08e6830879ce43e3918c8d3c8bf1506e51a6c747946374ff0dd0030e4eb4c11ce83deb65c25cf3f38ff1511a356507eda62;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h37486465498467b3111191eb2b64a0a04e6c27b71a772220bc52edcc51afb78af333e810b7e15ada73a328e3d86008cfdeb63e44ebc20402dd0cb71447df9753f7e8b12592e0fd06;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc718af3885d731d0cc1a82eebfd6f63db56e72c2fdc6f2c36a29a6e76049fb1ce09b40d6c8da6344770b45f881b028175104beb577a6e58c6bd52ecd0fa751b31e3e08e2340ca95;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h341918f852a2d6783f292d85410098891ef29f93103d98557a9cb7164e261a29a12f764c721b79efad1f42b40b856df3b3b4d0ee00155177559a924c014652f73f9abac07cb994fa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha9dcaf5225c2b325321a63924e3a1dfa60bbaa3bc99512b9eba95b7c3db42c0e4ba97c2a73088f60e344d3ff767d947686c6391b66f56ddcb4e9eb03ec5964ed6b98d083ea13a50e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h10ab3b96859c9c4bbd157117623a26fcc8328fb00af5c3df635606b4bd8968404adb8240c462b3c61759f079f7dc6e08ba15b64c9122104013cc6326154e9b94134ce1f8a1c0217d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9707b42f9c4f8524e50990e406282a6aa26c7a377d5fa176079b57e3a95f99ee820d61efd7dd3f5339850cccbd9c3042cc334db46a6de1aa5969550a550b62ddde17f4d58463c5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc5249a44f1eb87587b01e8d4f8f5cf5a32f97f60dd7d313a2e7277a661f11b97ce54373d2b9879ce151952670cc49502dc9d88de96a41b35fbecd6a403159d21a2423ea5f2d3408c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7cab0b38b74453316618c26911a0e0f13749f1b5348c8f8df0af761353139eac5b1e904b02ce912866bdde1553e202e892904b1f558e40cba15b39d1d42834be696ec3f0a0dcc045;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h527537aff579cebca2d78da363ed7981056428734f76e3b8cca683f1f26cc64bf6e54977aa725fc687dbad2cf6622c47f4b1cc5692729f32e1746818de096d5b35db8791c4aaccbb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h13e81f2a930dadd604ec98be47f2ee4dd016e63f103f1e719ddde4928e86b5164e5e4f01e65cb88c889b9ef6bcec3d3a4d817fb9acc0c524f208eb5c421da3253bcce84baf6bdfb1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcbf052a260132eaf1af82a44c405df87965a6e233447210b272f527480eaa9dfdf0d305bd583203303f814d37956c2eb2c9e6fa723996648dc3498a24157788b443ff71c96632505;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35b9dc865a8f5d11d8c97464f388e8f6815346ba9b49b226cb18ca38a127197d570f99b12de4ca112729eda3ba9736af6075d75828cfa15e2ff07e8bd40cbca07251fe516db3f486;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5415975858d67d3269d6f00b4102e95e8347f5721a4d2029a5c42c9ef19204c2b1b40e6f8eed6bc96334c621ea765f3d5333237521ef0b58c5693cef978b621a0ce4e6a0100027b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff689054c82ada39042abd07561521000fd4f89c91f05133d8bb510f8d9366b11434e76114f84ac4146f2aa0e33a33baa8772c19dfe8500aae1c787821d7975085bbb4018acac75c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29f3392e7c1865e6b426ca2d7bb35e8034df15bb03e6efdff119acb796b713d4c8535493fcc6dfa810d3b89976d8c0e9d0c054100655df31d40c4861fecc20e830ab693d1a669cf6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf6652d5c9948f297bece4074cc376c74b716e291ac37d5df5fd420032169103e7fedec1052527de91771b93f7e25112d834dd7a15f8c9d289d7b78562d9896e7829fb46e07957133;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h39ce23c0453edf866a87c6fa99cd6efa1e13d4b8716b495e7b3ffb9d57623274842da5bfd7f523073aff5d17c55c02915f9bd5594df77d220b52b6060bb896d2227ffbf99dac9299;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ff3a76ad0196d388699ccdb3804da9f383906c4f60a51463d1d8723b4363c56e98e7696d5641c9006fa71135f292d53e4932c58315f025373e82dbe409830e504a1d686657a8d74;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82f7882e5c56b69554c677461ed2b07f15e05a69ab29a370818e4588ace0dd6c6fd632bc988a88bef133ffdf5f023e802bf75dd54c6f698d676eb65023408761e847579c0e262008;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0af1245a63785d70ba6bbddbef70e004d57087bf3bb1213a2bcb7bab7b871c1b93d7199efbecc8c40d741efda7204902023a06721a6d1aaeff775970a44ed6ce1b72a6c746ac16e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51d84b640db667185780e1593f9c3d048ae987064d143529c4335545234531309ffb74ba37f62eadea255b0947a6754235ba15d983d9086204f2f01a3a80e77a5835f0e287a4f7c9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1159528f88c9930e91ab9c3b479d7e1936c6402f34ed6d72e831cc54e2a8e3be8a3ba104eb3592f6955d3fc18d38854569b91b3d6540390c93762ca1874b7886cfb925368d3b4091;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec22a942e727c099b5038231a4e7035fbdc8ea29ea3e1f4ffbe141d172ca438d3b1fd94b7156893663d11747aafddb0aa29d77ffc8f1e957f73a2422cee0df59c53d0c831862ea05;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb29f3a249a884cf44e0d5c5e74e8e347c848cc3e72bbf0e31e8e38b6bf4f1b85f4f376c02d83cdb945b7645821a06d587023ad841d1c5ee824a4624da2ab90afb31343ba7b50d542;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc8d33435da827a171a9b7d26c172e6dc55d968396a5455e04a6599e59dc991e9007ca8e5460aed8d6b8dbe4f02d8d085be71affbb15fc4981562b2e318787f566a20d9c8bdc14f80;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd741fbfa5bf384a33dba1f220c2929fbc1a4c5da7d247ebef6ec91ca93a006fd3153a6a8c4dd78074db0bceb9e2c1e8a7aa9d4c2ed83d1117265781d9661e3fb7b6484d140d7415;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e51d423dd6f5a00c92a44d19a746e6a3e9e32fd83224fcc90d16fdfb63ba3d3e95d50cee29ffc1a24e65a1c761192668e174723edcd4d5e0938a90b9b12206e6137fe47ec375e0c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a0f5b5ad0375b94dbe1f988891a32986eb4015c7d0a64693a1ebaa6456c0629c34e89bbfdcdf5e7a1db79ac8f0723d0487eb9324d7d4421d117118ca1080cb610cd6c0f199710f2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a3fe8310e5f0b73545976f8a92b99a50768bcaf946c350e59e39a7a14a99d4b961e9118f1f91ad73d5fb6cff5a95fd0422a1260485c6c622f9d1036d0bcb663820ceac366eea4cd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69925ccabf046138107b128fed1c6f429c7e83f048df05554dfed7c1382d072e549a58a34b9f78f56000f136fa6d39552f7c4d657ba198f4277488a2b4d0ee99154147e573c5b6a0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc72440a4eda0e3ff5aca33b26fa29abb8f04475d5f3c5b25247853a8527054d15a047d3d6f0a99ec4baf0eb5d251c0318c7db241b28994cfc3d2afe02ddc4693e1ee0e82e19f0f1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25043ac135cca07a755b90611f0e81b026fbe03414ebfa568d677d80ad55c3f7d2a7ce1dd32bf922fa0b0e3b998b050965fb3aa23516ba5de6d189232e703284dbfb9d905487d95b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1732005f7725d4fc504036fe18ed663dd7b03d52539a0b67d8a077919c5e2a00e42f5676a84ead689d4d39ffd683164f89484589561e1fefc99fb20ffe8bd44d39e7c7d47973657b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h364ed4cc8dc2dad2015f7dc87df24bdab3ea518bd3ee95d18a323d8ce495e82b59d86b6d268f5e4b3a97576ebe47583f2abcdc3907932e50f717701ddda55bd41cc14586385b870;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8be809648f9ecf176e0c31ed48a081cc362813acbce7b313618d18c5ca92578fec07eecd24938eef6731ead4ba607ea22b368c674e3e58ca89b2beb4e37cc5ec205fbccd43b008c9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd0cd83461c32ba4fa19834f880a830d239810887254161165436811506b0358e38ed625464797fd83082cabefb747e9c95c41e55c4dcd1e715b5cfbca5d1dba2e9dba7a1b5ac48f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb85e69a50faab10a89aefd95cd609384b71e3c04147f158a5578ca4f14e99555bb270023318258e5d93c2dff5d991aecd38b0ef8c388afc8440c4e07d0b2a42e944e7f593a6556d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdfc2351e4069c1849e499347363a9bca953e82e9ab304072bf538f6d522fc90c3c91feaa0fd456f9395855ae3cb62eb01857b4d46001b0b921b740e726cef7963992399664a08648;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb3f1a2f729b734641270e06f389bbdad094e0f8ea5f4c03966aa6283004fdb50a141ecdeb6db5d90de4fdc6dafbff607fdb284e611fa8af3967753e9e08a23dbef2d5194f91f1430;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf4bb7febe302cab90f2d74ca6265b8ba11411e62e027edf6ca5af509810eb0e2bde118d9c1fffd3432b952c3e78862451126824c81b67ac4290d1d51f6be7612a44cf9b8b62ab49;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8364909d4ade7c878a4d4b190bff155ae3e2715344a7ad5884655a24a318aaf3d6d243d924c7ee2f65195216efc5721f2a552a3762933b61314c4372ba8198a370af0a9770f354b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3a7f5b9de8a5ade77384103243edf1ece89d417c4a0f4af67096f49f1f5dd1be0180d24fc039e686fe98f58809cc8ccf1afcb6daadd82d6ffe921745da8341b8e90b03ecade28c9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd682274ee70e7b96b1b3f26be3551f15773f88072ba1bce6799059430ce7193bc5953f7d9afd3fbdd026bd36e1118230684b32c018ccdbf1406f96bfd24b81707300385a80144800;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ab8ad78b253c02d071306e4a1a32b7b99c0326cafe054f1f91d5ed0496bc0bc7c0735df50a3f7e70549db5a228f58d7ae7134484ae5986aae9162cef0093554545557457ddb09cb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb76b386b9ba9d896a3899d2357abd4d6ba3b83ec13d609be5f8f7951d55aa36ed2dd816f910f75aba7c53381f862eb9570c59bae823513ced72b2438d810c6affca4028e0d48652b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h686b9ce392dba391d7007292df02f7234fef5ad063c2f1ba3f8438b425567fa7a40a7cae84ce566d9c0ef669b0f40b499b3f6acb00f3e1f9cd9a0afcc4c17a3f8c95122bd992e4f2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b8e99ac3e7b5dd6a183ccf5bdd32c8f48152c1fcb8cb2ac38c35af48e5f55b3816b8f0bcb7850b04c51ceda80c85b925e51393aedf198037d9a06e912f2f93c5ead4d8ef8693251;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd1b642e9c4ae37608a7787aa368880cb6944e7d73b6d50a5f9e1c7ca33adde2e17d89f98c9d57f1eccb15f9a7272be951fbf04accb16b465abd4b04267d56a481e6de1a0b0ff79a4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4b616a887e4960c0b5833eea0bc70ecbedc72aca4daf83efa2ddb75cfcb72bf11372f7d6aa2aa2319541be7983b13d04123933402a5e2d2e6cee994cc7f46cb05de77eae64facfe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b45b80c268e300a8b1506e1f1dea0b7545c53e0cf1d374eff46b736742fb81443cf40dc5986d9a39b20709b06690cdf6d3e57bd4f4663d9f33509dcca64d3eb7f006dcfe8ac3b66;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfe86e0d43df71d7b7894e44f6cf259124e53fc132e95c5581b25052698821016bce29568315c89ac286af75dde9c569a7ebabcde9361c2f91eceda25665b834127b8bcffdb8b0cf9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce1dd0f5484b57299698ec4d63899a281a0e361ae04f920ba06329f4baad49509eac322f736c518cd6d9edc84b733a5cb6d8292356a7e20b751e5e5af6350fda00635cf32f9a0b42;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc607aef0cef84d1e6b35fd2d4f3559693d7399f623184249297fe2983988ef06bb9332d88dc8c5948cd5cc8c83867f85abdcc0801ae97ad1b081a6379fc9bcbd0d5544a6d4dc0421;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hacacb8cd23c9af73ba4c121665d29d22929ae62e6cada05ee84e08675ce082852748f72d1ede22ab18bf0c36da1ceabd68cd100075d40b078b28b794934e02048a8cdb988de636a7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b6820d96e347f5151c8d25b9ac2000c7b1ae6d2d896f241107cf7366c387679688f83cbbdfd620c6c7465162f55a0f5bb6245a2c053c2dfdeee52cbad64474db5f57a1b5e0c2bd8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb6f7b141fa53532eccd1f9e610232efd455d1075141094cca90a00ca2b56e89a0c3b6bf7e0383cfd2b2ce7a763c1f98a2577337fd556399d937591197d97daf158cdf32888ffcbc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57b530abb367dab2befe810ffe308f01bbe48456077e64e380eb0fc90a4652b395e7f76962578d1fd7a75893b641a5555d848cdc4d8681938eb4b45d29f8d1365d59461f0a468c84;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h17bcaf21f7458713ddce9a7362e7d5f217a16fa7e19dda3803216a305fa86b1122cb1a51a7fe276d2375ed820b0e5759d9dac06f2e08ec2420d2b7791e934177487c5a8ecba80271;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd75ade4e8f41cfcb47b1c3a73fd8379071abe36de073c6e822eb0185ce7a0d25309a38d6f62f2ce452963a05b8697c4b921904631b14e9a7c0469420db377d9f4e54ac5bf7ed667;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea1507ef17e1dcf859c2b0323f9f0cf28e6167e9c98d60fe3ec731bd17e63f974af5a5d320b1285a7fa5a9272a8704aaf2bd0caf3a32749630b28437593336cee1d751db9eca85bf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71ecb6ac46bd57031c77342dbefac33a4f963ae43f08ceea9f1bcc92d0c083e1784c5b258ae78857f624d28e32bb3001a18eccd08967e2fd608036986d908eff28aa5ab14bef0147;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f052ae9955f3180efcf26a770e70fd69b56d1c04e5885a3f81964cdf7ce1db7131050d215c21dae69e77039a2e29dc089424ca3095c49f5a9791dbc63ae6fc8c475909dc885ac91;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8718b006830bf545f6354c139929ce462ebe4f6b8672afd1f1827f4c3c682e69cc0900259e9a3869908409c1aebc2f5121b9208384f3ca3891002530e4b5b3f4b230337f8bd1deaa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b536dbc9b23bc8aa28bbe0f40cb3dc2f2e4572b69e07448a0b355b26903e666d18b45baa0978a9660664b4a9ca1418429effb0de4052aa4a8c86710079df83ca82398ca7039cf3a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd28d60c5fdf8ee3de5924c054889fcfe0bf6bd10c6a574457f06dfbecebc933cff955249946c18d9de996b3b3b55accc367a2c54b4a133013327a33bb4deee4e0d2b585c1bd1a0a1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35c1f7985f7cd46cc5a99709b579dd38271e17e1325dfcedbaa67db882c346c0e962ae4250f189529a8d12d49f6ca5a9166ad1a1b375672f5f487db9bed498fefaad14d46b769d38;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78e33a02ddef44ab902efb252bbe79a8fb74c18828ea144c5acc5d3b07734716d2a8d80336e2eba26bce2bc437ba70bc79c98c31b93ecf41008b51be51b7c41a8920e495307760ae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7bb5dd840258b1ec8dae541014902e44b5c134eaa6ca74f41f8ce6ff994804284f642a81460361b3158aa61f2ca06691edd91891d76fe04efda344ff3a99a2b7823525e50a02d7eb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7937da6ea657930c5c796788082261a78f537d68d766229617396b4dc421db70070b07560d368b64c689ab380f2adf73fcaa2fddc4117bebabe628aeb22cecf09e4c9a0e854571d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16937ce458e3e55d6117647da7eb3e8ba2beb269fa44681ee0c183dbfbb3296f6ee4370760e92dd7a65b400f6fa82271e92e36b72ffffde185b2fb0eef949c92c9bd0c7bf5e0144a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc13d6f3f5d73e35b5bf7452502881843c2e99767a07a71df9ef3f0f4c57da7fb329fe0d04c94d61add71c1cdc2cd4ebb44932fff4b42da934f74d7fc26cd6d3cd109fa3961121a9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h62bea3ac5ee808942d168cf9186771b3657409fcfa69f5270b0e14d15b58c99481edae42bc9e6d4d201569e210d1ec32a37df192a3f6042ad4882a3b102be20d03f6c5d18f531a50;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfeeffbf405bb01a738b8f6e8739b5a51f4c9357b738a4089dd3a6bfd2c47f9cc52849c451b1936759a5407afc0b9b8add521ae1d6766d1be08b8a5d38beb34a07c02c3e5d4782875;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha4b2a84d64247c928d45091830a447f944fda75b5c99c774b0f56988b25f87cd2d5032ca593e6a94d9f444d6a6115750005b74e1381a3aae5bda6a5dc725609febe3359372584520;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf091b04f1abd5a99774de2ff91ad5ae3613edd693330f34e1755407a0241f5722a5103cb2a0fb39436083189fc4ce0c6f290ce41e384a4e5072a75d88e5b93284746ee1867c69b9a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a59ba89a30c599dcc3fb02c246b64778f09789729e56ec6b3bead0c8675346fe8852b110327816abb1cf9f9680d25ee982d88642e09ad3f65188eb5a1ddfef414b35fca583412f2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h228ad09e3f9eea338f6a900f3d93b3d347702e46071108b8ecbf3cba745db6aafb11ff4d6ab3f9538ee32e80406cbcbdabad18a5c634090eb4a616c1504b378989d8c05fd9918485;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdad0121ee88011d2c18f047ce61aa319649c5a4420aaaa5381d75b23363e90b931372520f82528b7c6070d087d0f81261bc49a2e4c59b019864446e73ccc606a4ba4ea6c3c6aa1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26929f0cd9268364b1d3f6c2ab90572650a0af2b0c2d03aa3146922c64767a1f51cc62aeeb6a8926e3afd3178db9208ef547ac7718a640e5fe91aaaab756c53704766735ff2923bd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54e38410e4ad68505640b61814a020a284326a735e334ec45f8bd202dfb31b561dc5c43f73d05317dda8bfbf85c7ef9e75e2bb6fc9a7281373555b926801918e12f3ca843a871681;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1db091218a980632fe10ac494a9e126c63b2d5d733aad1ad8be64ac277169a046639eada59b5118d37fe3c5e8c124b8668a51a2ae64b705fb068ce5980bca171f69eed7c9d0c7fde;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hadd798f8eb7f22fd33baa6cfdbb3675a901e5957e974995831de567091ec916229a6cc418b400214d56f2c79c47e9c50b7c789d8883e1b575885c22e4b5d0dd42b049a9f0ff85528;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54f833de27454620fb4f01a106bbbecd87f0ff0b0438ea92f359881ecb0a974f03360a87284995a10bd12af9babe8443063e32b0ef670ff6efcf0da05fd59d335a05252b129a6a88;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hadba4394abdb11748dfac271cb52c1a40a5b1290c4ae3e9f8468cebe19beea24064ff0aba9eea8d31778015888e8789c42c6a5392e4da0a58ba8729dccf13df70a07562898cea756;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e9dd81f151a3e9d8cc13a6ed3bd914704f6f1370da7ed878f95b8ad7f6a80b6b05cbaaec5af8fc11940d0212b9cdf2bd2d8d0bc28f779e315dbc442b457b9283c5931f72b659233;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea607abb5d7eb05b0416c2ac750e1d4382ea78c4d3e4a040557b93c96e3fcf2edbcbfe6423b41a40ea1a27c82cceb774653b63bf3683aa856798a228b819f71244c471ad470b7fd3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ed6f441cd9e5d2b2367c176ea78aa6ad5c637ee8de1534fe1089b40388bc21ad69f49dc277e08bf469ef327da940e6675e9e0069e8797830fab0dd034a8dd25a97a354d6d8ddf6c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91af86c8f2abbe72e813521826ae3ced3a0efb6c54603a22c65299d6b15c415759e7e72f0635d133c32a57af040a87417c2eb9d6ebfc0c757ad05f83ce92b80939bd0777b86e9468;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h10cbd1eb479078273fe3971ff58da29dca18aa6f9dc1916d15261030bf4e67ceb26f66aebf7711fa47e4a0da1d9eee3746c3fa69544fc8acdf84ad0cd4c80185325dd0052f4d3699;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5d5e6ca7a3491d3aafae950d3154f133a0344f4ec8384724339cfc33ec051ce41f89f9bfb27e9513233ef12df30f79beb8b7b5c84d22e290279e0635abe9e7cdea50aa26b572a1c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h65f8098bdcfdbae362c5eb98e99909da0e132ba46dea0ee40c80436cbf5b3417debfa80ce99165caeeaf84c33f341a91e7766de389733a20077c451f41724c93eaef81b5a7e5ed7d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9abccc73a5961117465c3e85d51b064d31a24343776aee0f96ea2d2bb6c1a0a3e713a52f2e03ea7ded6ea284af0c9d6f6af0de46d4daca962a04579c9a227175d2f4970528a7249;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5d78e50ae442e4e6c33454d72da35da437cc41ea3049523623b2550cd5c7bb9b6c2ed1ec732290b9b8dc19fb1f9ca5b427aab5fc77b6816cd8fd151e2a08455f2f49757c75441d4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8be515f5fadfa030c181f8360a8f037008f2130669dd9158226949aa7d7ceb4e7797b1a7ed695d80a4ee71876b946693eb878190fdc9bcb4656190e600a20747273a35bc51fca23;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb04f080de2ff033bf15be66e53033c5349ce39d61ab340196121cbc60da9705e1b11f651ed25442d77eb8ec0ec7d711b2d1416e12ff0b32e308c2cab0052acff09e54009a633f4cf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5abc3acf5336b768d989577fe7fc1b1b258f98de6d54f8ffa6723b7cc5322d716d271d15898b0672c63cfea8f1ab1bf768b365c1cc4bee2b9fcf968f182f62187342fb4160cbbb2f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2168f4c515ddbe58a4f1579968d67df777e4f31368f8773f335a17b15a05070a693758326aec73d2754e3f7d92fc32f55880846a3e4feb3c504244ee324bddefec088bb50d7df4d8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'had22c8cd394c1997ac5df3173db933a4c3988c571f371ab804fcff5ce096a161cfd730a9c5153cb69a8093ec80d920b470be7181a59ff8756a2647135f5b256f30a14049bf9be083;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce9a35fa8b61de238aea146a6533ad6f6fa02a58395d0d760502a66a7b8c6e7c454137f892b119a87ca0a78b650c0bbd2bf59523bfba8cc9a35eb193465ba81b7fb67c54703a1f62;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc31977928c235ba00c6591aed906eeab70d46036afcb4adc05e08d0e05c85c2ffd0a3f4e1c2e0eb8324389ad7793619cabb120a9a2b56d00971075863de6cc4c9a729930693d2e37;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h300376d12aee2de25a3de8bf20599c6679f2a3786d6bd8992dc79e7c2b28f56a8e21290b851da6d4dc23e2c99e2041c89a75a8f346e4dafb14e22640603b67d5dd3f21ecc5c59315;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6070ced591b7234c9370b93c76d672e6f4d76a1abbb52334890dea85036d4cc7e50f217a9c02da121f85a9a7be3f4ec4a5f674ec89412c643f1dee846ec8b3c94ea480bceb59d5a8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6cf233904cf9bc0c77198d311f8b7400560a4a1b69ea3f3094169fd6e631f81db538a96e82dfd3ad59977fd9e39f344e6e3f27d25e93da59e74e418cd09f49683aa4e40b5365b7ea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1baa2aacbc02ae74dc0848b040e4c388bc868da1362192a37b519250900fcef44779521af05f952b096dee2c4932d4a6fe69e3ca01a48b45dce6183fb3108c26f4658854f594b731;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9bf721644554d60cccc89ba1396543c3aa612c696878a9c850ce8872ccecd9a7b9bdf199249109fd9153f23f79fa6e63eda4604029105d7004410c89f3837ff646eca5969e364d99;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e19a4a0ada13b2c57fe3019e6a250fe1ba0a2e97483ff77504775672da8ef712ab9f7a52e9f234290b1430872a05a18c5bb284b3cdfe658f88e020b168c3155d50920351d161889;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf504ef665608ba19806b5c9ad403775b60cdb5617e00ed770673baf9a993f75c56cc69eef39f257b2e5ea9a4800026dd5e0efb99b5fe8e05a3dd8a163fa076c08ec7969fccb3cd9e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h352e0de4c772237c821599bdcb51888c9b05fee95e8e37249c6b944df4694178fee2d06653cd82b08bebcdc54fac965ec2f61ac99b08e6237722bf15c562ba583af1beb97414c23c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20ff1f2357869308300697453c14136e25360bd8e9e34990cf5b8e614b8fd15a9be482196ed95ed7b239ffb586ed02b4adb6594a055d199ff576ab0249f8394db14ec6afcf7ebf62;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc7848b7cef955e6295785b2aa156db13245a19c2fbb0fb0182b22841c62d493192dca50ba27dbdaa3912a0a61bf1d310ed3d4c33e13875c20144b9ce1431894d593c0d7862e30d11;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1da1c9bb587007d0549594ed93b7ccbb0fee9da2c3177b03fdab839fea9f94af1b2327dbab910655028d386562a3a13361fb9ba97f69e3a2e4453073277f7984d82b37dc39f8b116;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h222ba6fab2a75e1a05c6c83df7ba5e4bd53858c3965df255732708e6967db3a948d8c05765754b70ab3e5cf63c899f9c740a6b90c94b40bf04a971cb517c47bfa00b9b50e459d19;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdb00f62eca942aab079192d124b2720a1e3a90ae3ec920ad5a911c2188d92160d1c5ed249edfb46c607c901d21628a1c8ee97dba0fc4cc1444d6f8a5cf2a17af69fa39f9e25c4616;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf1ba6a8843e9eda6b8350bc9b2af8479c14356586ca37a158076ee964d77bb0defb0d2544797779aead0bddfc2add8f5ff916c541ee8ba18e0b8851ff5ffcbdcb6ef8bb6f639c2c2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hedfe9b9716de258815672feddf9013c0f967a012af584254eccaad39a008c5394284ba5abea95d1edeca42587fd86cec24a7358a531ea48489b4e751db640e2c6ffb1c2918382b83;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h580a70db8f699a343c67cf574be389e6340e1d769434a9bcf87063124a95f5ef8dec3272448ccd6e4c1d087f2e9354e2fa6ac3f51ee4c65f24d7216be83055d6f07d2a1ad6ff0c92;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a608a7291a2dd5f17b1b7d2970bbea76dbe01190a1dbea2febb64ec6c51c4f992232d066c4c6b2c825d8ebb9629b7fb0b4ab666fc4fea43fe8873099a87262e8836b0266a075a92;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ed75200845e78eecef3da1c15c0aabbc2e58688041e523b0e8f455076db08f8cd51a614adbbc2dd245d7af093640b96efa82e699e42e077f84b879842edcec742985f4a0f6bbb98;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd266dcac67c752b1cb7e01091f8afdc4f7d015c7b9b3597fe3a3a50282bdefb0004e34d5f9d1b141ec0f21173c93927666051075fca64b2fa700553acee47b03ad48ecf081e5e9b6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ab9ee4c0005c6999cd4228564bd1abf90dbcb1ded68eec16813a6445a46f2f9ff26e1b59672b68446efcf9e82c6bf4ea1a50d2f3ebd686330fad0a9ed7a6f20afb4ffa06902680b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hddfd195192eb21f03bc08d0f53b13b712055bd5c3819fc665e4d37d510e0c106c86982267a607c446b1d37a3a22e1eea3544fda1bb8f325816dc9dac8469c9a015da663a811b66a5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4f6be3cf09c02541a1ed9c243464ef8064ccb22d966312fc20880686b587b674d86d75db34834aaf3c6ad8d2df12a7cac4ee4f0a49521c559a417054f719ee4f2aef3ceac8383b4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c5d7c365afef64d61dd4e7bb4e853332404fe3206cccdb26eaa4c9a94b6626cdb2840fc95ac973b1c84ad19b1a1a85b59bd078a24f7ca1c59fe34bba329572e1dfec51defc3f8b9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h782011561f7ded6bf83514e38fff43b25a661feff567be0d441bc650c0a2df0893265c2d401008289f256f84b3720174bb1f22f33231e043ce061c437d6b89e09fc9c2af092dc85e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba86ebf36d9eab900d7a597b3f9a586a00bc3a7e6f386bbba71e31f245d51722b2dbbbd1f40cccf8a5aeb163fcbd3b1d859ad00e21d8f43bd2998e98a36e877f0e8b7a1a101c939f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9e0d50e735f94c0d45efe7e7ed9d16b7950e90047646646bbb6883c2da95ef06c49f05c1aa2bfccc45e5d5b7ed71ea7ccb7aef8956de17a429015aa7e4e161d199bde35075cdc9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb4ce66d9678ad276e4bcad7f1bef53164ab7b6f1acea63506ac7e72309ce5a6a2423fb609a03de4cde6dab7833e4625411ea20c348a65fb2cae94dc5f5e4bd225875dae3d6bd359;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d264a2006ff7420f2d98cde803099a808dd5c430003199e287c101b6df7bd89e9dcc682c01785e39d99f92b9d4e4746ca3c8d0a94d735fecbf80c62858508a797dbafc0168b8ca3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8013633ee5c35b0aebb260ab618bf59ef22dfeaa05b5919f6cd1f179924d54596390c68a398e419d008d265ec67412dcdee64a52ae3ee467264572b9ba60920e9b20993c94eca92;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbc89752298a3ac3c3669d82ea03e5fc9ad785f26698a8000b8bee05a589759d2a7509f1eb27476815d80bda7e70bd286dc4b2ed61878445bff08bb6353a63d0c1d8647b0f130e77b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26b5aa3eb2300c5d5a32de5d3f7c919be7c4e2c3d822d497b05a2df07203a5efa8602fdfeb778abc72f8bc0ea710b0aec2ef782a1ea6bea50384b82d60162750a50829e6f77a7ad4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d6035fdec1136516f9559ab1d6f55a7ef465886345e85ccd7c2442262328a081574c649f38faac0904358033c5819fa68335ec1f152023fc746f6e62e9f1711809ff82e4b287857;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5963026d85fc9a48235147d8f43287d142480e9aad57832def3f9ed1aadef477538ef21e9e44bc2e193111eecc67f466f3450282527c13763c3f5fde672dd7dfc3a9954e7941d4af;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a827f8e4add592b45d49a3c98db400af327e025e19cac11ba0166fee7c27eb91262f8e3046722cefc40178162cd6ff15dcbacbd4883806a4ec0e18ead52856557208a85f19bf548;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64269cba0efed5e2150f3ec9f808aaf11bdfd5d2a13517a74430ffca41057faff608e88f8018f1be7153008e9147e9833a37e8036983552fbd0aaedc3d69d50a5e777941fde65d83;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6d7d016067a664ac71ffb99a945edd39ca90063973d2d358bd2cd998de033e6fcb7f0bff0366f4f51024c171d3256ff5b20ae56da97d080c3fbe64a3fb0c420bf2abd646bae59fa3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ffaed66cebdf613c8ff103752abdf42610c4f71dbcec0cb630b96d84dd6c3be049b375c7c0d2998eeaf98050a9b1e82238359fa786184579c6b81e294d9e013f43203a440484a3d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h636e8ee8b44bc3d2da64bd4ff680f38784bca9ec95113488a31aafbbbbd1b08b4be1a401ec7fa7d15d1381e5830db8dabd08d49588c73bf2676c2bbefb0f3e2cf67ee76c76c8e906;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d46d994310b6059cd65976106a05fa0f577babc60ee0dbe0ce5fcea269cc62fc096046c8ebfa230085ebb267513a1f0463e73dfe5033281e04a738a360da6ab3cfba2386c61e2f0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd956e2314a4b1e939d6ca8bb82d76c436fb49ddd529cb4b227846be35923f2b25315776a2ea43c0d70ddc27b3473393cd91de88767d42bc09963ca3aa14746fe998dcfc2bdecf04b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ae566a2e70d82e1b0111a30f4703ecdc0e9abbf752886ba6706b2de33f7aae37203c1456b3d433a9b324a779861450a50a3b61d59b912fed62e5057ab07f54a216b99ae4b39a9aa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf01f1263f0cef59c17b4727ffb49e5ac4dd6e49ac36342300426fca9cb44d51d39db107c62d7632a6faa1c0226c4afc95e4ae071960298491ce6e12a38350a48a395b07d05effda;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b709b4bbf21c3d77230713bf146aca58c7fcfb850ae42b6f4849f6f2e4b6fcf7e10c4a3aa39313da746e1f346f2fdbbcc7a8fa702bf952164f390962bd03d7b14cdd02bed88f3d7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha7acecfed508a1905646cd18f539e5e81cd25f909f9ac6b884711480b43cde0d2fe53becad9c0a5b92d8fe21af139ed91415b3951ead60fb127c93e196f3eda0ef05b20987e29264;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haac736d08f45f354d5b10dd1ccae055c0bc172d06e5fb2230376a95f9aae3c98cc758040d4b9f7d6d23044aa66b0c69d8f8aead7a4274adecb8e0cd3e911bc0db531f3c1b5c237ae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf09f9ce6199b9d3bb4e0769a3e41c8244bbea5dd5e440eb3f7d2e3e353e30616b0e1423205633f9a200214afb085cbbd6a5a309c0472200a3d84f65fc0958f271d5747f6c228bc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h139c0e97c77ac6532d3fe86c33c42d65272ce19ca5a12fbe5bc84f1e413d1c78ac71b7c99149927fcb71fc4866cb5953c4d7acd3005ae0b821b7af5645b3baae0d9f01cf1ac392d1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1da168995bbc9eeafc2b791c7061f5d9aabee1ae3e438c59f8f68ed9cb78932fb700c351a3526812fa63c674d1ac282db7d5172b263d8baf52636301e53fb3ab43c41bd166947c6c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h32974ef6d218b340acf8dbc2834e04780e54a71e80ff5ea884935c52f70f0bbb06d9a8acf50e28ba744fd3e9ec40dd82f33331e038c6ac1b1fc6357918f0fd9f7864bf32deea28b3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8005f67e4ad395c54d8887238120ed610e7d6bf74a852cb559220bb70fe8852525351493da9f6c57f5359bcb88d9024e61253fd14e8110b0695730089d6b62cb5de97e83e46eb628;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hacabe068475020439b49711f408f3c77a7365bbc41b64e6f3edc76ac997ce18e43e4f44ae6c6f8a772ff22c8e905f76169fbdbfd8faeaa05d2297c0ae922a47e9c6539125d76838e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35d9533b4cf11dcd99cd3a81bf45b23b834ddbe44cba4a120774e435ad82aa060596eb800c76426d044f4a28fd52fceb96daee18674471580b2251f0d5209ee0e81d83f939f4acda;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a8312e6f2266d9fb998c53969b9f94c635de1757044bac7cec8403f8a3bdf1e4b65776dca653e367491706194e0c8d2fa093aeb75555505a3a3e00c853d1d22a765568dbbd55513;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h274a60fcdd63f29e1ab58f07569a49ca6ab24eae227caf2ac24868bf5a143afefd582c6f1984412b088bdba6e404ffeb79f68a0c33423769f074e20fc1a5a2850afa4102487db55e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h834d268b4b27c88e553f4a884197a3a6d2ba8dcd16741f15418c07cba8f0187ab582e0135fe18e096d8faee9c7e54b14d1551f5eab73b25e90918f10086d12d04c5084443442cbd4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf13180c500865e57b38d357b1c6a121546d3f62ca86860096cc634a8d6a8fe66a0a2f6d439dcbc6d7e36c3a34582f0d6bd3be22f5cdbc83a92d7da6f83813ca6e0df20a4679ab61c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1271934d9d94cf36aad171ece35dffcd11c704c1f4ef7ebca9e1e2d72a369211e479b1353bed81f69e511c83d8a267e7c16bff3ccde49355ceb3fece85220f2971e74e40ec3af50;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf00eb7fee7ec9e3de9b2ea470b8b70e5604c33e7588651477d7984742a93acd5d1958fc3453f1a6767f859f7c0fd3a83f01dc4640ea3466bd2ba5fdb5a821d7369e8d9146fb742f6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e2595a855c22d289433c0eebaf8719c667cb2f12f0c69120bf6aafcd2fe7b9f1b95d9c6cb0a3a19d2e1b8a16b5c70abd4d2ae32db283ecdf15558b7e913a550ff996b92365c958d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h475a9d4d093d5e0efff55fd7cd36a504c4cfa8656a9dbba11caa2e0dbd504e89cdaa6d781cef0113d3ddd92fb26598773bcf98b0acf9cc033cacf5cc7d455959a904ad6ebe98be85;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h756593b1d7f6762513ee268bb14889f0363448d42f758176287f46706dd3264bfccd8dbb9189e1d504f73c13e7534f25d3132139eafd994d0000b6761b85895c25b9ea638f9a68e8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a1ccd235b6aca0e61438c6d817e0c46f077a5a1531ea50bdb7bf24960bb9e929539a84606c87d8501296a1f17395455e033a681783f8c10297f50e60b03481880b6b85f5cecb81c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9354aca41cd171868be762c6c4b2c2e00188bd5fb28165162f76b313e079a9e0cc8b5ab9a3511150e07fd605ff409a4f4effa7aae1e11ab953ca348d5d2c9cddaf41f4deadf6f6a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e04748583aebb6aa63ced9a2ee0e82bff3e0c4d17548cc8bbf0f41dcdb45a4e01e1fd1d842895b2c2fc9bbac00f5d59423fd42e6fc6c6df23ae9e512d5e9c3625900a096fdf722a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a37df9b473b1bfc31509b77a38de45221b3b48e5ad6a502c81378357afc9401320fb57517fe4ed20100dc04d72be142415ec7f39ae79f05e6f537d44640f7c0fc0cb5183dfc5187;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he55a4db032cde28fc01bfa2e38e0684bc222791a6693924ec71ff5d2cbb70dc6d28138d297b6b722df06c5952419c93f59dae2b424b74874b392c6e42dfe114e6ee933d2be04ec6c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd2cbfbb59c9560b5c2b641fec0499d2aa47078c2698872c2dc6c4000199f6afcf5c29b2ca10b9f6573d0093877d1277da0adc3ca85e0766766d4305bb4869204e3ece4b319d4bf7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58f9863764b5120d14e496898143dba08bb63c69c90a6f07ac20c4d99c5fab219c8ab63804734bd6e25ca27045642f1ab09f6f9c33f4f1ae4b1cd9d6bedfc76dd8e8dd62f5531746;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb36c333c026d9d0e56666e7695f12aeca18d2a366e395c2433f36fb494ac6674f90d6f3523ba6a8a8c918fcf2da1455afeabdcf67de4c2ef69ac702ca51fd5b1d6fb2bfa4dcefd2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6ce3b9a6ab665eb06a1f9d6f044ab0dbb0bd80f690e9109a10d4986dd24428c3c4746b92fa997d981941c0790a3d3c2a55126a1c2b572d334dd8dd789ad253047af28da44608a6ee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc66424c0a13bce0434b418aa99216cc14ee815ec97b3afeab46f5d149e8147adb7320046f1a14b97c300ed01eee1c8abd4beed8447ca1e5134ace1698e09ae84d7fd844c44702711;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e7cc197538a2cdaa1c365ac63fd74d958f538a44eec37228e38a80b8bb35fe8fac44082adf641e4377c32df719574f9bc8630c2bf8354b52bfc8c44f5370c71a37d5dd35a5d8ed7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he1408e6d0120d7370d3550e7523d810741dbeb46611d0dfda74ec51f03c336e8df45511ba05c564a620c427d9eb9a10faa41d765dc00b914d9cfab0e20c4601caa9d34c7e6d6a35;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48027f28a200a4348ae425423ad9f5ec5f86da37a962fa2835398a639af6e8677a88d018f5d172fd3505268a3107da0d81be62e4d6697e2ff4213d63b9e9ec6d770806ced57e6dea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e4c8f0923eb75cc21801ed9aed9d2fe4c64f46d0610ca13403e61c4bfeddff2785e97ecea6b881c2fed89ef0a96110ac5eee0050d23278bcdde0774acc97fb481d867001d5ee346;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e58a53d28ef4cff0c66a24d76350ab59048e11c1ebfc5e9794d07b564ac729565cc70f59c0298245ae5218ac7ab391522439420d268ba72d32a6157ef44bc62a4352233f2ce7b76;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h97ef890e18d1eb130e2993b3ff70cd0263a5369c9fb263fbe82cc3500e36595f8b3e7491630b6bd6a292425fafc6e79050edb877a71366407628997f0b0d88afe848b8b2ac43fcf7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e792df6aaac6f754ecdde91ab346bfda721da8c282938b39bd47f89c26802ef8ac4a7c89a53ed189d1f192a4e4b655c85a1e10db1720d59cd20430b94bb08d75ec599e003a30d2e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h620c59cb950e7595aab27da81999f9c3dd7c54ddb90383958ebd475dabd2ff4475a22dc8d35f5120d2e7077b18ecc82172b218f9139bba93e4daa2b018c18484867c9650506b8ab9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51fb06877dcfa9a125571ac55d6d16c35db305afb8b003bcc50d1f4639ca33bb150f7eb5aa75a05e3df2d65bfb77e8658fc2dc578e10c6c98c5bbf9de17c3d85fa095b4f4ad4cad5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87074f0c4189565c8654b55f72316c600b0af1add4ee4610dbbbb15f66467552a1307fce7d1dfc7c3db96f81d00fa7e5bae6993a86013e5b3e83982e4c1af91676fca75d1b83e44;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26a4b42a364452fb8d375f7cdd589296897a50b5588fb139e81aa92ae2d97c4276b5d33d592e45aa9e07b027f0775eee01402e69cb648771d12208334fd86f5888da052f3b5a642;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he83600dcd2601d659fc680d30eb5db9e5c41039f034f61dbeec1139700b5f18340476e91f02fd1080e5f2c5af6ed9ed33f6f8df95246a6a76326e7410369578ee4e2ec0ebba8932;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd4b01df5510173656230739ead52ab361f3cf6e2b1f4f816d192482e7418eba448c908a986a5ca82afb64afa6e9b8608715f9fc681f7d496592d35e5c99faf873728cd47fe00bc85;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b36a94d5ed20f1edd16c2bd55b9054b7f01de4c20b16ca43a1a46371795639fc4eac7abe5540a9489a6aa5131e8d9c7f56f480815f92ea3c64e897d87d90d4cb228c9a8669b881;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c50e49d8b2bb31b451aa1dccc5cc85429198d9bbe9cd059130ca095abf30ba77ff1eccb34bc5a4a578dbea5173bdd28dfc618d04043d835d6085459095c6805bb0bf4a91e520fea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d5412140e9a3a2b95cd8e2ab5f9f646427bc839f8b629da72600e5d738eebc114fb3ea043f2e23a8e345b935090dead105b9fb4f7ad19b6e1e617586347676f78a44458367eeb0a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h38b6ec64cf0b0190beac4047ec8bb18c3d0f411892a853e78a13945a219bee2cf6940a9d8b5e6cc3aac7d05081da36a7cd9aaa7d1db5f5557e809b644d1a15222b5578d3d83d3b1d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h46b1b39c4dbb5e0c782af0b5a8345ef06bcd359ce6a1f345dd07b6520cd94df931ad8c9300a96a0809f4616a683b8cfd4c0d9770685308092529ad80ad26c5f8072421606c414152;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ac5d8162d9d91d3e1dfd0b2c384121ed36669623ed9d86a607c4a2c97a448070709a1349371e8c89a52d63bf9566a975c152b9e187966286e81436e0987e4fb55d90f68219fb7d5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb3079bb747fbcc368def8c94a342fa8633047c43a5a8777aa8399af71b84af6421cca64b7984a1fceefd8624b5f093e3f9d6c26998d3a9b51012321434e466db77a50a34565e1e1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48bc56faac88edb64ef4d185ed3e2d44af7beff4de4644ef78130e89a82d3718b317ecbb65f7c13beefec6be5cfc5e58427c848a431a89c1e2af9a49785c111a63b8b0b7d362c9c6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3fd25cc0476bb5628328699b22fb40f523220c919438c2c3c1699035044fe3db590f09cd243cdf14fa040f13ae914e6b74cd6ed9e8c0843166d0e2c8ac21ec4f2475058f4f5ed104;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h22ad13bfc774e0aac66a314998a8d481ed0ac1e615446e820f1c16aebaf73fef1d9ac372e61a1cd28e02bc2a345a1a1cd07fdd9a13f8bada0a9edca074e67f59c2ad3ea7b4ad0386;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h532c47dfafb3791cfb9c7c8f60c9efc5896df1bd5a8d6270b1252e241c9a37ea544661eb93070560779775f237c28ebe87c0a5cfc5847a65fb779956eba84e4cabd36a04cb3819d7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heccb4a5cfed56cf3e279889caef6afbd76ad55178950cd9ee624c265bd2725141e7bee5deb700c2a9cf8d91f66a560cd9eb34689b3963c4cbde279152aefdceee5052f13738aa63a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74e77eed397e85c06c44c2c9a0fb4e44787fc88ad1674362376500c98a702fcd62fafdd68887c21b27e1dc87e7e5d00e0b12dca138381d5a2b3ee1f2c4e5f4ebbb2fb784680a85b6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6850bcbd67f1733809ab04d232c1ee5bdecd8354c52b2f0f6fcfc6bdcaa3b67e39055a93cc441a7ab4e87fea35fc7dcaa8d23fedc1ba9296a664f567a139e13d3b1ca67e47a89e81;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb2127ce7bc7c5fdcf2d6a15b15f77f971ffd02704946c01d762ee698c9e844730bdf67060f94f3f54aa3f552d6f4038199154eb71f5c33fd37f9b577113a0bf609a34b5f5656e6f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h931b53a525b8cd1dbc7aaccfb1a504d2a63c038ae3f8ab6e19306766a592004c9cd4711b0238720306fa1a29cbb384f1777bf27df6802d360d83f05cfe57fe2c2c45cd0cc2992827;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f58369e6f0f09de3bebdd6c91c900a6ec5cdc58676d5182ddb39db08fb6f06c2fdb09bb2ee2f04327044ba4bc339e8e1a2a383090e6eddb060cc0a98a06247283a41fe886e74c57;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b018f8c143e85ea86adeaa9398f877dd040993fc4b0220650c56841daa24314b649e655c08f3d416c0fcc3cd8c6d74ce6730da94266589eb11d9461fb07db9cd28209790189afb9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4714b38a9f1fc46110d573f0995f6c6b989a360b53e4d1ec732dbdf780ba3715be6eb62b18b17040453b1c1edfcd2a7737eb23029f8364cff26fc9020d349f41eed4c5adf5e3de36;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4daf83bdb4c3e9ad2525ebd84e38d387d42eba9e7484619810f3753f656ad553e112fdb503d2aae248c921fa6cfe5a24bd98d3a723360bc2b040010ac42c53ac3cafb912465bfd4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haae72285adeb21f31df703b2d8ba989fa51dcdd19d398ad1a779a1e1b31994d0e689573c7199a4510e7cbe520b818d00fa0ba6a9a2cdc9a6b96b2dbcafd0c7d797bf156a731790e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1bd332947cff339b7301e7ae20e6cbc1a23803e9467c2394cc1d1c2c545cddeb2b4b0f3b369fffa171123c50cbd9ff7953a4718fe0005d79e42ac99fba646d862fe8ff405268194;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca6c0094dab27b882a4923802e80555ee31e5c68f6fe7f1e05cf05d550bac92036a364e45f7409202ac59c44266391f8adf83a0422d259b2c60f59cd0809169c36f0eaef125489e8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb6505da67398305630c578e2b763ec2eb8932d11e38cad391cdc70f171afb3ca73db5e2dd1d536ebc5884d1a8c12cb334d6ab8cd1df679c11ba033b5df438859fb15f607abe3752;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94cc461293db0705df9105707c2c8210cfacc26e6bbc0d7cda429e4ac1e659c72e403e0c0b4a5e8960c6b6cd3a68561be6c9014ab9104c331b10e10acf931b01bacc5645442d9a13;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3485def920c7e856fc00c1fc7548c5508355abb77f8ac2c8ea1d3a2acc27083a73a338e5097ffbcaefa7f602408e4fae0e611f5a4c7be661ea2e0cd1f0e0fbd80a70ff368d2bb85d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ed02404c46f3fd2710e021ef3843f698ae7c6ac144ad1cea039ee284a245b28d86c3d86c81cfe4212b52337f5a9064dd962985912417babe5c1f9f63c62235da7ef0232c4da1142;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h38ad92efdd7f6756ba2d871eec4991eae1eddd97f202446a2cf5bcf5e9e9b924e5df26dd9fb9991602ac3a7c87bec68a91c956edabd7d227c4e9a26d6c7b7330b7a894ae3333318e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h705c6a2612d5185b179d101354583767179284430d6166f9c01bf95247a8601f889cd3ceb4164b3720322aea9e1451476409d0336dfcb19f4169c1c337de265d0ca24031f1d01e89;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a998ebc108859dfef9ca1d9b0179c8f4777846195c355f567cebd52c0e13e9919aed4eec9c58682a5bbaed93717e9c278a9c610454c248e9087a77499fdb39eaa2cb0de873bf14e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he65e128bbf0195a4e2a380b9c3e00ce8d62f03c336517489104c64fab8b000e90b4549b537a8ed82021f4308ef65f48ff7cf251601cb22c88002a0a98f95410ab70111b5f1e689b9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc981c42ab91ec94827905c54285efd112a124a451122956e10e7f48728cab43ed7850aa6642bf86a99c692d2404ca288dfc6bfbdb599e11eb81304638492a9bcabf75074315f1eac;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h37531f70be276d8f48e136d6788bb89e761d96db4137084cfc229a3601f92a42be7a2340b4550210985d5b69d0086ca40ba6d5a4d21a87ebb372b7b87788d48ff390da8a7740879f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95689330e8f69bdd823e702ef53e2104349ac31cb17a2c8c77a400221136493495222a39a04b21d77abf9f2fed737f6ab02a8459424c3457e8e9874e78dd036a368775509bda23de;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0424bbd94431086c360e15c79d3bb9fe94060e8439ff9b687e519b35550c652af0b09b506b86b1abf7ee2de5f3b37637a22accd06aea9bcaf0346481acd216374e707701db7bb6e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e021ac4d066ca28c3dc4fa1e2a6f419a9b535647a6452557f06e35e8f3000e6d464ac9223c0a5227ed5d90dee7a70c54a1a3a1ce20a757b281f5642ec54d704ee5755a08fb2f800;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hefa7826cf451a18c9c66d0d540ce174539b1e2f3da04e1e4af659ad94f9fa50e2b129774489b366750a33bc832a437464da7ac99ff6c65670c35f460a95cbdffbcfd267faf1170e0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76a03525449411301246eb41949890a804c2556f939b85fce7dde0da9a794e07f94032bcd76a8760050ef1b18c1ac3286783b779254ecd887c47ee6ba6c40b18272b7f0d57c8ccd9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5177411e59d484b491fee9b2dc1012ed1a957cfec68184118521cf787cfcac5d6d57f17f194878fa128fadc0c2ddeb8d65edad8c0681ac03fc46a008ca3afeb1ac626676d382ad7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6438e389658511984a49d990c1b801a82ae7b2ed478aff80247e35a11a9090ee2aa50957a3071e4ebd3adce0ff8cfa59254174555be72db68eab7d07fde914a7af6ec6f81f21a638;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hac426a89d4aecfab67dce4fb85bcfb6f848534c5737b1aaaf7e24513f7886f63682abe30e36ab4eef6cd50ce2717d77dd714bda0ccc7be5d9b0985bac39100f47978bf27bfc01c56;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2dcc507d78cedeb288b0fb0cfefc7838432dfd441597064410c10c47002bc02ebcefb8a79529a3e9dbd96859e1ac3bb3851e911f3649c54419ec3f2e075b4b5c25dcd055fe00e97d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd5a0fb828286efd2463e17c08ecc85b782404e1a1cbdc8e7d27523dcf2c765fa7fad5c012f81b0e404091683aaf45ef27de8a053b91932a404a337e538c5a30c121a1fbe88eaa17b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa0148e7d80f14efafe6573b24cd5cda5264aa933096dd0ae0c63e5544d265f0cb07d5a2120e20178007a1ee6207b298e4f95413897e4da0b1f5091b1d70b40a3fb8a5d28f8f168;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h431a7377c7f7c697d204c1b164862331a02d85af0703327a53229c636a4e2840dcfeeba7199ca81d81fbfae3ad02168d648cda6d251a596205a3551a0f48b989d19904a4c0fa3da9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3dee5c4366d968dde255f9d41098956480cc1c5a57db39fd30743b1f5e16c6d961169c05846f86392c23a1fb0bf0f218c7def5bddd8d0d843986eb382323fa27d3b01c15a205508b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h10aa1afc008986b004c41d2ce8b0a6ba6d76495b5e057278a4ff5d81d6c589e1213c376de3d2e739eb87dfb5532433cbb995c66b6977c855fc24c676f836543b5563faf32a940648;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb374b1c6696c27f005c2e8d7aac313069d2c2156392ad3918ddc6f41e5fbc8c437e39fce5ae962e7c6a22e03b9515b449244f87cbd9b069362537b6812bc6b6063b59f68ad8f843f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f602c9141fa99f444d540c57297012d473ba421ad3fc8343c68f7ba62d507398bf01316f4fa254fd27ca3d769c5a9e54e07b41c676e23c30929be2eab13f65f5978e9a88f541420;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h15b3052b38402f608431e3ad6997505dc6f28df00d565880c9e842f08c0290263ca94c814ce3367ec3addef14223217fea6bba094c1cdf6290009e1132becdd479d5407266965444;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h868ada6aa90932774bd3f2bcbb5d1a2f8cef6c786823b934bcddc95a834394dcff94d683c84a6f0b7e42f7cefad1da0c6fa22ac496264704ec984d46b300d82316a2d7ec64cde9ee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd50328392fd4c833e584e694593f685afac138e61e2cb08029a81fb86bbada105abd3f1b0bf50bc6755110c346fc2e93546c1842c1b21ebaeb5c7ed7264e7f4310cf5f4ae6f1bcad;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61146e2672192f76348a591459a60267463c57f7599ff6322dcf3a4df842c84a24147cf24af02cdc387413f03a0544dd3d0fc55fba084fae35a3976d8c44703346dc642d994668e1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h638b54a61985bb0f0ed9954f92e656eefe6871d5d8c6faa61c7f7ee6fc287c755cd2503aed913d72fb63adb51f196312452677f23bd400862f35a60b29339938a490bb764d8905d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc479d1cbb353366e86a2c76ec25a7495b147a1e0a254f53ea56aa2e4147f0744ce7588d3bc12836cd2803bd6abd4cae01bc6900e3f39d1a64524cf388dfef76c4ed236ee3009263;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha9e4227d787cecd000accfdbd9696a84b9751ed07409cbd621155a30f26ab5953206f114b2ae81240d48d77d53df8fae6e10f016592c7b26e7af8eca2ff91e85784b27ecbc908673;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74ecd3e54a5efbe09ddce501eecd22c38c513d6cb2d0467a744cc5d18fa381aef5201bf2ff04c54f74a00cbfd3dc10732f0569dc2916a4ea0fd9a5ddd5370c72b6cb5b9d5dee03f8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6879546f7c241a97ff87622fb8bd17d3c49560a4dfde7c20dcf52b35a0bb7a70e0a83d207294eb078b1e7f5759a4493c10f5f7a858d56c3c2221f8148fa3650ebfcab5e79f224608;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61b57bc7b54ef96ad87924af138924f346acb460e0e923028742fe0381b4a91a39a6de88fdbb01ea25fb13abc380040d05f415bc5f1596c39cfe58a4a5a67030adf5052d9f1ccdeb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h188568ec10c760abbd7ce8a7f33832194ca56ca2286dfb7bb3f36ee2720da12546c56879cd9ebcff9069009fdce2381e629b7fb78fe6029d52f61b4cf00ebf998401e4bf1db7054b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57b52a5c328e763c17f231d2bf34e0c5e5d53afd4b1ce434f7624e27c37906299319498f357569d34ba753a976bf308ce73df11d36f1267d0950e6d3d902519882675749a8f69dd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53a11c221484b615f2f53e3414dc61be12c91406efaefaa60e3a5574964975429b35f3af083a4945b7b0a5095a6f0177c12c343580ed7d17e9a7c12f7ba36f7c33444ba4c2ee2fe4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1bc2fe7959dab3eab73ce9b4012a52c6dfb6a3ca235aa3acc6a4639009bf5f15207732fe67960cdd025d05d545b7417015b1b4e953fd228dcacd806107b87216b60a893bba6de362;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb64e3f83c6639e9c276be9890b63821874b7e03d356b0d8d5eb77fd8c5dafc5c8746ea91ffa4144b43590c2479abc97cadc97351849a604216dd70f91be6c9a6bb8335d05d0df5be;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h93e73043dcb3026b77a1d28b07594c653605a1fb74159382712b39d2790ab298625126055c2936f6763f130eb8af31217c62704b3be78cd9606ff7928f0990f9e9882f76ec38e7bd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcc17b5fc8669552103c12f052c54da4a5249dbf2bd688043c9e1360268e75aaeae965e07449e83635491aaf88274c40d72eb1206b7983303aa553633f93a25ccfd19a05607dea74f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4934412594f649dc3f8a386ff89818a0c344a19cbc6d7930e77cd9f12ec95f8ee15b6c2c08d1e69ed189b78d0254252644537b936477e996eb15cbff4f9d92aa3c0531b0b8c6598;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9897e0a102c0a674bf48545f7159d8182221c37c9a8d3443dbd72c8e344655ff0bfc27612735723e82de296801f2d092170d7a94a5d128e9be65a4f23b262dc6a629b0b87f90d8ae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc1df6332299a64c5e042bcc100e12f51473a94e44b27473f681eeae95065d79f2202134d3f1f821b4f16e9ba4eadc6838b2fc8b0551568888ddd36c8f468e733f7f662419537e5c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h49b17ee9b7711a118e6660ebc6d18ef6040b920aae4c307d1112eb954d7be2f0dbe28dafc7ad1d3a83d72fa801fb386abf9b868a65642d651d23cca5c87eed2a9d083ece194b03d3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85cecdcd2e8ca37388e69fa63fedead969557110609b5cc4685e6ada9132d2df64d0d605f31b8a4b11ac4472bfdcda77794882fe6f773988ae41e74a6883ced773db5f78cdc1ee8b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd4044a825c6352b4eee23423fa9db0e530fc864090d15dc68eadee2c36bef62a3134bc2398ec738e9e45d26689569725d2e6a652bd98962942f85bebeab0eb2d30de46fb3fdedec8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha843bfe311b929384d5248d143f4ec0df02b26e04a70f892d6350083c9ce807cc0104a19b25af0b62d8efc971c547dc935a988089bdc6a121c0bc8f47c34ed60b80b4cc93194e49d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40e953301b11336db856927e655300287137d060128c01660afe06ad4f7e3bec3accd5515273da32e31665d20082b82e2b2c2b72eccab192dde6450ec099b5d8fb20e37cd3e5b18e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ef6996017fd6099b88efad5be72c41f1a7371ff94a62ce689c2eee9137a83363b7b4b9e939084bdd72af9477f6bee5f43a9043b27ec535c0afe15827d755f9e1d7fe0ceec7cfb3b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa379248104db6291e2ce263115ea33aa6a990044adc8e659c6ef371ef46c831eb1d6d01b12376c54165696b7fe9809eeea9362032b464baaad95fc3409787b6fd69e72e26f31c39;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h830e4646ad8a23b6c755e325326baf3d66ef1455e7e73e725bdf4d9b3a92f5d290f270d636aa6d527378e46b9f769d879ede0f3e7fb8a13a4257839d253495d6414edec565f2794c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4591190fefe6d2c8cb5143e8b37e8c7b45ee3e72c6c7aa8833b6eb8b474dede75e92af31cbd2e4f8c1b76f22e11a8e868450a1577ae2ddbd4d2510affb3ad57e96c46ba1b465daca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h81689fb36dd85c630d40d9029c7a748b787c75725b1f6fb2db7017388389ca080bbd6f8192b294f9468657c91208ed16a08a3417781ea610f5f309ef25dd0e28676ac4fd2b520ecf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25892b9de4b66191fca3990e70037e91665798aa9ae717f02c9b57015f1fd1d0e5dc7e54d7919d5a72e2a1b4b56b6c09e0901023b33273aacb55075da81805d70710fc4a764de92a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfdba8948beb112fef3a003fc8712d416fe7dd57e373291a85bd3b23a9fd21c9525e6dc66c5071bfa7e264fbcf1b1ce5b54ca2fb3d5c9fdf7611ac5e9be6637d62085ef886956dc9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8d1047325d3079cdf9f41f35bce52270731a52f85a3444565ebacd88a9dc2eed27ffddd28deca12fae3fdb54f195f34c6d3b7b3bfdfc5739773b2c955680d20b58311be4cc7f4539;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc876b3f7a1a052980cb2fcc15617389648c469d0a6ea642ee5e617b6aa0775f50828023d9ae5dee67aa07bd0cadcdacfd5e6db9caab9ae2f208709b107b7a36828910f306a661207;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h51243c96443e096c805428db35630d5f4f0e221d3e7a7b1ccf6fe2decb729c19202c6b658d7fef0f433a567a5bfac1c13091189229ed412ffcf5a08dea89973b242456a9f14a2322;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h147f0fac36666964a0d7e17290967915cd8806c66e607c11898f95e3b2b86941460cf7e2fa078a897e25879ed038b346365c5e920cf452574cacf3afcbba21535720ebd07c0de8af;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbe66b493c1c9ec07fc92499ae29668da24ce7fec25aeecd4a07dac8d74956828e36516c4e11b10dbcac0a7f317e62996eff5358e349f0b4b8bc69d5c8fc4e88a0c8020fa4512f7b9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbdca532a6d171f1143705683d0b1c96c715ae6f8884f1d6a68815403accf58142bfd0d18512771f7dfe6c085bbe7fefdea305952e539886e7b65c078ccddd630ebffa239d837f886;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd96a6088b28046ed70e12ab27d1c325059640ff4efe4f3567cb410578e0d73fc7c4abb6402cf195c1d227bdba41a0da21fc2fbdb3e6e61dfacaa7a3ebc78f95bcdfea574462732b1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8779d0e71433078495966600c755eac0157680b479a99d7c9e48613f30879f14a61d4c1729d03b5832ba0e13fdca0570a089ce6959ce7e8c60d7556092521052d1332348f18a295f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd703b64dd8907c3a09a6a6510d24659b88d0167f3faeeca1c93cf5718341206b60427983d24b045ee35b2746c0c49b1502411797b1fc235728a10a374cc0044e0133f1492944ede8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73714c83cdcec39f040aa964e3eecb4dfe3ff7ce1d567ceebe7c6e4fbce53408782570912aed2af9faada0225863e4992cce7199ad74870db0f9d8c30da6a7fdd0706e2969ae7f42;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6bf1b6cf18d578b8856922d3d278248b0fc1ecf14df41f6bcbf6761cd96b576502d6986623fabb88de274d3002b1fba8ccc47c69c9fca53524dfd9ded55d55c1d1cd97b095f29222;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd54a1d055f9a3dc1c05ff5de23897706ec26d3e4dee5164fcd5dc183f2b9c7194eb9f08b3ad2a2c400ea3a8adaa31151587b8196e8c647f5e551dc19b3783d02fbaa50b31616ac1a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h70510caf0b6637d7ce6610d215fbdb0f8793b075f1adecb0ba231f2c796ea141126b53080148d42094fdc79ca5c3ae069c38b8432947615d522d91fba03b9345de9b280193f38c9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc112ebde22016f5716402be23be7eed2558e8481b8a6fa155bc6fe89ac9a5d0e6dffe98dd608e56168e529e5f6b3b225a84382f7c30573a5e576897e3620e2b5e6209f2c542683c0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h30e1af169b0394fd64611d49b3a98468fc5e6728d78968c45e1e15235d433cd3804c3bcbc89598c46621af95f8c8724db1282add1f50b707a9edcb66dab9607a8e1ea96bdc1f660;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9a84de932e3f9d9e98561060c40135c49d2e8afa6a76126eefc01a05c939b5d4f473e9b4d2334419413dd9178d39b7e89c33956e3ee160fc0a7f3fced02a9e358773eefad2cc10e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf8ae76a982ccf6ca3781d7c4d3916e05ef60cdab65447fb8928f93a93e92cd4fe6928b1c528dd532dc75be7a527611c2067691e9965880390eb600e94ee1310d9cb710ffb2a5781;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd65fd74fd78ce5d03e51d7480b27ef34136cec7d864df630f5ba1d997e7662077be0deafd772b4d97d3ee5ba64608f2e06bcaa60d72f4081b86aa5e5fc8733e3e89edd2ff89f090b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h717f3b47c27cd74c0be7f6a0d4332972624f679a8bc3ebefadee8a530cc1f7e83b3bb8a047ce978fab638d493a50839fcbc58b215b5995a3aeae987d42883036f0bdad784aadebe4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7ffaa3971b2edbb7105d46aed31c625a07fb53b160ef361b150b4b32d466017f85995fe999e47d756b0efb592396325b7874b44a4965be8c5583514ae88041ad47eaf148f73e85b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf09f1c27148cad3fced94edfd9af32c378297bca14ccf03ad7f77bf12551422525330b3f448b1c6c2252c149dd5df929f02ece14c8f03b4635f8eca1aca6531608cd7a4a14ca80a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0c7a678cb3a4441947ccd8bda20a84565585d9845c26d567c952f2d9543da8bb9025e2bb7e4f5f5deed574c28745835dc048e3d26091f839ed507d0ba3f427bea12b442eee728ef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a1a2d16e982886d20b6454afa1bf1d43358465aea4171d9b001ff242134cbceaafbc8a9186ccd8e34b64951dfce479acf3402af502be0b7d7db693fe76837fb47e15038e9c38c77;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d86cae41ebabdf533b87db0df9d6d67a1c1c88a0ca4e72fa097cbb2f204d056ac3c0efadb66cb1f93c329249ace209a82a07f2d277fe927ff22ef382ee8fb16cb57d9c2742ab3be;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h36275e5019fc54837098a22b116658f08f7d094ba8c95d6f090860d46d3c60b0c225dbe439d717e7596db82cb2cac338072c5ca904f5997c8fb39954c3f35c95f58d2b5e317b3226;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h247d180ec67935bf06082a5ee5aecd020e3951bcca44a3028846c5cb10a4eff655ced3ebdb9dfa9605d49c001e04541ecc3c1d4627295b81d2ba58872768df68ab971c79accdb26d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h178dd45532147ed1e71f8ef007c33c6e02c1c92712169a29e27c5e61d20280b5be0c261d8132f77938112c2c05e157f7d310dd5a6dae67b292c3980c9963ce3449e6ed85448aa4bc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e9aa4d79567660379fae76c9b0dd80befbc1f988fb85aa47e9206506cad251e1fb1ba380fa903ee3f3a499f90c4d08fe4858dc618c7f883c89f9b6d639131b0487226f8d6b5427b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h597885b2511490545947b852556d6ce8eee710603360b375730c67f7c3bd871048916c15bae85e1fe76a0e0a64d597e6cfaf81bb79d496d82e8ce4adbed467b9072eaa1877d2237;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8086fa9becb7a2c01b3967f319060549cadd6cbec9929c8b43b2de2aced6b161ce47b6564e3394070a0dfd312942bcbdabadf4c81d70c93a3fceb11b477f80816854845ecaf4c571;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h144497269b7c766a13a79253320337f4c37f43e6dc24a39b37ca6e6276295256f969072cb290c4423d0bf9a95a1565adbf6f98f85cab9b3adec7cba50f4fd0a00a8f1d66938cfcb2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h30426477f47f8de7e2a889db6a68e9bf25d4741b1af42b15513b0a99321fc0fc33e8d51b38c3ec75729259bf78381be9b45dc992e2a5989d6e2c020d98bc508745b4f3c1abe4fe76;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h884bef2e0ba032df0279a95e4133fa5420b8fba2a13aacaf28b5b1aaf7770c108e8857d08ace12dd8def2dfc39b34f1c9812a59fca314db7395b74d21f58935c44ec15ebabf74f3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c7b3e41fdfb6a8e5639e442ccbb3666183fae972c150faef352ae2fb215b97788092c966e315242f4ad9368b9c8f2a250576b43653ab4a68d4c7c2f2c2ac4caa6910e4e898f76f5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h962e88feb85fb9d1fe136dd3ec8bb861b4cc777096f8be79815f300a9edc892087d077ab216c11c2c429ff0a812730f69ea619336d405d25be5f664f54e5f2b72c1f65db8c3cd59f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7ea2c407b1e45e3b016d50706798fe61ef2ed0c26b5d724fb4896227ba735b85702f2b3424593c32c0a5bb11b1ad37abdace7a0428221737fa81cb25a44e8f57c0e5ce88612639f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb4e5a80e7add8323ad2d0b1a3eb77fdc543229e41428247b4ea5c6c52c2bcf5e868ef7d843ed655dbe268fb62c0e9f39b06393dc402dae11f6094836a92464525dde9beff1ec41bd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h64f535f8df3840970b3f5089cbae1650b2ced21c36faa4bc9ab0a42b93f8468427791757b05d57c498bee413dabb2b863bd87cdd3fd5984a98ff9e87dc5a7a3a566191f44ec360fe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69b0a8761a641cd954651fd5daa664e5091084840e00657cdd49c9b0087540b18a2045debd47047542117e8947a7077921ba17df94c2b489d3ee2db6a57cab4f16d88ac3339de31e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3be9ddcd5b0e09ebc11ec3ade72e545a18d3c175747d32c59ffeec5e6f0948bb55171745f0ae446aa32622c70eefbb72514151f3a1d3b421bfdb8561c168b997910ebda34bccc3e0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb17727c15753ff562318c9ed982a3ceb30f60df83e293d69ca99e7616663ad8711005690f6b5bc6cafc3e9c969f3784385207bb53770ad2bff39270c00d847f0ac1b1b9a6b480b07;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h557631b7430cfef3d7dc314cb743905daf829c24e7763b8aeec06b387a1b345a1bfcc5a62fb86f19daa46c7b8e9abf487117480399fded9b941724c336ff2dcd9da6ee17fd280dcc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3cce1b19af0a455268e7bdeb182cc1081196fb5402dd34d31ff9cc1494b5721d171daecd18ed4373a826b94d3a19e28a05d604011fd6f1b02db426246fcaa7aa26a7355111f5866;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14d738ae07ab0e5f0a6c386d18e85d76212f462711bdf4e024586636dcc03e7c845d32bef0db1bc116baceb5a6a74c45b7a2680d48264d9046165062bf42b473b24c913611b2b9d8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd27b513c4753eaaaf90479f0181a3ade160362000c13a4437064a178c6f812a5c820b5a8131d537d4a278558dfd617dee2eb2439e87de86769db2ea389b33560dbed5de50fa3220;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h828dfb14a0b13ebce00f0b38f2ebb1c1b082beadd463ac48464e42bd665d94e0cd97238176797de215dbaac02a088cd35137fd2722d3a92b6a04d7e6c4c8ef2fbe6be6a642b69281;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha43193e87ed0208bdd612142bab86452920a085cc0c066ecb3c19b305e2fcad28b30a2349ddf893678d7a092b9896867b97924be8f188298aeb521081881cb8a58a72290eb9d103e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6275c2116bd02f542ee6bbb9785a0541b6b9a8afe97146d82638186aea3864591d57e59fc1e8a30ddecbbce659ef3ccc57f645a13a0f647d4397ea6620b6626d6606fe1bdd3b1ba2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69355846d252f9574025ae1d1e6e1e6f7d67f262086cfebb2b13716cff8dbc5a2051806a07c6a9223ca4b033926925ed778a5a0079dcfc17423a10ac60817355f2538e2d27f3cf80;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h989985681b66cc03e895f4ba2f08fd7ed75a98f6b44abb262e897933ab26b8eceda4b9ae3b30454ccc28677facd32d517af037e754d48626031e783df65dee4c14bd983c6fb1e875;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h66a97ad1325139053e7e315ada8c7729e6d71c1fd457acdd5380533740b5ec950d4c87f74da71c04044831ccc0d44be04407e4257bbe30b07c0c99b785bdbfa9fc086045242aab01;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h972363bb9fc8852b502a44ed57836ef81c7a5d132ab9b13a0b753b6e8d9a79a5db21739ce7ec02d6d3af7c6e49624e8ee9e1e1f1f95052a1195f86b21d4c9068a454c26da01f1f3f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf18b4862091bce90d670e0ae03236bc7a6e5f0c75447c79303dcf953cc0e14c8075bb78ecc13e6cee50cde742b521e800a4e1ebbd782a4381d979c5156924142bdb43cdd27b1b530;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b461e417fa169fcae1902c1d03ce189a42b1293c12af546d44251f23e55cff198c846b4f62969b429a9eb8de3008ccdba182d4b79c2d5387308a2e5e452b59231cc7f7260272868;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf75c22c9ce3da08a630e9aa76879bdf461e718e912641f66ddfa67f847b15be2325f808a0c26c2807682dbb609364e4b5c804d070db505c89abcd172cf40e216bcc485cecf7a6684;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4aff54b97916ba303d31b4e29adf40bea8f5e2f22d4d40264647af2d0423f48af16ec178f6ec8f77e83a83995ba237dad27f00a185308ebb4f2c6bf37a4ce233d424f78ddad4e47d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a86f41501c584f670660ff5de41c1b45f9c0573ba4a42961bafb46375d57c4647326a41fd575417ea5f7a477666c41703c017e5e550d5ae25716d39ca5f1dcee38a03a006bdff80;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h274fe030803dc66f794db19432f07bec9af6df51ace2d4bec6d0b3525e6973bf372676f312929e6ab789eecface1c8e327f4eaf7ca9089a7e3861ea5beb2b57a46ea75aaaf9af303;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20b839a1639096ea17a3e1ed5d4563106a1ae5c56ce0d3e816616a302ecb95c0ed5bf275fef64ccd9889309fe3b070dca269f54c0534d6a4939f99dc5fa25b297903b6239795e0be;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c2229763d399ad0d955e3fde7cb06dc8dfdbb6c9f3b7f24906a8c1f838e7ed65d2e2281e20a25c8684e1682c549f863e4256c20bc924b70b0e1d3ea00eb26c85629793a19a93a9f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc545858f4fc52a9c546c9588a9bc85e5acb539c8d27a2ec3444a3144754e8f704fbfac9138fd42776f8048dfb331ac63f5b154fee97abde6285590f30ae0b727b6262a342be152a8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h379f85fc04790992397bae81650fe2a0f1eda7b059009aad2b39c006558f29dd12d460cbed3007721404215738eb16550217429265fa26732c697225267e1b22edb6ae0950215245;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3429bab9a60546256c94949726c68004a92df1e3aff808d4de02691ce632d84336415ab10ed3cbd1e5e89144bcd6c42cb3d4f6e3ac780cc24cccce6e672edb2b5047d554a20ceeff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e57062382a35bf6efec823cf8768af0f2a08d0ceea8397e2ecb4a3af38602fbe895d49b2209759b381d3fe975b959a1c5b2d7aa9b1c41cd17eef1f2f41531f576c9d5f663844f36;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf923287438797eb65fbac70cdc9d76e801cf8305656f71cedc0e7b1326b3d4103a1d27b2d4a5d60c823efe939d990984f7838055c57e5e3dbef5ac5586d6e7f1aba97ccfa7b952ea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfc9743cc3ac88845bc829c5131f73e08fbfcc5323428ce7fe092fb60163de9e3bcbfc31fc2eaf84fb5a3fae1e47e8575b806c2240eb287760a41148088e543df815c8d3bee1dc299;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h695fb3036d6d05ccd101b0a14178ca2e91290aead8ee32b32449682858b89d874c679dd25d79dba65b124ac36f6db5774512868428080f53b2fb366576cb1649e2399bfe9797f482;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ae6862034d0db4c270ba5c20bf2a69fce22484c1d07182e94829e0b0f274a16c78013ce62c3ef9d74409c267eb98ee397786d12bead287ce574c463e099fb6b13c7a368f2a08485;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h50eb33dce145f87dde5680a21cc4e9b0487fa4643e2b0d50e0f31af58dd6a36a8b51dbba7f7e74d5a318b681dd17e12e6c5b4cc7931a80f5c31c1616a9ae89ef66e13fcba8af01d7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfcc0c32302a6bbcaa057efabe3521249355ec8f0c43e7819ee2a330d0266aec94b20a9b5d563ae42240d48158c9486ca64e4781ee83361f5fe5bf7e1426ab0e21497ba22c0005ad8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3247f337e95cfa5d33d72873287eb2f38258ca4def3e19d853b4ba58c8adbf3860be7334234a33d9df47a4e8192a2a0acbb1e995e68a812a3ffbfa0d1f9c7059353ffed82f513690;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc3c0beb48ed368e5eafe6682d673d1669d498ae8d280a0333a2dbe54a7a6db9791995a684a5191eccf52d83b8954315ac7a75c5d3e7df039dd45fe42b3e66a3bfdae76466f7167de;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ba64d23f07634ececed3b9473a27efcbf2a208a02d190dbc916afccbf95773ac8434217e18a9705d84dde732f122269572c1f80735104e0e093df6f5b872d0e7b83fc0ab528753e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26c2990cc8704d840d7c5e3e7138fd9b070ce6e2a775ae967634bd12a9ea20296ddf29e4691736dde2b72a2c9ac044a73d09dcef65187c2c5217a40d5f4ec5ee2964d164a0e5c6ff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c0d4e8246e8db1c927243b28a66314241d19fa96ad7dd697977999d7019c35c57ef14eb01e6b51b35ab1c1278b66d1dbf60d433ac354d9a510e8c7694c2e3ee0879f7f572d07f1c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h31b5e66323b2e74dcd20cf049bb2cdcac5a5f41b9d38d25655d3cda245a62eabc91d0c25061d57dd5d145cbdc95a12917033ee95f388ebe11229ce65f48a3cc217d475c443b68036;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2389b9f33c562b5266fb7af153c8a74764f45b2bcc0b5e44cd921c7797ec09299193670e8a2db4cf8dcd0586c773bfb2a8adc144df10ed3afc594d287c2b4bd33c52acd41ce486b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8cbbec9d66e4056824262833d4a9c562408947282de89e567c08454de6059fe46069d113c184955b805fed9d11e9c46ab41748017a1d2663877b7322ef88b0546c024b39a21045a3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c0d0ad209ca7279392b79c4851f5179ce245442401067713cf70dcef20b6d3a2c77483c07d7826ced19e09f9361b587e9d1a1b916e59b8f8927f864cda92c13e19fac896b09aece;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf995e228e07b5150704a7822f1df03527ebfc753cc0b43215271f644f145b80449f9a25c03df7ab974a1291e9e0c24c28007f1c645fd01f19dee4be333f3d13b7c7229145993195;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb825748683f02faa7a22740313b46f750cee46de0edd1c1f5baf32565a7fb86b3742fea02788ba10dfc5688dd0acbd07cf5c79953edbe822af7838c63bad7d3412f1e53d401d91e1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h473ac37eba9b45cfa19205ee0adbd2a6b5a7c6da06c10b7fed60740f61f8b0659e85f17f668d6f831f047231146fff4672705df4be223718672c0f544e1c24ce1e84134a6d99ab4d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb36dbe84728c162e77fe8fef629d0c84862cea432e8e24030123ad4a069f37a5ad5385f148a3c48fbacb28728f66d24f3da21f2108e1e8aeb5d2e5ac91eeb457cc6b5801a5f0a6db;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a4f6a6e2c4da3d852d18e435728e6dedfb25d60f57c72a66fb034c47859b7f89008a490a3d234d2c5f24e72fbddadd2a2a3dfca3a16f329c9caeab2521bf576160ceaca5553c6c4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff342aa28942267ce0525b7a9a6c23e3679ebd436bf27280a01d4cb38bd0edb61e307a13aa04c4aeec117176fd5b482dec5f49801bafd05c54ff77564ee2be00a9cbae882376b476;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5a7eaf608f331f8ab031e5015e920d33cf0bafa96d1fbb2c09d76fd9208963a6cc61e6b53a910e7b4e2098e97a70c47b5e01c493b6cafb88aa2a4859b8256263836c60cf9638a016;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5216221db8909a70d7e3e055d2b90050f315dd06bcde5b6668b589a982ded4ba5f9734f775e180adbf11319a4ffc5cd8c829761decf39c923a9f56497114a7a969de0b6ad49664ee;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf346e4985895f2e9e5d6374fd96306aa47424e5bb3a20a6389ceda379f9bee1c1e953d3cd99179af475b3d5c2a8aefacbd2703bca8159600765e06eb7d41e581ad79a57c6e8641b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6759b69c767873251e38a345efd47f93474a4e42d406fbc3a22fac1b16665ac070114a4532da6e2a38e4a8d3c89104fc57c0cf53ac2fe36e5d71eac713271961d72f5bd13abc3eb1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7ab464d49ad946f7515158ec46cffd67efeb9ecc09c26c5d7b13872ad145d5842634cf77ad04e55aa881fba900dc1b8651d5ec9ec0308f9baf6cfa403b39be495d672d7349eebe28;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55308e569a95e3c5b53bcde426d2f1f9cc6a2c134a72ab4fe19977f2e35c232f9d0ff6dc3115b558d41112a977e8b41856ea866847d7da70fe40e15be0b6af031503e69c2195b771;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18ea20437a7e7e59152dec283896e8e2d4d093e0b1fac41c4d04c3fb8176aeecff12fb62887c61cf36f74755d905e65813467eca66aea9535ac738268a31c3e57ca55446dcc44a85;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a20b2496ea339172d24d8d1085ee6da8cd9db800d3974d9791dfc312b59ee390394a7f0c99fc1ff494275465ae2192d43ac456cdc73d9280f6ae78b5f31ee26d5d2d2f75e40938c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h10017ae35c21f315d50973f5373bb46594ea4092479ea4ae5e3a6323ae9a466ccdc8d212c5b159a1fb6b50e42cc5c2bad4c251100e9a66a8af83ba79c1aa191ba2a2c80c601ca815;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6a53237833d397bc070f24f234d114e666c5aac72dc131f0b02c0ec0dbcfdad2af834a02c176a9e7debff649587e9ad2ef1fa69cb1861f517c4015e0064b28785989294761566f74;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29e1fc6049bc268ce6129ef93e9b383d517c483b1189b26ccc1e615c2e604536ec287d984a1a1eb0079a7ed9997b24e94ab2fbf608694fcd58ba5320a809b31389049ce1ccce7028;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26128b44b45969bcaa3d63568d555606806dd5b7054f069f0199b6bbbbc3d4fbe43641d031954e495c1de6ea36273bb1825b40a4c912f153e5da9e16ca8d51077e5d141fcc1e1240;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h10154944b737074a15c306065b3d3af844e39d13edf3d01ab4cf38d29b7195dfdfed27ec5320bf685bb678ca7dfbf7287826145cde691b6b7ec221b6e2e7f583c0d3b4a21c5ffa68;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ea3f818286e6bf5251436d74996d04e5cb867c6d917b4d20e3b4d1135b52f6073d0d75305abbb187a23929f9d893727dd3c084e0959fca26d01eded7e3394657a55a67db57b263;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h707a5c4f27821f24a9856bb85948a24199b0a988a2e532979144d54777be7b86b8e84fcf792599e733b172be45671c7ac2b5f363acfb1d006c3e20e89b26247aff282d52f1a7b13f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h88d9044e1d57bc698df9e14b574f6e6a6e1cafa3dfe0ad1a5569e55b8dafd888fa33115bebe1e679ee49aba67041f1f6d2e9d8a0f41b633d38352e2c5efdd80b0c3ddfd436a3ddf4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d594a272d0145191c54607a9e6285774275ec95b628955942c6960801bf29c212ce7383c698962adebde7e5c6eda0a80bc6654a1ad89eecfe57345793e6b6af24e2b980ba9940a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h65764e829826548a30c6bb1e7ee84973e401ea6dedda1085a82090ba8c3c1e272b025ed0155054b7d0213c373087caed2fd7938b48322ce91cdba8d1febb5fb319c80c14765ff084;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd38f029312672416378c5f415fe1a18a97c508f9be26f94845c87fd2f0fef41c360e4875d705186a12ffa580e0d982d3d445ab987a03817a524305915ea95d1f871cb4fde0d50e77;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3926ca3812c9aec5cdb3e75a5b5363b1991defd8bb4abcb4942ed32d4c399677aabf0d9441e22c8658582789a0d6230cf3b0a5060a21aac1d89eec5c8e743781986ae5a3df424f7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9255b6bde30cb9fd8e08da33ba598f0c1e81c89bead5dd711f588ce7a0303497ba1d1e76b9fb4eec33f405e4e29aa4dab1339f44843d26bdb5733e4fe11ac6051031f03a2f3a882e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb504913b69771df03befa01372fcbc06a97892dc0c7aac4c797cffdacce58e2bc142d703d15bdd68d120cef43d48206384a92a64fe6283fa7b8e2d9e6f8632fd8ece3c5c7cb74f0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h725a7fccf2c66ef44c2c5e44f169271d63a4e0c3804ba54a9fc1ad36ef53512f4501ff3b851581a559a6193b9aeee44c17d2fcf8ade8682bfa4ee4be1d0e7fabd0c5f1f64a6b4979;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a46ff1fc4cc7993d802b876def140a8c531bba549e7783bc72f9a80ab9642798e872a2403b0989812bd520e61cb0f4928bc98f1f7c57ba61eb277068712d250d8d5090072788ef5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc66c6d38cdd882e1debcd76b7b12290c650160f54ad7c03bd72e924975b2c57de4496250f6050520cf09f3b5d41c7620f758658056c5d827b27c5a47deea81584041bc89c49c8a74;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf01bc41b9c5d342844ddc1360780cdbf627d7be6452019f5fdcf7614984ecf03c0fc589e6b25223512ec599f919d81ee6330218fe959ee18c422da82340d80d82dd1e0db9b8241f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcad82f8866d5f9e9ba4ec8bd8cccabc9c9ee6dbd356b978b1ccfea654bbf34c8b5661cfe4820bd100425e67ee6f7bcec971a00ca4253f307670e78962dfd193687dc66e9c3b85d56;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdea8afcfd4eeb1aaa7912d97892ad9d40467be77ace859c5c6fc910238274aa6d16ccd76a91f36da92dc4a79b03a2bd053d52a65d909675821f7ea9a6fd156c5ec682a223c361bc8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78aa59edec918f994e9bf94969fcd05dd308d5ac65411ec5f673b3a80707456101e57bc14f6eeca05c0b79a01acb897d0c2d4866eea0886cea106930a3ca612a70270925a61b0857;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd81e67134f18b1dfd3c39fd2c34ff09aa969ed5a5d47ba622baf9446093af3571af3ef77d3c76fb18bd13597a03168576c7de330ed08c3f60858a504c73dea07986d5be2b8c9ee6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48f1b84303a6b05b671e66e6968dcc92c923e6357db59f084b0da53f09575c831020d3a9e609bf124a05085ce5abad68ddb36132d5954c134d0653901683fcd1fdf0422e49b19018;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h218688c71d3640c9d5668e08f6a51e12406346e0e591b5dc88d1184a3fc05ff7838a4074ab58ad41b24981296084bfaae9f976fbee40c75e58717e318f8d3ad99cb8b14280d694b8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h815d101551afb700c3d827ef06ea550eba7a1333a15760eed13f48b0f69328044a6b7962c61e60f4fd0c9e68f1ac5df0a16ce602d8329ccdfb6d624ede991644ed270eeb135c447e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfcb8b89eaa1e1149ceaa35509f6d1375985ddb3da05029affd13a181aa48175b2af6ffbe0295edf43bcc8e4bed1f2a08dc4f22710fce6cb7555f431809c813c073c5aa4917a0c21b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h709c5208f1440b9195991ee9876e98b7c5b77c77e84d9fb34378c3d33178909a35ef9f5f916e24c30e3736ef1e01f0ba94b620d0e65279a51d2a09d1597f81d90aea8466b7f88baf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60000e597248f0f3a8b3a5ca1c6a9f2c2cf46c962b845e7d14edd4fab2643134fd9cc06e26fa8e37d096464657994c00a06806eb55b49d62a920c693d9f10c0890820b0751a497e1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h860c1f45a9c4b43d234688602c66989fe5341973ec7707982ee2ea6f3bec950c17514cb53eb94bbd2c2055a1eb7f7ad87297a939b529fecfe38ca61e79c74b03121bfa49d2bba2f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1947ad7d09be789c904e0e0c0d584ea8eaf27093edeae943cdaa8a35efc38d28d9ab9014b45b725eaf95eca5e41779b2bd331caae2ed7fee49021e4f8a2326435899dbf89bc56c3f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdbb9f4f8d25fceb4efe36813fde47d5abba4c73784787b472743059ca2d742c60fdf6ada648fa2e182fc5f89e640205adc24bfa1e2a22b781ec6272cab54f6b0b9bcb99e96b8a926;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94fca89515a2011d39717ed9453da24156d253b47eae789e5a64275346342499d3a30ba4094960b5281a60a81d184ffd973da1a1ea4b32e9d18e28ca89316f45b4dcfc54683f4c7e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1940c7193197376080636a08a721d39dac54db8cfc5ab4b5544079578d4e0303d076542fe3bf6592eb75db1092e27479e2937b8689872a918e49563109e61f83b51d2b7c467fb95;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h488b365d6e06dd8686157d9e1853b23a32a8572db7feee7f619d8213755bd319c43344ae03e953864219496beaf61ba2d6799210e0113d3dedc9ebe595ebb5d50af36dd2347359af;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h69b2d0bf0a4eed965214b5929bb7008cc8df414a98ba1d325a352d8f1ccb456cba5524bb6fb1bf73ca56db04433683c8c1d092886d8790aa39e76a76f9d9495fe84c116a4744dcd6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b114fd910bf27ba17a3f52e0e1e3e9b47d52b71dfe6dd8e6b6a3b78d66e480dc7c15b8b80f0710f35cbb545f47ca21dc00ce79136f8add6bc26096ed5813973b6b4937734c9d43f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc07ea3a7d7be298e2eb8a2b4380659a5a259c1dd3cd89561d19390116a35ef4173cac87c27f95b128f969364de843ce2ffaeb1089b15a607b7f41e38b8f92ff93e9a52fef557f72a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b2d0a2eb97f2d384d0f28191fb293e53fbe6c076596ecc02cde070caf6489f951ace5a4ac3a9f9a9520fc4ae7d3ec165ae32e8d4fedf7a41c66a044b47531afb78d4b1d3d8e4984;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcee5be5857af34294c1b910dd758bafe133533cfa50d7bc0525a5d82825dfb11c901573347828bfd073fdc65f9700de993631e1a510fc28d0f214c40300e725b8d5f933f00b17228;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4c4fc3b0a354e487e5f6f91f04a1286d8fd3f63edf0d27f9ef8e0228dfebe3e37f721a70ae1340dacf802c9d97b9cad20929e2b40354b679b41ac0a1331f8bcc4d47e0605cf9829;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha2b45ceed9a42e9a8f8649b6f45f541b266f9dfd030b534ad09962a4cb482eb46b2eb2ea78717eb688e4e0078c578ae634a2354e67ee99d0cd27ef65fd2b6f149197a18581ee1d5f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54224576872ff194265f8cf72a9471b38887d329135ff261de9c87a4e8a72c821e044e0450a85dc02a993a13658787af1575bec73bd915c3f620f2deca1f02a34ea9b137a9fac03f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5067c5aeaaf725e0e0315d2fb48d5bc92cba03b1450086588af9329dea82b8ade249432ce2fd8c2cec18a6fd67552fbb0ceb1867285ccd8621175fba6b981020208221a82bf6bae9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha066593414da925efa53353e3562ba0eaef9401dce6f0401519b62992be84a3fb8c8f4db3faca6bd0ca00e13ac0daa19a98b114811fe93dcbc2e8bde28e4ec9d490e004f7e250740;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha563747f91caf109dd3939bac99ad57eaffa115a8ba0fa908bcf314ff2f42b6fce1196bcc22f2ef73595c9d2a00eea58b4918ed49b18a41e72da8a4388c408e3ca9969e44eaf2d59;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec1577b0ef07798c6929032c084f3f91279cd9b87db1bb4d745bde984b5ae9c77487e7b3ca9c03a8fddd761e9f6f9543a7869d6a3109a472a1eeec9dee656ff6eca5455969b7fb9f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdcb2c7c54c8318c056f8ecf27794643acb4dafe6866f5f843eb27594675d8817e71b47f93bb0810d2feb16b296485d966d3be99fa99981c5e2d4e31bb2e5ee8b87b063ce12a46565;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a8826b028767daaccc055e19ab8fa5efb689272b3f1737ba79c0d8b231e7d528538e55618a0146c3ad2a57abc56220c073ec9e305468d104b076607bb119c2f5a9c43892a0a8a62;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h189d8cf8c04126b62078349788fe985e3c49014c3de4375ebfb6bd9c08ff1d911b7775f10fd64bc0e753f6cfaf4212e9db017277ca6d7fdb93708ccb2fba914b2f9ab7b6b633e9b6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3e0a06806f9d23c5e8b370876f4d5482bfdbf26cf358595d4c328566d4f73ece489605fd37a8f7e75658fddc677811a0d5424dbcb3689f9bf5f3ff4bece4e1e2d53ed0f7710cb13;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h695f90e9789a1b8118001138457606c8b8c86956e992547a50894b48b61beadbff84f0327b96a189c1e714cd2e3ffd6ef2919308293d97ca3a04b6d00eeaf1d0699fe85f772cc9a4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f841b3c364a387706d30a192391c68c454e55d66409383268eeff8b94879ab9b817d4834d3fed318fb1149c744fc262330432f6e96f8302b4b18c2b97cdacc101672e4a0978e763;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc28eb2688a7fae88f76640f3a88132c6b34df9fb8d25fe085dde1a4f88aa29a656a5285d8f5dc4369a4097680fb3c2300ed0bf0f4296a50d63883acd8b9497825a86fa695e3d5337;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f3496d9ab96113621df7ed6219a26e7716414eb4df7bce7fec92fd7e2a24bef2fed9b990dbdc6fa68c15a43f0ce41bd5cf6375a3888f3aa5d42e9127217f5436288da7ad39ec994;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7944ec465dbc74cbff4872d6c191cfb4ec248055894b155e8f5d8b2d69200dee76c2c35916df6b5cdfe4cf306c8a1e655fefbe40c55ba66fa0bef13738e1577e5e89565001830abe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha2bd0ce1720583231e08a9262eedfff409d4f86f5d27e164063a25cd89400f2c8d1fa054c42571b7b0f89b9f9556661763c508efad1ec5f30d18b74e18513c7263c3e646880159bf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1b36228df533154fbf0755318db82da7b8c48a6cd45b3a0945fa7c38b4d30210b95b15bb77fdd235bc0ccdabe97e42bec2490beea2a754a2b6337b99755b4254a120b817382f515;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb57047465c8175c13b43e7d542ce33bd792a9578d375fc677c0e56d604cdd89dd18240ef5d18f29f8b01f57b20ff0c0728b864876fd2613b5ef2760f7229ffdb7bcfdfdc859b0f5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h72974c57451faa438e0c247944c5c9a350560f2b528914b65deff7186943a7775c59dcd53b8f485a51147c584c7ad0f82560c41d58c06a2235e165eaf4523db1eb6cbf19b0ecdb70;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h600ace3591bfa2bc2b75e13a4421f1d5d82a45804dd7aabbf6110d325d5d2b2d935b701e9d7fc74b375edf66869484443a94673fb0242d2d1cd9d460e5dc41d367d698e558fb11e5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haef2782940d140f03f855bcc9a37f41eb338f0fd1004f02ec9438e5209045c46e1deee48dff14935c3e7ffde3f42a8d8c24fdec1c4526bf7e18fd6b87499825b00db5306270ba7e5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8e5cd05f958c65b30a48558c3e1449a7002e04d7cc89c58a854a6527a0c99997e1cddfe9d0a8360923fc6baeb0874341d692158c05b63d38e1ad3052c97a3f32d819fe568018a0d0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea281cd093a53da0872040b4f1e065fb3f4b78b2f18c02089d99f15a3cac8ce0900f8ebb9d710679b85c36e686a2e48f4e017ce47f2aa3496c4787f47aadb69465a56cfe88a3a6dd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f5146b1121d3088ef020c7d8da5d2f8c897fa3e308b4f4631908be462620329142ef7273dc5c3d00f36458a67549978e564153b702107871d0350e3ce1c9a91e99f4c691860e179;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56e4878c678bf57e663e77ad7931f93e76f79d366756e497c30b2b0fb41e6f71085ce662564ede79f8656cadfaf9fca2323a154c56d4dc87ea153fd13b8832881eea3f77364b7f41;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4abc7db6d736c62ae58e65ebc45fc108a21028a35a371d587f871bc9f98585ff732177faeded8d63308784c91e07740bcc136a0e9ca60367d03aa17db481311c0f14d51e1cdaa92;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e19953f0707bb6da0ef354360d99fb74af7a0f37222ee946f145d13dc4e9f30d1ca270bb720d2d7d010c8f5e52c07f4b93526704fbdd387e5a8135bc401136e18948d5241d41ba9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he5d95db24681b7295fb9c1948f7074d4659a2bf5344b901df05e5fb3409f5779ac601c11d73bf7eee860c953605ff936a7e7f7cc2383c70da05cdc77d1b32eb065313c6e1d793782;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63bd486909f78f42b3167cd3f1b37456b7f35648cc8a7ced6385a9d5bccbf0842e2b15d4b5442d0dbc210f57ffc31f065f8c9ee3746deecca8f8a9313522e6414a21a132461b831d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9dd25a264ed2536eb834289a9857ee88775e00867e401811d9987330999c7b24dc93472d08026adb1f33af257ae785e58accaa19e39b2c121c914a88247d5bc61231d2a55927fa7e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8978111fd2e34964319e41219364b250fc9636817eeedb99f3328b354ec3f9abe487349e989e4a4d1453498073727d028cd8c253612d2cf2d38f3d08fc29d030b153dd1e8fb2a1b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68507fd00105dd45fcccfe7695b92d53bc686ad5810cccd3d318c7f7ab01a845dd412d97433bbd96bf3808287909a8181f453f4a74e968843184eeded6468eef826fc89831a6f9ef;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h494880c52809987aff804426ec7940e4f569451eb812c5055ce811af41235a17f26ea68bced9d370f99239001b0aa0deaeaf784de22a3def8ad1f9c908db3e868aca39f253f13931;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf2a65bdda0b31ff73e64734b04152abc0b182d7c4714b93334ad42fbad45ac0f34d03ea1492172373a1ebbe1b5e842e4a17fb3b29fbee705316253b290e67c658374cf145aef12d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8eab79ae0f0eb487fef23fa3b945fcee8d3d1e8daf8e6ddc5f6645c251ffd32accead713e880084cc52ebdaeec7b291685cca52408d839cea40cd65527c235d0218cfc902383083;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ba44c5413d8f6e99b0703338f35b87134a2349db5dcf8c95029a6294b7f5b8894bd1e2b3a490aa7bf529fcc879817da082db1e8281c9b9b3e57f01ae9f74cc08083f62e4207e1f1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d07e6681671b4c9453011f47da317bdf7851a26748012d1fd6581cd26eb5bdeb7e62989f926ed26ace70fa8f0a0ea47528a2656e9a5804ec884d862a6c15202d859c2fb5b3fd238;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec25f20629dc73bb9655bcf4e65fe337a1ab20044d35ba7e2ea8bd755e2d91106d1f82dc5f0c2d2f10f14ebc04fe19bdd0144eba53837c18e27c9799700451b9540258f1a71406d5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb0a41a87e6621fd5d7224eabffe9d338fceb85ce97ba838e2ed7818761d0b98d4633b9122ee6a52dcd1fafe44d8b46ded0c177de6d0216cc445f4fe01cee87c6062f32b7974bfcc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd44b164557d2574067cfd011503b253a4161819f14df0c167f70e6fa9d94306cdcb4ff20857ab9127457437a2826f9d79f4440a922e63f711d7f2be3abfea084c60361005aefbea4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc66684dd6734f53d30130089642b48a2c011491262715683f6f42a8c38c8bacef9767cd10cd11bf80f6bf7c353bff29cccc74894febe2fc379f3ea4ad831d9e8038a569c44f7c009;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he511286d62707218bfbebe206f510992f6d2c3f0f68af43dc46916972223927b5ef63ab81c7c0ded0d505947016ffa7ae148af32ada0a33e3341c310d85e4693186ac2507141b7b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f2e186478bded2edfb2e3702dec76bb41a0c31f054fbb66f42f21baace681d13f0116d226aaf4372a2226023f04c100599974d1f64c17d9aeb0bfd95b6c520ac730dffd4773845f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76775838eab8af3f5c9e223a82063a3d29fe3d04931606524959c55924ea56d24d96b220da1f0cc6aa5bad066414b39f8d2e365c0f73a445c18dca2d33560f91b08f13926c4eba60;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde7b3c1252c9cf02a8ad579e4f87a98eb35e126a799b66b61aac675dc80a72843403fd92a15fc533f8f3d2144502632ccfbabdc47f952ba4eb522f20ab168d82f218fc32a24ad3c4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf92d6de50f3f40de0f24980ac823283572aa9817e83d82f67ac24f7b9be7ef9abb45a84ffe9a577813dd8bf605bc6a70d8305f87d9c31bbecca2e57e113e7175c407e48f591cc156;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hec119843253e28edaa331874eb0ce6b51a275b25de5011e02123efa80770937ed018ed86aa892a86bfc51564d3977cc08cc6001083c9af8b7dd183e241825fd3e53f9c857d920ef1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd9b5c776d5c4c522abedc37cee06ab2fbd97ca0e6971bb943663dab662e63c0b15dc9018c2a538d97e2898cbb291e17776090f4e2e0952e13e9efdf190e0a034b1380a873788978;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7f72445669f02646e1659200d88e3d7769ed2459c98e9bdf90088fd538e4bbd67734114bf38177ba0d9d3e6b2fa3e7609ac774d362352ddfe736acbd55504e8c9da0fb34c4210866;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0845f0a32b23b2393ad21eaacba64027962849a58f09028c98800e2c74d6c70b4a1162b22b34867c748b57b417bf79ed19c80a97ae97ccb676083a79b42237e189a6f483d676a95;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h14d6f7dc1376b1fdd7a4f844cfaa78116ecb0476a2285e9118185cd4a77d7da2746c4a046c537e132bb37bf625a234872db065dc7ec1c11b0e6c22c9c06d24f88d4ef5bf80a4a32d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79a8f45d38acedc4cf3d1ccf8cf33a6c13430e75ae7ffac1e1ea85cb4428e6ddcec4cf4c99b766fd4504066e4b66f92b17326ed65e1f4c83fabdaec19bc03456393b90a67fb46a0f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5af258e9af4087777fcf30c18329b6bad255db9bfcb6be6d23fc8c739e31b437c3e6b44dd1ab3cd80090fa7848017e2dc31af9de3025c7fb6cb7df1aacc5745924d0be79e538c3dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2677600fbfa2c91dfd72ee3cc57ae2a2d577e05f76bee20062d8fec0eb2471b678c2a02c6e1ba019412fe5544d9ff75502e75f651a3cabe220cab2238485c9b32646f4818f48c1d8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3aa13a4e246c4e69ff7028019fdbad69dffb375c6624a65e48ba15a2f72f2d2f9fd0ada6234107cee4b479b2c4e5f5247f94e0b68193f11c4543b7877eeae7bc233cc042e03654e3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0649591804e385e6f45054a26f40b82e3d4e16d167a201a2c11f76882c5f5a2b3adf1013dad5239a5a6a138a367f683168f6ac7b49b20f61603830bbbc1949f5f56f72cd47c5eb7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd75d1b84f26ce7a30f479e3e040e980fac94c499c030690c4f907cf37f883f2feb9d929f71e11cbd24c1ec9d9c188f83fbbb3ad79b9a613b52262ca1734f0bf5c3465c2e4e9766;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h128625ac18223194de9f0bd38ff486cdf26bdee9b38aad71b040f56cc0e032b9bf2476a8c7a1079cfab71d009d5406c025cde4c1b6f3ddd26cf7484417d29fd3d92d4405a403ab39;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h103fb5542a15886bee3e111fc59f45f1148666e3e9c291d94112e03ceb4c476a61be94c04747b55c1ff1a3ec7496629f91ae842eba9244c7a4d4f5a3b1190a778adb30e7e48b9e02;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf243d7c4c07973d46a001078d3e1bdd5e0d4bd12fac971887c89a0729d532f06211f3bfe32cfa52086dad36f43250b28cf5dbe30537f44044ef596b27c101fe88936c493a0aa33fc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9369542420b4d68e3e7e6cdad21a7b2687727f7c329175c5b2b8aa44edfeac9e7009db84c71af68d4fa0123b3dfc5b7f367db65c6be1fc33262761259e89ee79b4d39ee9aa503d85;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82a25040e4de596e3e472f2fb4b1166c10f672a4479ab9327ee75645e276899cd3461a64bc52ef731c2d935dd46b445d0def0bace4c8edac3eb8fa369b9bb2c9a38c1e4d7077b9ce;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1c5cba217b8c3e3fb67ee93adadf8ea7b5eead0011849b779982fe8394ecbe944a5018a1e73a552a0499d80a726881fdf34170d982d871547de9e1d65f370641d4bfb157734e2c8d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c21c9cd63e3caac40f700b909f305ef15b8e97b3f6ace748ead84cd2add06df1b008a354cbf11dab5305dd50034f2fa2b65577dca35e0be2bf4a420ee2295971c55bc245ec1a57;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hba0776efab3f6703b861c09eb7e519d6aea7962b1e45ddac6662f03f29b1c302ad263fe09ae30adb8b4d7fb49406f7dd1770bbd71fdded95099af86a718661218e080b342f7c7dd4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9ce415e5e26b92b24df7a267499d8eeae26c10ed24e7a97df2ec0a5981fd5b38680f2521c9af664878b33ed5df2574e478ad7634633bde26834af83bd7ddf3440afb2b827331b442;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha9df4d94e7fb63f0d9040fd161c6ceffbbdc1273c4d0e509516e1d9b6a5a9ecf3ca4b533f385b874cd1da9901ce1f7c39f890911bd69d5f96d1e1871c91b2066edd8337dba3c60bd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heff483fa99fb4bbadec03e5c154f0014a7542f57587f4031931292115a12b045aee34a8a93ac929488c26b234c1b583dc1838c20384b2e7f205d6ed84aaea8d58aee68ebc0a8378a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbfe31b701eda51a665f2627aee5308fe925fd596a688b610f59bc1a1dbb1a3427fca3c494669005ce4e11b18a63d0b06a36f83ad04edcc8d87547bbcc95f4fd47637f8118287af36;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb4b731e6dec7f8d4c2b1de2123a7b0de044ad825cecea97f279109fdb1abafec172019b619207f7f2c3cc11ee0a742b6ef4cee15f32b3fbb88ccfc9422d7724ff72b67ec7c21aa0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8d993dddc3e9811f8aeb9d11c8f580d541e7b2807ceecfe20ac66b5608db59b1097d84582fe962583b31d07ace295ac13f92cd7f07284361b14b41f1306ec4ae67d8c08671405625;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfae0fbb22ce4c804c0b89e4a1a89539c72903e933cfe90ea5f448c08f245e045e3c1343f13fa0449057cf433495f2cdc75b4807b312a3bbfa0016a51be0ebf9080c6880d7bd4ce7b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f88115c3e9862c97fee262310dde838b6bbb6c0e0927c531f8a88e03352944c7424251761e18916aea132595acfa10b4a44ca33c39fbae185089bf72eb1e95cd72d0eb5f7d0671a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf30455f5851461b1f9804a7ea8a61c7ddcbc5e7f9939c4987f694418cfd98d64c3ee3555cb13c7a7652b5df7541cc5e7f839b28ebb0fe4c27a1eaa49c019b4074ca8550feeb35a57;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h62c1a6b9921ae1f032011cb44006570e26282f847a57523d4cf14bd9bf86d59a5da353aeaba8a2bd4227cc88fbf5f510cb43a78fa9a966b70d80caeb06468d8da01d3d59f196a577;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c3948175e19486437bb47c96ae3f3ec2844bc10bd1c60a2ac69544ba508d1aeb4f7ed80564988997878661251f4f7bb22ee3d97d238724f26861cd9fcc3b9364ab3c8d2115d703a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5716439f25368915b4f8a3b37c3a37330f08d5d22689385e3311aa87e8d21eb60795edda3c01a502f17053a33fcb31a21db1e762b48a5f78f083836db98d594629766272fcfb5452;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4832f6d27b292e58e46303b31f94d8a76eb4aa3524c5eced9693509d6de62cd03fe168a40e0bb09dc2daf5d97579cc20ceb1826668288d3f3877c3cb444da4cd40f2f998b276b44;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h63dbab76b8434f7396e69b986ca4b0cc9a9ae6c79f2c61b180122d3790d8b17b5023852bcd611f2d1be7b466f0833cfbfa9d8b47c7c4becb6e621da22604aeabcba841d591af1128;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11d6b3124e6434f6c716c08ccbff847a0e3b8de1a7023bb0b7c5883a6b1274a154a1a3e5b32572ca284d7dcba4318957dbadfb9a0f28eb92ae0a34b909bdf97a21e5cd1a0e082c12;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heee15fa04cb132e4bfc178e6d5cc6c6ba3764719d8b3d7b29f2045238c8ab8cae7cdca5242dcb9ff4a811b39a8ce9c63a5e996f8c324afe653b7604532434e16b87d5f4de0d9e132;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce5c3278b5e2823a3559cca6210194e9a873b8657c6633483fab4215cb6f80e48c5d9f55658fd6053d889f8a93663d38d55d835312fc1dd26665279a3dbd21265ed5e8abe7d80fcb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hce4a9521432a0d7ac776835b9e1b2d84a090f5cb22db3809486e92f0557e69d9eba876ea8f0bfe4573fea95f5a2c1e671c4c20ed653ae85061d2a52ded385c7087f4a536ff55ec95;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha0fb6893016134529e1c294f97aa98cacb5b3f5000026233cf0588f87743d48722fcda4b6203c67679ac2651e9ea33094b831ace52717f2d711e2393a4a3f37d33ade56043cb5fec;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff40730d81910f37367941d79fc253324eadc7a9903375bd6789b565e6767c7b28030b83373b948e64f568ab6af522653073a670362effc287c27b0c73e91172706386fd2733229f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3228460f9ceafc7c6ff3c9c92461b1af17d44739eb7a55fd6d8c6564d6f5c5c02db49936b9275bb4cd2c8f96a1d625e20d40866f9fed9102f39ea8cd4f10e3a7cade1ba58135e06;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e2c921c47eb22af68dd3689ce7dbfb6f529de68e784c74a3b0907aef62fdb09968c50155039be0efda7709d9a556a1cdde6365d777a74e447ccb3fb4ec981dbcfce2404d6db22bd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h29cff33b9ab0b92e63d3f1be686a33842f64a75cb054fb6785e0b13ce1a5000de8ffa9a4ac3045e1b757c654c27c325fba975898e2dbf0b9bc5c08e1fc4e44f9b52f97b6499027e4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48fb4d619d34e8fa1eb48f82e7dae65b0729dc6af34240d2128e8bafeca183c85eb2736fee5fa1badfb184bd67f67079ebf4d99bd68e40b0d63066c1eeddeb368b849158809c4031;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd3bc43af8ef8b7842bd7da016e9aa07d4f10eedc9eed89f2935d2a0d631e1d2f5fb1d4aef67279657562f805b6bd07d54a2025acfd3f9721e4a10bafce09a1e98f34352c1750108;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbfa68792070933b471cb389377328348642eb8c30ba15fc6922d4bf513781e2d3cea765f7ac840ed598c5d79ca2bbfa26a52fdbd3a1ae2d5e8eacfd487b47fb8b0b0c48657ab04a7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7dae03e3faa454b80849ad327bc8811414f15e9f80090d2522286396eec9094fd4ac0bf6eb907879290bbd84c39796d3cfa0d16d188c4f36fd4119c697b18acc7e1affb42bc08d0b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1e1587c1e5ae85a3aaa46a7c59da1f7d5783eb3fa07f8735be81c2517019acfaa4bec01b1f2aadf2d0532c0d15dd1a4bf2de72df147c5ad04d106d757a703bbefbedafd9c12289c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h200d2ad2ea9a960d1bcf1996161cd36d540439baf60c2d5c7e60af525f0974d9763dd3546169f09e9ab12ba49910597aaa22c37352b114653a90dfd907da83bf92eecf277f509009;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e4c1f1fa0d48dc184f049618c757a99c0be71e4038e4cadf632215ab651297ed88e568625f4d4b27b5001966d1e40708e20ae7ec0fbb84326cd062a5ff8db38c2b1ee3328ba569e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfba9e70e92745ac1a0d5e68d2df7d86d324ba6aadf6b853ef0b372e2713b76b71e9e09c038eab4ce5f0ea17e930c40e3eff3be9cfb600e20b48297f2e0bb166ef63c23ad5a8ad7de;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h84cb22e947561c6f1103f7059694d0107ae04bd157c080d2b9a4fbe4d87219c366f2b3cd0f54814b83ec61fbf352eaf79e33f20d30972e9a85f3b8b8add7edbfcbebd4b45e37d4e4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf28512e3a215484fc75c21fb672162650c68069eb3976ef9fa39b9260c3991e2f788ff9beb876cfa493b2d97814226800b99ed3f529058063448660deda8bc4697c62e2b80dc67e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfef05c7714af30800b6670d3a9ae0874b386b2d2ae9940f925dcf173c51aa384afa5df0ce72832bf7bf031623b3787d9eb71bb322084d47c6ba3e05a5c4845da9d6f1572bda686a7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3e961603baa607d0613d23c79253ee8fc73f66954987e37ecbb38b6a9a264ce4b121c8b943b0ca3ad9f18a0c148b98e47f23f449492d926ec40a10295d010fff640cf64803868d29;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7cc532b0b34585b0cc19629e93de59f84f484796f31942eb651a46856720457869efe48b2860a76e186836525edaccc8d7d5fe4acfdec30a79a25b8b82de9bcaf8d314a6a220edd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h244050a5882c8fa428ee6581cc84a95bbb2c28e8edd2c61000910a5f35cbcb26a0f1d0a2188a5408a9dc585c01e951b092f8385d96f8c8c7607473206f3a40dd9cae92aecc44df91;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha19d29b9138a6356be1262502f861e45abe34ce22ae832b0dde625d5d5a838fb294e004037f89917fd468781d44028c35edbfdbafe17d17df07e9dcab6a799026d6963507c1c5012;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53bcbc3d976b45209f7b2e4ab2144517f6c25b916be7b05b5bc28126eca22d59005b2b7cd36a583d0e83084b7b6e831bca257eca65399183a7fb03adb165d7c4c78c448536c8e33a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h71bbe04e29200987dfa775459e83874d74540cf97d34df7c774ce8b9fa55b8b566017cffde9c3e7c349918cf6745f42320c0e8e7cb543b7ca3d6f12684b1986b29fdae23a42ef614;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdf102d76d81e4fc0df3761cbd36e6191abedc4686efa576bac6e775653beb3dd05e0fd00570625b5178f3b9919b58111a37e4689689694a87f6840ae4136b31ef7b14e9297643c5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57ea512059db7b2342c462e58e6af44de9e61ee84021e5665f3f74b6517eec13ca297e876dc8ff6f04416ca46fd5f06ed204d7fb789ebbb4789da5de198a36e8800997202906034c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h698f6c9cd0e61359fc48e46a6c294d06e7dcbad03de4fc41900ed89fdc3f2e15055fa2ecca909eff45ef97e268a838f8ce07bba112114b09d27bea82716b7ae1329f99052e506528;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca3dca9655f6bd35bae69d113cd510de970d51cd6a43bf3409902e43aa1505da3286676b64042df7be20228a721518226cbba6556830ca524f1fccc1c506561895b0e502ecc9317a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4245cb157ccbe7806ecd0949c7e516c18b95826c4896bcddfd83a2fad31bf636ae2dff5fc71683e2e4571b48ba4f7955fb1d6f0421378c55972599a95a978ca76d30088b29533297;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h548a28748f9311c235c8454dc2b2e04ab550e374e02e05da2f700ab0466db8c53bd00a819ca46516c1366ab4e95f8eb3c90f47cbb575d0828da1d223d22a233c8639ecda763ae2e6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9081b3c63cb9b184fbf31cf1506edf4b6181d746af22886e16a73f65319661b5eb6b43ccb4c898a576d06947ec6780a0565e0233fa69888f44d0182bfee7bd3806df54f5819da3b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f6eadab7dae38955a8ad174d1a16e7139294111b203d1a65062b3795713c5c22cbc3f4295e31c4ffaa1f1478b948aede51ac8610a2d6ddbe62ee628c37dc9b7bf23bda8ff51eced;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ec191da218397040e29b341a77a96ece14d90fd5afdbc405772061a4ebd0579dd16c6a4032d469af81724645032e6d383dd0a106614650ddd56cd354f823832960ea5a8c276875a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f38bf7d57fc335d13f5c9be43728e4acfce6d643fa1dda09d11b3629fc17c0ab00c3c13da997fe434e204593383fbf8a7573179ba53bcac5810cf7ef618ad473f54d5c5ae175ae0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd125dcad1b8afa84b30e0afe5998da29dca590350c7aa61bf4d04639a2b8e59484cc3d4a1d4640d6c12960fd2e71ad840bd180eb326b027769edc2c72831bc38318512e427d0f44;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6dc64725d1eabce169a5c99802f65ba2d49ec5e728a74f9a94804b1bb3959b1262dfd32df2e62449b2ee4ed2e05bf52ed3b9748a6364ea2cb5df6d890aefa9d937fcee4f38b40805;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h84b5a0e8441ee5d2c7480d75171da47515d5d6f18afdbc1d31ab58f6974524927804cc9f48e4cb636ba2174d8e367641a6346c4b2504ea36b144a3daff03c8592a063666be5855a5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf9f6d3ddbc0ee672cee03675f5b33a6c3c77f3baeec704b5adce5c272aabf11c0136c87ac58bd81eda55b44ceeae2d85dc1bba8a6da866fd738cd0f1a855912563a1f6a6a3ecd047;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h259bbdea8db6f84c4a108d71a170837227512bdc572789fef26f3afa748262ecd8f445ccbdf5547fbcb1fbf2b66bd7f605531c821240db1268f9a26782b8f158cbdb7355265d965b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c4741042ad91862310e9d508bc5bee2ff436ae6f0d205af9b1275a18e239cbc0a1dd27808263adbaac4dc434d17dbfc3ecc14e0319d02d098a002ed49c779196b8073c098fa6dea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h397f274982c9981abbec34d09f99b8ca0b26f1e45fdc3ba4ff90052165e13bbf66c62dd8b39b44874a8e16e3bddb450c8fec896344b2235f58ccc63441adc64a54ea0c0dfbae476b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h508ebef7c7b7a44ef58eb037fb6d98424589b0ddd913541ab8dd208fcec3eee22c34d8e88b670a3b0603b3b2ed13a4d9b852706eff25d0a8b5444283e93306fe7763bfb1340dd082;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1410781e960494010435154485f0caef86d2735221d245f4105d68782aca0e69ac12830ef6455cb7f07ed6780e75177305374f10feab42c549996622076389cefb7fda76612e5eb6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h16145401a6e2d795a0307d473915a5288fd76ee4f46f11f49a874a36fba74fa992f6b6a16082bf632445f420637d5e7475d0efdc685a78a89164be6ea78054fe29895acdde844f63;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6f581729028b806ccb505a565da790f4de0f8a1487be99b09d259c04cd25b6cbd81bbb12780f5f732f3a2882a04e9e1cc6f32ca75fb45f59af5e12717ff18513319d720c9c85c10e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd57cb136252fdb24ba8e077f92843449c741545250a1934b2732c36db0871713f064309b3c96d8ce5f6653491a70de3ba5cdec320739596398bd42434a2a9003103b8b55b84ada6a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h784ed4e026985e6dd02c5be4e8b72a57ca1be37bb4d19ac6319bf415ed7dbfd12e72124d5a3510abd11bb662501b74d893a22f3744cba79675653dc160bc8068b80c9c3c9c04c11c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf275fc0fcce4dc2c8423896ba6751daa80b373264948c4e7b9d0608ead6009f552fec8a8fe7fe68f443fc63eb15f208bc431d208edd308f727546f6826640298340433e1f62e5ccf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h61dc13f0ddc7c0714ff9869584193b024f383b438494be1750348c8fb299f8842afb23d1909ad89edb99ed7e49f9be425431ecc441c0170f592519f7cb131fa8864c7909d84be6da;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c011350b95db1403297c4af391ec88c93200781630f82ad461c30f1222cb9b1bbd3d92decdc11f6c18edb124d1aa540f219af13d4d34a26a0596ece1131d412c5b47dc0c37982e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d0eb685122edbff446f06f4d3153e66f4ea53d91e5876e4bb08969506c5530d4a53b5e5ee3362b82b858133c609d9530495abe4ac24e39d7aa95a51d412d50ac7c4e0bf69c13d28;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h11e27ce7eedb36f3d32bba636538c5e8860ae4e2fbf6210f23d6d486429d9fa63991e018f608ea0ce001163987858997b0f4b91423cbdb52daed28dadbee229572c7f8a9091e399c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8d470837d6f9dd80e963501d05452c7b17e484212f81b5371c16a7643bde9f94509e186b97c10eb93bda52d727e17bbd12cbfdeadaae0559f82e1274a24086a76058067ba1744350;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8ec31b8686962b02cef014eec2e9d5c40926f49dcf9a57e4c37ea7645c2ee8c1be1e7c2efd9bcf35a7df73bfb3d67cfd6ebbd22dfb73c4c2fe93289eb795da57d523798f4816525;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h49fab422daf016bdbb9b934af81e669ec51d4867d4fd19e54cd9a8aa26cb86c9e3d95510bd8ab4ed73caca2448c149e35783d6ba8e4b981d00e1c3e6ec89923e90b242aa91afbdff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42cd67a1287a956a8384941fdc5102aceb7e42f64cb52e9f2e6d4c4cf715a2249835853c84117545985e88e5a9fb318c2ab28d56822ef13a9c885329a5a43843fdef3d6cd06675a6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa95e26b7c9cda046c19e79669ec005e4ab8c7d7bd25111f123dfad9b3984a0701b453ef7af4a7ef940e72414553320bb16c3f0764714ef7c52a929e5d851a19be13a8b9999fb4c9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha36f1a5fe6ae804774ccb5a7bf1ec550f1f9fff8e3d98a2cc33b54d77e6088d47cf987ccd44a129f41a0d5e618574c214019d54c24c6eff50f657689487cdba216f988bb3d0ae8b1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc8c0a2e791208237bd55011b4ac93ddbb2ca8b26876309161d0763998e2cbf9dc0161e90bf8e3d30782172dd7eb8e388af15d8aca8f9ee9f2c8fcfc9d47c457e99d2cffe1f1117a8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h91e5cf3b9bef1b88069e08d7f551ebc8c4119cb5ace009498b21374e8a6fe73ad5a3671989ed9de1f0e8ba30936b22aea706ba4961e3e60561a4007ce369efd6b34415f948101192;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he413323d6c1ab1909ddf606798ff54fe795c5d72cbfb3c96dfedb7424080d9fd22ee13a41ccfbe246fa77ab7b574ebd8680ba2a5a83d649c8fbe0b0f53927a473b844b8f9cd9d518;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h376453aea52458e4c6b248fc64d4455d60517b97379a14736dfff77ad5520ec39c674df21cdceb04e486437a3699b15909428e205c0d3e2b5566987d0ba3c077bfc833d886b39cad;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h60a689ca478dae367ec771c308578d98512b82a86e906a7329526485535329855142329aa1ad86348cb67d5658143525f7b45e82febbdad6d3bb90258b68393eb6e8a7e0a5d25890;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e2008594d9123c405e7d6bf5cf88344808954ac9de5dada0a3800ce8c939f25d707d26ceb403becb1dd8593d2173fd26bb3109998223f4e126a61e25f6c1053171d8a7820183787;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf1504d440f1cd0173fcd0c32374391232d70a083ec62bc4d19881c2864c1d5255e7ad846d1632c78ab16cca54e754e9cdcad6be3a08ff1bcf5a647b13e844cbe4abe0fec6e4fdf6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5cbe556a484572e938632525d8509d567ea9fcf0d3c16afb0cce7ad6a4e793f42bc2a20abc061e76cca29cc25a3e4a2b23e336b1aa78e95acc0124b87d7653d5fbafe6263fee5641;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h137778ab9aa096133943c0bb77ea157c3994bca6cd4e6f443edbd75735e48f751ba8ea619e64bdef60efb4ff2a52a1e01f9e9d56c1218e418ccdb867d92a9740de1c89be2d447c27;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd0926407292e9a73f8b4c40bdca07dca098a37865e80398e4a32ef9deaeb03b17d2873709836d4408ac499b47df2b94e8530f13e460dc7373b93c79830e3d1d91eabf0f069fdd7d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd24b4f14adad96704c8e68ffa5c36fac2043eda9f63b39d5603c6adc5f1eb6235d869410bda6dabd10bec359cad4d72696e5db78047283a1c6ef181c0d1f72cf6e465343dd4b11db;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h82196fc7e9c4440b31de1db1f5ceba6428f58b3f9733d42cbec1c30d89d2ad4d204573c1b3e6765aa8da382331b5e17ec18704544174613d1e1e7af3cf95006d2b6cac679b24da9c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ebbfb57c4588b6bdb203ef658196f426784f3f40ca0a74cd535d25128c136b2de712a5f0b82328f38a0545e07b71711536f35de60e358d59dc975c6939f5da65a4757f7b9e8234e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h337dd59b877db8dd752b72286ae5f22873ceb762fc6bb034ad4380a9c7de10333fbf413999903936a4c2634abc08bad682e1ad4e7856876adbf848fe2c02fcaa8fc0767c7a648faf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9948ca21dc4e5587a1aae861281e3d80bfbb9db231301c639615a1765b9e6407384a735791a6ddb5f5d2089388d3fe082310c2d59e0c6fd86afced1bc2c88b75745854662a48e1a4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8a463e509d26ffcbb4e8647f1745221f349882d60b972d9e1d8a60330478b3b0355ca39920385bc1a4648f174b5bde4e57c3fc2a20ec9365f033b090be9ae413875d3ebd642fd0b3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h226060f57fb2492647bc5a76dd16b0bdfab7308c5ef0b52530cd82101b40e8d01f7bf0ed549e4679101aaadc16979b475015e4810d4166529dc74568f4af32454f85ef5d542b3311;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h78ed57b7e3399e3a68d054da8305098e4b5e9dbf9bb58f22125f9efbf01423553adcb8dd2a81b1a94fdce7d5ac2f6c8c47ecda7b2cd5118a9ea721fa3a06114744d5c6542ea76554;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed3cb2b1cfb77a39052fc1f13d437a0e6759771d4727e00002d7c394d999a6b2507dd3f4993ac2aae4837ad69c1ad1f42d825b754f804bd7847ab551af2ae1f51acc35e14193c018;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf260933df1e84e2cbffdaa25d4daa68a1850fd7d4edd884ce85883773bd1e9a974471896f7f0bb1d6b1ef5893722e9ae18ac7bb32b92450c7916a426df6b54975c43b88b8b1c9e0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h18b696c1cd221607f2c56dbfd1349efa6199fb4cc3e919b8436dcdaa85f230ed51b583b3a0081477618f81026d48602b10932281eb4ada5e8d2daa8eb49aceebb7a84dbcbeebe5b7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2257f9e18df61d6d91b471fee378bd6e99b86a38c95de3161c555da1b00e1eea3edf525cc1b8f6b222efc18b908329a1670b3d94fb90bc7f987aacc7d8f408f2d5bc71895bd6ecd3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5891cbd5de9de34540ea7ffe9470287d2bd6a2b68405678e9aaab2e3f28ccac8a660cf4d64d71426d338cb36cb8c908ea9b3c7cdaad781d32ff864e50f305e70bcfaaef8ed7d1885;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdcbee3c9981029a560db4ecfb73a69e4143623ec2d566adeb85e6d67a6b063afe78869ce2abbb10c2f515df62c9c5d139e5ea0155b9364ff6e3094e7a9fece5ef49488b00c19fa88;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h48ec6414bcdfa909473ff078db287f964e799ed83184cdd0006e34f22c9135cc8d663bd0411539460eca477ef7a16a507c836fb12df54d58f22725682cee845a1d128a7654b499d0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43b8f786f59e18d8351505fa9b60e8d6eec678041f0f771eac4b479e38b6727eeb671f976c74ae95e91d1780639c3d83929e58de375aac4370f8ac0a79b6b7902bc7b0e3e7bd02b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb0d7158e3e2231d1fbd38cd394af8d03757caae0655e6aa3ec7d90a158da5611e3c95e81d4c242e7edda65c1543124668d9af47908420b53573bf288487ba9983be355678234985;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he3d782c1a8aa541f72f051e09ccdb85f03db43041a4ed22d77442b3eb6fab2113d327ed04789676b100128ff6bf62145961f27d0420ef573fd588a9f7ddbb1d22489e4b665635448;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'habea27b99fed71311e4b8f33c7ca7a24af86df9ad3f39b54ea606fcb42c12b84acc6e71d50ecc9c3f91c2e8fd0135d4e7458f190d5eb782d825d41cf5e4f82015ba5e0a0afc8666b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h890b6104ec77e03779e2eb653dfc98398268b558691d4c5a10a1f1bc24e5eca3ec1f7adc11ccd89fb0afa6d0440ae3eb6d1abe1e6a14c89ed2d231ca2adce04522bc1aa066ff1596;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcd03300c4b3ed813bdcdfdfa5624ec4c96253f89ea3a6292f4ff79f2b5bb2dd96c7ee5d85d81be15d3fe2c9af217218cd3baa3c44e573e2d9b0732205aa47f6e1e52781347f445f6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9b2a4e1e819390d068b1dc92672e348149729093e78eaf5242b5ed98482b16643bdd6235926a03083f0a573535d2035c5259b929765ff89a5b7159b177b57a6c2124c40fb3555597;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h58ec9a4a8cf257a459e54cb17db7425028156a10a579a9a030377e90b680fd7ae6bcd193e72a3cf0f44f77f9b8334c7dbe40d3908fa74aafe35927035f36448952728bf16d1349c8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb2dbbea4e186e078c788bb2d03e99e24c80f52d2a49f6dad2c918331a16355989889dd49c3ae507cbc0c5bb544e2219e4dab8dcd3ab3c5f0685a2edc49d6150afec60ca56bb8088;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf5739af1a7620b8c93deaffc96f9a9b0f551f086c78cab40354dd186cb193236f62bb72408eee96d2a63e4019ee7c3dc8fb2822ae647d072ec05cfae03ea0a8e82276c87a662c921;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43cb394dd729803c5f7d6988e8c69a430e03712922fa2d2fed3f8d73af8344d563178454adcd4ffb322f58a3f15204bffaea398c46d3630935d84913360bfe6aa29465342f2afc58;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3ffdbd11ee842c2e3330eab47bf854d87fc6de5577478fddf86a2f0fbb31ad375ffb7360fedb7c853fdc870c4ef16ec4fd7e0cf5bf4e69b0a940800c9cfe743ba558f8b73cf4ddf4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf11b2727d3a958a2d80e6382d5b2122af5d8728e074c1e724869cc14111c9a0ff7d22da5fc41e519ca6770806e584a8a9e9e96af204cc532b4eedc9d192e6bcf2bb8e8449b744177;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7be70b721365ad03efb35e7b7566ef80c5557d309f329fcdbd0133e0439f3777c887d4f8358dff47e78b1aee5445ca49d9aff533ae2d82a9159827465ed9d9b09a37a5635ce1bf15;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55d5c4656f0c270b7372a4714896f8932b49568d79f5e595cb2f7779f2033f685d50bc4ea46359b7b0a39a96532e1319e29474e0ced5cab947eab7debb46148ed66467406d46853d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1808cc0a3cbaa24a00c38af83df26862a9b7e2e9e287410f1514316af686efb0f9552aaae6a647193b9bd62b27c4946651a9e0d062d2a08b2ad91a40bf8a96f9836802ef2341579f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf89dfe9a50cc2a9d3bd09b4a14795eed02a7c106f057dff269e58e166cba888ced92fadef5d149b423fe755d57d010f220f6027a6de24c93ab715a78b5e9d73396df61567558457;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf674776bc16ededb9a65e45f5edc78e3e2b0fee7dee3657beb002f11ab240b312bbcfdd8cb5c67a8f028b75a0c809ff7efa38cad784d17b1c92c3eea101e53a1f7ecbc9cad459d9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h493117571502cd52cc23814fb37669213b3ee7bce7e3b5532bb151f531e3c4eb681c2783a6377a57bb2a8074dd9a5df830461e21f02713e90515b642d69e664b53874e09620c41c0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ce2ed991a4a74cc90b8ca46b4dc5a3a942474b1e6b36b00a06182ab2d9ce0bf83d319c4d6c45db95bd9b28a1036a46109b3ef782a5c5c6d814ad37914d6c7ec389b3953240f8b13;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd05c3d99e5468a40fad897e110e83d51c5f5a16748d792dae41f6ceb3ccabc41c918f2eb598a63f234c86f2cc76f8ddb5e6c2c24de3850aa20576c3fab8b1e0338995a9f35495684;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd701d36f80dc56a447b6d18af27af70458f55a05cb429683b3cd44de7dbaba31aba726d48eb9160f8703e429a187608abd0d8d0511e83fda04d808c27e4c572293a8d43a015def7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h34bd8c4d4656881f18be4d2e5a388256ffa1d52560e3ef076aacde2de2eda07c0073888cb5f5ed06b299c372d3b113f64b64d410a01f742ae9755d01771ff2f182840d4d1a186c04;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c55f4b47962b474bfb331af328091c28291d37017c36d571670d6979d54abe6d3517c3d535050aa8b5a27c4b01a069d7dc4e4b01ee97e577145e23f68ade3c110e54dbc8849a97c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf3b22524b2b4593ff85b5751e046d6c2cb6f9cb8008023e381a5a84b8a8dcf42932d0c5d3f69383f4b41488a46bf6738a67ec548095b205c39c7a888884762ab86fba9a0c36a1d01;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1931f35e8d4b8eca00ce05184dfc8c92fdfa7428ee50849e00508d6093341f774769749e0278d4e053dba5506afedf3b65336bad8dff71d19a826984c6387cb077832697bdb538d4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf85ee1d3cfe4f37516d861192d7161ebd6064acb56347a505866e577149e89e22c2196f3844456da50f6ca0e3e1919291fe7d62d7e46d495a744228b0458ebb2e1c7e8b6aeb69546;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc82e3275ea2499a63a1ad5f1e0a7e85ac85cd32b1d3fd1e99e21b48e65bbe1b38541ab768a930c4d1c292d0e0f30247eb112999f7867f34abb330cf7b9532755fca169ff663dd1dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99d08ecf2f7b99288bdf82cb719f67ea4a524422fc12d735c9b470b3d79e860a6971cefd3460effc5e3a9e334e0ecf08917755702d2e60fcdd3c206780f947b8ed0ce697e0882219;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hebc043b66d66de6a715c292406545a80ba2decd3e71106f829142c3921057aa833aadf07d570ae4c7b2c3ae0b4c0692426c141db47e86d3da3e5a269f98106a52b4f4b5c8d794661;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc31a1c8b0bdd29a6bacede40b77e1f559615e412ba2433623aeab142ae87f2a4d3276efb4bb3422e90e28f96fe75a6b1dd648249980acba1b56a7cf1a5ef30d9e0c4f271866607a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf2f1b78d60866372353c52153f11f8faadb1d49a3b194648f0367cea168cb118f8f1d8cba74a879309cea4ce1dec3cde38d2a16f56cb7883baef867d0c21269fb59e4f318d1e59da;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1090614ec29c119b0aa6a5a6e412e3debdcc36e4d56e64ff656dc0d22d8c1188d9af15a16771d3e3fccf546f6e052f68ad398f2e4d6a6d379410cf8d1115722450ead49b9fafa769;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h24d8bdc1be23de255dbc34cbf1c41676e9bee98ec7f8f3ba691e404090fa2142d7ede55365ac4d6d737abfbece959c8d82a0125d25b98e88ba8b05ec529eddd0e7f07ee0e982017f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h33bb15fc79d865baf8c92da4087af377c9d8e88cd76f906a645856e657dd45df44ce58b4f089748e38089f57808e6611f64969cba612eb08558ff60814e105691f57eee5b0c65860;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b1e8d7611ebe9a3454bc9758475ceb00c6fd350f1263e8ac0740fb5bd71a1d8225c67efdb8189f6633ad4191687e03b6508678d41b77a82946f83d5459124e017e76191e5eb763a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h799a2655d698fe966d0ae5025113a87d09a474683d9e54a4f6923ff832d0dd7591ca625b82ae4a959efebc78ee24f36081ab836515d2b2ff506a25899a196acf1d55fd8181a4a682;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c83c6b3b0be94adb72d93904f6e22c5dcc114ff041460f8bd502da3f3b19e89705345d18482bf5d286bcb344c5e2bd94b2968c20930a01e8af7cb12f39dc1259fd559dbe614c196;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3a4d6947227fea5525fd3047a8950009bf18b36c9abd21bf397d73c170a868dbf2da4b591c052a53e071c27cb0f5873546af16b4f4183b44d3477579aa2851754ec05995da8c036;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2d29e0f32deba447da6f7c2d4bb09e9446b3e94763c33aaf2e9ef21e63942003856abc291d034b8c7ac715e279e23eff950d66ef27f260838b81c2b57c6ddfaf5843be1a5b2ec9b4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee75ad1a7f96257deb6a0033a85f9a63400bdc1b83c42627fc772839b5e6c414d564a250fa3cec76a9ec1f7b356166a1b465f02293ec69bdd3daf84f508e38c0e03bbaba0d524dc3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf0e3abf037e13e67ddd6b7248f75926470dba421e7fd92b265a1d1caca5e207dc5ac773dcf7a49edc24bae7057f755d6100023629adb4ec56542c18a2d2dd6991edf20360428f1b6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h30ed6a00b5701e620dcffa8006e5015f90bf058d3d87e86bae3126933d789143e6c547f88bb8e4cec79c8a41e32366273a0291dcbae25869c12bc54c9149588e8457bf186c65e838;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he770073b343632fff7749ddc51a0e46d6e1e9b963cf88b0d9a955a32b73327be85dadf99d22a6b59c65f6b5bcc275b3519f453f8c8872fed6b84dedd957b83eb912cad69d09eafda;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h98aea3162657ec18597174f93369941bf814ccb021f27f6b824bdec020543fc3dd2334a46f3210ee2aa95eff8d484d8c4c205982027c9cdc45dee948c96cfe6b6cdbe055f08df26b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hefc1d74bd8784505912320e36104782908da2aa89aed73e8d2445f1e9b4bd5acabb90835a64c16c5ca21a850f09444ab8df32721aa61d5507a3356b6d1cc5966662465e9d1c7d17c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd093c3dcc608cf47167e74c225df6cb8152c64b29ebcf95c546b0e26afefb7383087f3ba388fd4f90ffcb01a116aca1e2bb0d3f1ed35b21784a35850bc73ac207b8b81382ee893af;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc08e0b7f5c24b2f002ed924d59343e3be6189bbf287335f1c04c9f94e98e22f386c3be6e765e1dea2849a1c75eb1b223c9d07c8300f43992dac8b3164ebdc16d622088517e8c6440;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c41748129b6105a0663a32a6adc8880e8978ac803dbde8aab597f30ecdcf7426364dd4f7f76d686c0459434fc3ff3e00408ed39d74cdf76d36621baa06bf86c37c4f15fa20ce0d2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3aedc6d2ebcc1f1a02b73273aa530effd01764b42e3fdfc00345efebb07bb5cdbe0e12f4e71bb37516802ed897ce52c2fdf14ca6edecd2f049d5f19e38acef6c007f0804f9928c48;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc4534f6aa0d853b85095ff8fae1310bb42ab5bce37c1450bd4485405d64c764ebf12eaadbbb216e6ddf2523670123448f572ce8b706a6b72c7fbd633d7d0ad83c53e26f49e96f765;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6474566ee662c0062d5c2f150e95d40e53543836ea45356140470b6950ca206857786b00b299dc3a2efba9b761ec3d6d61fef3a9029de2f7c68bc8f4e55c07df11bb196ce963d6f5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3e73481d48af9cb79472295fc5946ef9a3cc04b1a579450f99030189294ab70c3c3172ecd17fd625b195db8d2f7bb37fec9099e21d999d6a72f9e1b8e332cab8e981aec82e3922f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1d9247aafccd3deb0c5752e37f80d552920bcb4291209b3b67382d288d2ef34babdc7c9bd08859f4e1baa79e338974380fcc47222216542972af271091ec68a0fdceb61ca2f3692;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb104251a3445e2c8085cb59156235440751909e688b5c09ea28ba30fcd5b5d995f2541092414ad76d489b2dc2a4d332c0de346d39b8a89e9912cbdc7e7a1be84fd697fcd12af131e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c1764d7097301036290bf8aedb49338df758f8ddeaa44e837f2c3fce32894dfe44d98d55d358f89992b1718c26ec42ab33ff3d87fc707900b0d281acd7acab88ceaa743c1f0e3f3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6159131a7bb11dc5418ffc045cb3a5a26071f585ec451857e2fbb31c9289bc557d09db0cc690c12637af4f8741d7bbedf891cff75d9d0a4cd2dfdafed56d043349048d938db7c7dd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb1500bf11eaf71cb0d6980c4becba1e062e6e33859254b53cb8e8a09e772777eaf182916fade6e93a5ef67aea06ea1552da1999d93830dbd17030aa7f3d89835b108453f317bb6f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h25b5808e94cc2bf4190b5d3e2d29c0accb44e091d466d4f0ecec69851e33b15fa0e91b95b5279363b49c4c5b8303808c125ca597ed33b00c65bed8c77fde69459286fb0ad363b2fc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3c83b6dc88067987e1036a0205d399c5dc6e43f01185361c55a0bd68467677f0cbfc36e462b581543e319a835662be73da9b21ddd2335f0032198830f61a7173ec280c64b91e94a3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h589766c9b617bbae49352e2433df3d66a15a3aa9b8d3e8ef09b7578d39a9b85a9d5ced2efea7aadbf7b2f2379fc7f1b69e895b9ee93ce37b9bcf1676f9949a61f4ee7d4e32c3e44d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdee02561d21af4d22568a9bed85669994a8a6de8b6d9a80bb8d5ccb0f1f6be0a5eb029780fc34af7b6b58d48b3d12b7a06c1e88dc2bda8e321cad0fd2234d30a4f6fa2375168d2f6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56031f02c6c5fec4a5518b07c56446b195f31e8a63afe49091d64342a7e2f23698ea6f3dd70ef9c9afe481be4f56e5d2de30607ca7e17a258e11027592664c7f778039f4261edd86;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he4f30bff104d232e09a9debea85bce397047aeaae49cbfa41c11040aada404acdb9b336ceeed51a9ee17243117d5a353c2875ee83510134002a1af025f8363a132bd8abef4038339;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf30d71ba53072f2b54903416ff5776f6ddde284ea1a3fe31dc488eba27eb8d25b31d77fb50e6a0694d8b6da65144185b475f84a319773c499c2dda7af8f6c9311e13115b6c9744f5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb3a8ae0f3dc7d7acb5b0687bd7fbf1aa8b3af4eb43040f7340a20d833ab12ac4a0fdf5016149681393054af9c02bf15f3233de42ee35e5d66d006f3f13ad5cea7c0d53685b3b45;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf391bd5493923d8eb8941e47d8f04290330544d26701a914f73c941cc069938c608c64525f330debd2c1b03521603b42c16f1e6e19f8bd86a493cd6325f6faf348019406d4a1f057;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h555890e60b01b036d7bf2fc87ff4e121b992e7f9ff9ba2b1e6c050e578d67b995dca9cc5e072924c241dc3edbaf23caf3b65996a73da8632171bb62bd3b8c3d1e73d1977fa1e8a35;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7e942340ddb829312f3535fdc96ecfd9069f34da401181861bcfd7807b6432ff52b60c7539d929dbdbf72a80cb32d6e6f827893d965cc6f7ee221535c701fe2537087b62948903be;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2eebbf8d88115ebf0ba7b0c53f4b120c9acd6a0ab13688dea5f8c25d5ae74a773d6a160768295cde9d7872a047e6a0c8820f91d883bdf7180239f5aa79f7a668942e8d861341fb49;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca03f568b17474d6698424c2022a0c67c6ce80c4c5d13629efe3d7250b12b07e767362711502156664fe2f842487f436a0857a579659ba17cb4edc16c59ae675cf760e5faacfa2e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb474f9f6bc5c7f73a559a9bac76373e3be73921af39a75e480fffc0e39c7338e542d2f5461f511671c1a7c6b6873d6d336f8203fa0b22f62b6863d205f2d2a7c0781dfe70df8c56;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54a63726d2863a730246968b7a8e76e6f23b411fdc5ce0f90c38ca7c75cd1e556fd61c7b91e556a673efbdc1613a04e25ab846cf1bb334094c29340702f8b3216a62247b01a5b26a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9977e87b4323d265b555128a18a907538a6f1943cd556e5ce157567d19c80ca9132d5cf8b76a8ba770fb2cb7b4926555122379ccef7841b4468f740205e12643d6f0f3e2bef4a938;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1dee804fa91c0dea7792fcaddf0b62766d98445b5407a97243191c11e61118a8593513909520852dffb84d087673a006d58c1ef451a36a9063e24cf46c3fe5dd37fa3b79d632f5d1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2078c91e85fc62b085b347523072bae6f9cd657e27bc0635523b328e4cde24ba09d6fc7e7208ff3e369f58b7049424f38fee8a41670f1b12d4bd1f5b245e8196c640ad4e6734b037;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3610ae6a2bfe323c31c7a7bc58ea9aaf83aefc5ce1a980bc6b1fa443511d9e0ee573adba62e768c5b2620d4c65d33fc0d69925f4728e509a6de400a740054674568727ff49c8dbc6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb0536a1ad7bcfb9456fe2164a367bfea6432d4244a860ec74a9f64d08f7f85c59445ba47aed57f20eb1550ed37fe7bcdd70ed9f94edee14a73559cf4c753297d2ab1672106b1ef9f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8b3341e9768a1c675e01b49a11de51dcde6174b8349fc5098f9c8e1171b5299b8534ee2b74670c970208bb2200c4bcaba56b9e35a18b99bdb0feaf4c4c3f26a2524cb2f2c665d549;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h804dadbe8c95c818082be2d09666b034f2322c5aed47e476d51bd0a749d7a447306af81159a677f6536e2b81e95a896b974e7772dda6b689a322f427d686809de6f89037d8b484d1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha3a44f64c5b25af45d37fd965373df2a635a8448576ca8d3520fbb7151ce84014fa584945202fb24e79631544e1cfe65ccf5dcd0745c9d0f5462f47a4805d222c6f8ceb7671a81d3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hddcff1a5a71fe0cfef0fe76989946c5c1a6250f1dfd70e37e7addd24cce194a4f0fb00e212919a679846b7f052cd3781b7dd3e9451d19f47d5e0f723d00c2958a4903da206bbabfa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1acfe7af91054db79d65354ad07d06a64f4d41f22daf0cd5498da52fa1c924c0c9be1605a5e8b1bd6aa7839f32aaa91a71c6c21c510417037fffd4c9c9bf8628813debe801dcd5a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd705e3732edef92f2d8f84940b65a8f2c43e4b9411ba0fbcccc18ae2e113b18685f35ab7ae5b656a926f7930bddcd87378dd0188bf4ed37ffaf6da1aa044d1149229b93ab321a74;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52ee0e0b43d06d1885b0bc5a75470edcafec64e64489b6c95be58df849d03471d396c961ea233ed1a707736b7b253c1b234e616be5bfbec487879af0a0b0648dad638c3fb173b271;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf63e4d6d8b69bc766dec80cb49e7b68ab35139e0f392f29e7a0b41a71d60e352e5a9083795a6821447caac5a8e8d609f9765b8c2623babbdc3a371577c4921ecaf2d9f9544322e7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7a3dcf6da9274e576da958989c068d2d9e6540f82db57b42035073c5ededc70578f09cd733dbe4dd8a79fae9b69532e73ef036155e804f8ea77ec02fb65d6ee0beacee20e7b1c2c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfef2758836e622cefcadd3070595ed0ea9f3377c34e6962ace4adbef52c5dea444959f1cb69e07a0d4dec6b52394f701aac7e865c28258059e06f7a5047883d4cc4abc62165e4462;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h79fb595aa25655fa04c8384a220aa42dee79e75991b1bceac0560088fb078c1c711abe06e873b4f8b19f122d3316da147865c79fb010ab664a1397af3d88fdcbd047dcaa8b4a8a7c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee200a57557fc4ff4825541e4fee629b857f2d53b76d4ffa1306e274a8e616d5435b53f14e191388e214d661748cf5d6fa18944fc5a7d087ec382e28089a9ebab22dd5ea420eaa4a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5e46e8e8491df3ccc38a88b2c937f865e23409456791c4af90fef2afbc4836a717fa4f1e14d43191caba78abeaa2a607706ea03fb1a621c584c8208fff06fc21adfde6235e9ce02f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h30d2b285b084215631e310dd5943265abc1da82e6339a953fcbefdffbea67520dd585dfc34026ec3d9c8fd7c0e088b2768a1a4e166d44e2b21ae644f879f0e3cdc79b3d7de177801;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hda005dbb4306a4d7851474d424a57404335ef7d690d0f363be649c1eb1625e36325b5f0e40a6b929bec423ab97f7caf9e0a6f81791e18b7c24cdf8b7dd16ea67f0c9c930e7f586fe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha2096adfe4ed529ab5c25c09a36d04d77805bd87ed2da776d03da677bc4dc51c56ac1e6440faf846dacfd3c4742d291e5d7661e211e8a83c8af07f07539aa6dfa5724ba7a0d15659;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h704807bfe7185df6fca8427cebb89715b06a15d88fb4ce9ffbbcc4a8dc76f4aa5495447f00cc9c65e294b4afb1b622525018f473a966148ae645ff1102b6ccf5e656307e52bff0e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d83b6befd0657ba2cd8ff98ba0e654db50a1027d29c4fecd43f1d10701330488db50ecaa8807852ddc0f877657fd922cedf7a4b2d6c0711e56d05c727673d3405b8e6f241f1f01a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7010ff3f022a3c81a6d3deaf5654d2616a22abf1e5dca84dd127e8d1660ad5e2946ae730127b62476e71c2b5b4ac67e69c58a9a2f2d87d3171a7e3f6e267cb1a778798b0ee5f4df4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5aba6357bbe2dba75cb442b90e1caa254a696e61049b5c887301ebec97867408df5137e1b2705765bf880497572cc91df2fa3f31e2da7b387fb1cbd29b939c46a9de149c91255007;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b5b077d4eb6a12d0b657880851125d1415da2108793998c9d35328251bbb786a59572812277cb81bdd272c0fbef739707ed58e0d7f7a183e7826fad7c2696da0c93d25db4a615a1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h49531943907b44dedc0e30d63be659ff9d4e28f8bb298407c70ad271d48dcb963c8fc3cb60c7552d9b7724a4f550b0bee48fb590a62cf7674c1361512789f6178c775089605c7c50;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h37536ed80219f605b44245778692784fc363e117fd6ae7f9726afc483b5eb39da0132a5962a9a0b90764bc58091b5ead31cb2cac3cf4bc4e5958ad5ced93ad5c271fb310f92deccd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he429824954d83369f290e1ba3838254e59899ca93edc18ca755ee25836422aabc256a3244dbd37265d4dbf68ba16ad7ca619e4e26b4e3a9d639444d8d4e4481e1960df7e521fade2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h26010b437e233cd529327a1d91a1cb6c0627848578a4a083b343a054bc2fa0851238177f4556d7d1b2dcc85ecb224f361b39066efbfdcd5bb3c662aff60137c0ec509ef25ad70c88;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf69514327d4abaf2aa250169a61baa128d509b2f0b7b44532a559b62393daee4b3159f8d76d370a614c904343dde2afdbf4c80e52f791daf7b3e973397390f29674989c245d0dfc7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9413d4abd12a934590d11e0a75afce6d81ceb3195acf84e9b1a7773297e76932c793762ebb6a9025d29614978f8c49d24488c2350a82731896b525461ffe09ef82c0f6414aa65ac4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfad0585da970e424955721d76c2542f16e529cdb0f5fc13f7abd68b1be12533bae9a6dc045c4841ef73607a11d106a1081963f65683254d7bb54dca3da9b34ff3ccdde237b6c83ac;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9889166a0c92d386ffc007fe9f261d35c4e725fd5e5c468870a29709c89a670dee6a01d676ad86a622bfcea6283b45b0c87fa6a7118ea53acbf5cffc1f9e009ef80a3857999ac08f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3a90fc3cab6b43e43bdd671fa14818584e22ee7d53572e1ba220a29438e0c96a4fff8969cff43e29524e7f92a246c13012de4f77a542d7669998026ab899e0c5727836abb6009b70;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e51a3f0a93604b736ea6ed8d075fdc8dc8c855a1e1f70480f7bbf2ff4fa3897acbd652a873af8eccf28c5205d47e121670ca659add5cfd6c8ac2a550d9dc9a2a8b0a90c6f76d3a2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6fca58b36c98363cf82eee5a288461f26248988cb5dbc567c39525adf8592881d34e0685cd02e904b226125770e0c44747d5b358fe718daac01d65b87e2d873b073315b145c789cf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd947afd4d45b3cb75a6fb2ebf1dae2fec490986f86810075b417949d82d42b4d9ce581e06b591f1e4bca5091e3faffff230e1903c7ad501d53433a78f5ee58e8f4133882896d86a1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94f2c2db80dc88e01102e3de8515a7b3e4b2bc2758f9fdec6cd61eb13ec281256075311287329738eccc7772528016be1559f8da80dfac8282a454984e0239efa6c3fde40fb3c10;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h576b46f00981f2793d358b831e5d549baac7234fbc1948e9f202174a1680eac2b60a22e4b1ac64679254d72dad39a5b1209d97dbdc547fde2cbcc6db96132787d1e48e710e2930b2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7899196c8f8cafa19c908948481fc7a6eb26fa16c0eab2d20158e318943ff1faafb461592bf277ac0b5d83f07dc79c358c8b3e0218385501c0075b7b099118b7db854ef12093351e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he9b26140a66f95809b88100a7c7ab7f49b216f3b04ef5aa484fc99cc380f05c2848328e5959b526a8495d58d935c27c5d7e2b2503b52e6b284b201a6048450be74bb13b9fe8198;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbd6b4b1e3c9aa26bfc08ce04da98873d5851f6bbf6c29934793a094eaf1ce29fc04889b8583d4ba48bd831dcba204d807056ab140c419e84f89761661fceababf79a065af92549eb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7783f9329ff35601c973debaf491893a13cf58b3bcf33497abbce1738ffe948ff9d0c9e20eccfea8f61c141c01c4b6cc5386f6056779ecda2955c3f66a24bc637b958cd23e8e49b1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55986a77b7cbf1d14ba32fa953703adbfe0fcb9cc87e63e36d747db6f28d31b5c9371dfcf60bb669bb0ff83035941ad958a72b7a1fc73df6b6934501cdf4e8c7e2b6eb4ab9f106bf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha59aaeb83b50c236d231add7898083007fa1ef9e30cd814726b3f4104818c676e0131b405f623972d151987bf7808a98cba9916a81b34f08a665bbab28391cf8bf189f7d2ae6e727;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8098e5943a1035e384d084110f8021d009271a1127103f3ef27584ed57034854d8e5861a95235fae09649895400cd22f3cb2f979d156bb841562e504a0162198daabeb45ac655442;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2a69384e28bc44e70ec9ee21d4d23ca1ca9b6f8b80e7f9b49396169cc7eafe03ebc4bbc0b36fa19cdd82fea40c72e591bade2b6669770affd45dee6d6c65a26a6a0d38e232f63c4b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h80cc79da9552070d003829be5d178e5840b0e042e67a02c0279f53b5947c672df0c884a946d33f9106033839e310b7c698ccc45036a1e841718051ef70e714bf1481ba1cf68b60cb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbba6543e9660633b612b74c142ae234d4f2ba39645fa77ee1fdbf1adb2bb96b125b70ba9554395898a349fe4b6cadcbcfa6601808331302161cbf93c1d42bcb68fe59f08703d3940;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9982cc5f14bda6a999e36f5d9c1c103f3fe1ce41a790956d43faa2f74c3e6c2eef7cd9665986821efb5d0f7bd180e72cb245053134fad3948815219b1f76bf9678e5ac6fe9827d3e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h986df7b7186466fc6a809681c3de4d5f37771d564fa12cbccd4787eab19e8ff811921e5f63df595b0f385edc7cd5d2b1c55cf34d927e31f31802162cf8b0b8420d7c645172facb69;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha18f824a678d98c7637221e8aafc7a9beb6837dbf0bff7f98152e0a1a62355c4f703cf936c4ca275c49aaf09dd6d3ffd8262d7ee845fa27fc95bbdd27c70287d9cf2e533bb1be658;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc327212c817bf65e1df29d9309ad9e687c7099a64dbc8a0e977b25087430cf3eee2e06d34ead59b676d0bf39652086078457a209e12d72b5d3b6c57685a9bdfc25736f3706f6b7d4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b99806c606ec9ec65e13c8460eb2d6a9483c5c98c48db2f637d6457fdce272e6391f8031fc5f9457e921d9c1acc6b195bbd5246f9bdc3f856fa5fa1a1b3da79a2b60dc99bd3ddaa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcecc6d34e32f69d7a6b7d81edf6a0f7810dc1a0ad1d2cf8faaeb432714cd1feb68a96178185964c6c6330b0126f0bf9b3329b4cc0ccab8115857e7540571c80bdb657cfd5218b7f2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc7cb61dc093d1aaf49cb604778e77b6002adfe7f4e4e8832c0c8eadac9fe758e665613bf0e49eb719378663f6b7e386bb69f5aeb709ed2665972900df643eeaf519294cfbcc8bc1b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3732f2e08511fa2514b7ed00b969849742bc1cdf103d1c5b9ad0bc84d2fa41bdf884600f9fc9eb994fe1ee09d7c03cb429fbb3ca8687995a0931574f33c0aed8b82752ab3c800c4a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9bb6feb861d6e8c5dda35b77fcae9ae1fc695ea4d2c8a73fe72ba9f1ad6e9ee37db5164873a53f5418a944d6eea207380cd95baae688468dbc1fa6015661a843b3c5a5894ecb87bf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h947aeea2dbadad36a80b161301f41bf205a147a41d4399c1cf310c854253e0b0543340a934c6f92c2a0f0f5ae769ef2497bcd66e81568f5ffd76ee883baf646c68e0a19cb8dd7af1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4e8ad209d7aa8620f1fedb914a7829bd69ac84e4d2fde16839b92b8eda9cf50f6fc621dabbf2c0c40767d451503d05c7a1792e4c76915230524a4b3b308aa3a3118c9a84238cceb1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb257a6be78ecdfd5dbb1b9fbe09530287df09c7d5c5399fd02435039c2cd52d65d6d1eb81ae68d9e35064149031069d1ce903358720d815db480071b308ec64ce7281d72df3868cf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde199fdaafb190f4eefdcdc154b7edea465852ad2875cd124e3dd2b1f1755cd8b420198b106997bf07d0b4c06ab5fd70aa25a63f2e467c64b18e45a8f2f20727a220e15d3b165522;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4f6394aaec308d7e45ea2121474d68942d3acd071280256e314b731eb0f4d56b7ec6dbbdc32d0c8ecd72c64695f4f479efbc8b01963169acbe5ee476fbb14e5fd3a72e02355e8d46;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74b85e60b56059e5e4daa8bcea77a14fa5d3a62601cf3252433cbba9385e47020aad0bd8386c6bd0ebbb81babc96c80227f8d172e968e7296a2db20f4dcaac3bc40929575fe7740;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hab1ff10c10118a4f1afa9969bbfc3e91fec771682308ee1bdb0a5520576be2e322b7e21ee5d63db9d76c247084ca3f16ca79c96d6b7199d35e83c98726074b260f7edf181dde0d20;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd38fcb2362afa2806c35f5996084e74c66ff09c96640ab49f5836e0522478a816231d177b298d3b50cebc61f8b1099b97cb17cd637e9592a1c66d3a57f34532ba93df36e0f41e420;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54a3c2b275bb4549bab4f49761f050fe5d63d7c73df22dc32112ad0700f5226c75d9a037ae508c85dbd202d16029d619966303b79cce5041f4683b3f0d49ba914fc4e2552ec5a3bd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf47884034003ad920d2495780262808bfe0df1e58db493302a8e74b5e6d592e3b9a28fcd410bcef9271ea118f95900ecbd72f4a3bfe7f371f3565ea97ef2d7ce438fa09a500c40e7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h124e80f34ef8cd4456e17fa17e07c5efa89cd5c1ae507504ee3e9008ba3b76fe0b294c68c47d1330df2f37f2b74732a40d4388e269573e81f74c1a64046fa6e4e01aa43d64a28d69;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27d0e9315250ae36fda326ccda1a69e16d6189d9d843858d2a4058fac262edafb66033c8d040814f44c66f1c7d832ee891260b473e64b9b21e635fc597f4fede986a086f511eba7d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf9c7a8ab9b96660f417c06ddcc262c7fb4b89049fcd2ce9a1d7ed73a7a791619dbc59c5db8689eed11f5b7c6451fbf3d7022fbe2943d884c0fc83f7ed3b46863f603a49767ee5fa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h67dc8479911dfd37dee6549933221b68ebd27245b1570786b2e5d2fb79082a3c43189e2a91ea4584d99b4bee8bf1648793ff928e92d07df138e67ce0cd72d5dd2f8860dcfd56710e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf70394561a7fa3278849513f5b0e59511c379909317011c944cf929054c0822529f4db543f3b4efb7e5c3c7427b45efb86e9cd0d519942efc8796471a7b7cfb9c583d64f6f8c36b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h816ea70a981f9900ffe5441dfeb86a9cdab34817076bedd7103ad887d551e5ac8183ffbc5a79c0866068e4dd6ce9ca1001079ae1fdf79551f9bcd5ffe890bc13e379c4fc641c46d9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45b81a9301d25c1ba67012cf8ba373fefc8d8af54b845becb7cc5ed6cdea6262bcccbeeb214925784cfb1c5c20c7467bb5d3fbc71226279538701fb9e03a46b1d4127fb54fdcaeae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8f97c870c6a2c307e91d2ffa831f29009e507635449fe1088f8ec709aa22ba5f1db9c3e5f14ea906c2435bc00f7ace98d75f9488cf2b687b37195401abb576f6b0ebb58ffc7e1799;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc0aa26db1f080cf1ecb043244488bb2427b1465955c7baac61772947b0ccb71cc2cc950b7496e5e1eb619710e659726c5f2869fb35819136385466f4138e475d57f26eb0a94b9a70;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfb78ee7349e569b54e7ae08507e021c5a75a7da13e5a3f43e685956acc8fb7cd9a2b2696116135b0806e7362aef872e73e310fccf2776403df1d6a35081b5488dd8bfa6be366b18f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h388554ba2c6893ecf8beedc2cb029beb49be1ef21024e7876fdb832317c737db26fe6c686f46b8b417788b45ab34732ab8902111d6f5f35d10ad9fc86e13920483ef0134b6674e5f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h608f50e157cb022cc31df46abbbf92945d9370e3bca54d01fd4628b3603e3bb4cfc23f2b0140bb1b294874de4d8dec1df7128a4e53a68342e0aae46762c86370ddd083e019e4239c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h52c893c2175969928289d0650281b9b1508b64c63838e2ca2cf64de1974ee4d543e099fa5efaa5251266f7b534b46850b8baa5d92456bffaf8cd963b7d127fe1242c448a4278159f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h201810cc4b071db7894d71861c652d7b9982cd0ed43ab8f2272c95e8c2b210ab79829a89bf4298697f460c9ded10faf568da74db9e2722753290ae98aa6bf830c5dbeb810518b97d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f25adae3e9f95fcfaa64825fc2146f38b836feebcf05c52567d39fd2b828364d230c9b703b932ed2ede6c1d09620f3180b8d6b1d07497002563472ac4ddbe51b8926954f38882fa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc6ab0188790ac78b9b7af9fb196d8ffb712bb10ea3b5b5cc38006490f6cb8e1c89b708e5264bd0ce8ff4d79d8c90cb051fc24a8318cea38a027a8768f1ce851383529e39b9aad5e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haab587c762602d0673217ad412cdcc69ab179a90daca0a6205c73420190c0b8efc50ee48342740e998d5c76325bf40af4f44e4e9485e0a0831c4d5f49d73254de021d9723f7463ba;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h45fca6a31292004bb0b8dbaf22ae9dd61bfe78489c74330bf6e681a054f9c0e93ca553de6cba1e3ce7edd8eaa5e25992a10f541b013fc07bbc3fabad4e9aa16ef9216c4c46eeb7ae;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2709235b226e43d262215578da1a4a32424f36587713e48c68392bca2eba958d47ea63226e4de62193998238eb68a4008ce517aadeba23d230294138331ab7dbcbb0a358c23f8f28;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h829412de7b95d2f01276dcd28d4f70117b741962d81979e23327bd4b75c95d619687a72221edb2fcc2d9827ac3061bb3bfdd0d8d6c4589303041d67d9e016ba082ff3e4efe9052d5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haed2a4b107c2e00d1bd8c9860e6885fc52b61b6044cdcdd879cf1deea8b498939d40634f7b28910f4476998684de4b46fd5fd1929de8b292b790993aae7906046ae5a56ab3e8556;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4a4983a627c67f878ace08f1c960c5f828913c4c912ed21b27d1a13574997a04a143ef25bb7979dd69b169bdec7aad43704af6be46dd2297b3c2e30a636e976060f20489d33ade25;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40c3459c8ea737eddf6d0ef858edd38b6da696b406ab2076b042c9de525b2f71374f69aca779b370a3f3b14815880d2fba12dcfd9c62b1cc6abec26c234d36ee1b4def39b4d1578f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he68dbd452725480fdeff341364dfa202709258df78b5b6d3d5525a675d79edf68b7048fb83d4d8c517a517a1f8072ebf8896b2aa448dd2cc996d993772838e81aa83669a6cc67457;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3d97301bfd5f47665a6e15d35686062ba437ce59704cd650b484127b6acf614764053c6005c7dbd1059f5c3ac9b53d90b830c7fb08028a75028922642060dbcd0ef6eeb598fa19d5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5028e6e267b63f462163adfdfdcf58e6aba35659b1f23cb195a0fc6a530177e2d32b254e076b994112c0adac649c2e6327895b0a1211dcd35921cd484a2ae68282bca1f0a36bba75;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf7805145dff035f2ec35e21f3685c1f076c1b4804b0d3f639d54281e4b568eb27ffa5fd3921fd26cd5b3bdfd9b5a8cb9bbe8942936fa3548c00cdde18d82715fd6b88936008d7f3f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ad140ebbb6e9d3af1c610ee40dab104af23f57d0dc1c671c0e0c3fc86237d01c24d0aa28246e7d4510afe17f92f3542f37c2b41173bf9a177fa50ee29f067b46cab65da61615227;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1dbd616c9a10b62fe752e01b36a644cc25539aa552e72ed7913972f96b65278eba4aafbd98b1b76f5deb2515a726c2a5f035d9061f38bbc34b30f254969f89c1b47f030c06ed5e5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h86e98f8cae85a7074b413761b2356e9586b486788d79dda57c9dc829aa69289e75a771660712fcc69958ef1a019e738405258bba91b02d6fe4b1e4a50164af3af3707f295cb5a6a3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74a18a7f0da1e5eecd6cd593f01664771dbad86d792f6286b002b87674ebfbb3cf48a2ac44deff4bdfdfdd800a85a4d26003b7e723325ffd9c6061e5768a98dd245d09b473c0f63f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h33ac6cb6ebe1e0038ccd7894445dc6b9d41f9e052fa6e797e7a648c22a235ab3b7422e366c9da4b23cbd6996ca9c801276a76b0a9d00abb0436ffbd26b1dfbaf02b7f5b18b76eb6e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee252f9703e9bf778c057bd96a269e27cf184788ba0d1114ba8cbaef325159829cc969496d1acb468e6755dec180c3969d15d2338ca245961a9f8a0d8384c46dd6d4f74f02cff125;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f5efafc76342a83dd0c1c8b8709dbdebfb320d98561e73a45e142c283123e456995ed8fa2b54b33928d999bf55c452f70043c58db41ff04a6dcd97ed53c7578152dc9d8422076ac;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h57378e3c2629d40a16c8a946912289d88d5d51696b5231d08918f72393fa42c9957f167338d35c88ae39624db926ad80dadbd8a7b4623d403d53378a1d4f8e179ec7299a765696d6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hecd6547f65751860c3f3e5d6ad47a8242253b4d3666ea01015e236dcbd2b38e76eddedb700158a4b09a97864e30a93a456b334de865c1a93cabc6ea1137ee3d4a29e30d1d7a7d97b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4224b4c071df2516eff7509bedc48a9bebcbbd8f7abe465f780bf7dd7b167c3efb63edd7ac6947d4be7f542afaa9a302369821e94f53ae36cdec5223aaefbfdcb52c453c2046f9d4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55e70027694f1c6b285c6594e2728e454442ec801d9edca89ea289b4ad9299fe7625b9cce3e664a745590e009a3c0d3c6083b9a229f63ccfa17ea86ba9a08935ece2adcb51d35f2a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he482fc14f42cb20c657ae58248f18c5ef5efe2faa87ad82d01de9ecad37864e320d1b42715a5098e6f08821e6f622440ab123dd691a4475f1e164707b1f109e1c8b441bab138f4f1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1a9eb1f220c410b824499924a50991e3f12304c767d265e786c83c893f1763d044f252ecf2b8e3c6efa381ed3298bbcbdfa300d36c848dd27ea264067db2632a5b5d9089879ec86e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76842c154016615b51897af394de82867e02034efbc3e08d32ca95321d0e18021e441b84b2413726a2b476f8633e22bb622af22ad78343313e6cf033aae9c4bda947f5973db34323;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h359d944120809a10a7251fd7b010780835027033a76a026ccd01b31a77ede4731434184b9746fef6966961e5a3499574b8a2dcbf6dd6f6c1259807d7433deac208ebca8f80f57e75;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c87c8f68bbfafb76e78550aeb35d03c1bc445278d8455ad1aee12a0a40e643468a2d26c54fed96d10ef8fe543138203eb6f2a3ed35cdbdd3e4171e545b6465a9185e59570608ec6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hadecd4abd613641c86eec853017b384d5ade67976b3aaff0867ad115dc8e4f4a3837b923a39471cc976868d4590af31d46e52ebffa6d1bb57949c0dc4a22c9248fc49fa66c34a903;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9975ed85dd644de38541864eb5fff4f0672f315781e1f958c4dc9382fc3028f4893db732471021f2d14c8503e7a99e687f63d2296aef83248f1a26bf8ff7d494bfc66c1e96689684;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa88dfc1b5d1f755429117821b1ac7552457c171a85cf93d3cfacf3d6afaac7456d3d06f849c334073c5bbb17e9ee6bc7c8feec697d62a7f8ee17d406e12e0c8f11ec13c8cbce14;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h829fd628a9a78a52cdbe11f72e10a136670bac0bbf02d8282e084fa217589120a546f0d46767e34278f68a0598a916d5172bbe42590f59801880122ecfa772f82348510e80380f5a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6588257085a24d21fabcd2ba553410b632647b7f85a57798e884b7b1e8f32b61467ed8060ce07786b2acd3d9d773f839465f837cbcc92f5d664f0e8c9fbc4f22ddce603685250c34;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcacc42acbc8078bd6bfa075ff83224f67d61552bb46a3a0a1a8fbd977e86a40617a9bc4625743d01fcebe32bd0007de025da062819d5e1b0de3bcd5fc688bfde672feffecf62836f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf10367b5e3ebd105be9ef8e3d1dc210a82adfeaa50b0068ff2f1e7f73951eba8e86f0ded091e7572b0095fd951b2ea251e78c05378bfb6a53bff1292ee5e402ee520c661d649c295;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h40e4b61da4e2f09cfc466dc0a190071555bec44a7cbd932e87b2c76a6bd8348824c90428bfb5a7b7bc8289c3ce33ef66e4a92148f553ded1802d8f5508d817de6379152cb494d538;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h21c9fa0df5111760e97ebee6f21ad85ea3793ffc35190b299fc3debf207247cbf589c9157d5111fd29874c3fd638d70627583fde9a105773d1811ba4decc9ea0b6f9ed1426392013;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1d9a1d1111a4c64a00498643965815c2e2c6f1ead945387700836b9689ef64b5cd2caa679d4a642c00b15f8ffee018ebac89ea6c0b6c51d42c99b1fe6a287eb20f8ddbb52661d8de;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2f36edbbdcffa8f48c258fc5be0521eeb4e88d8864a066efee8a65eb243ea3e9c6f493e053e3d46511f78cca0b053a371bd61ff7087c441dadf082d42d150d93cd8719cdfb8c39a1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h92991dd04ef2361e1c032b52a72e3ce7713dd3294d49fd1cab5f4c376a05e48a30ebbfca435c92f6f8dd62d73b87215efd9f739d9107ad05bf8ee149b7b1d46a856c7b04e9c61c1f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h43a5ba7d54411f952e8b0da6af302897dfd08a7aa3d3a943e55b17da5981c0aad54571be6fdff97f8e765e24f1fa2a5242682ef05006069f2764511347877b7d0f054eb98e652567;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42488636ee7ab2d0a95ac2118d10402d63eb0e6c9507e396dbc833078edbbebd7ae3eb3497b614866d86e14c2947b2f88c09cc9adf10e21c5cc5d3914e634e7a7113d4cc721c53b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb593c3e602aaefb2590072c1fa3eb2c009f6eb23a28093499a2f0b6e03c44590de3db48f640caafd02c46f9200198e97b07530fa7dba8b0b3c0941341524075766816d6d4c2254bf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1458ac0ba15e61c15a1de868c17f32bb37ed69dcec606d34b978e9eec0bc3e28a832d000da2aba0a5d78ffd66267d854a48dd4809c6695d5fd793d118e9dc9dfa724da79af0ded03;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha1aa7fc227d7a95f43af45765ada4fd46b2e82ccf7e9bb9b99f99ae5287a75c741f57b213ec29ba9ad0675a36f412b8a364882217037afff953aa8f52d018e1f99f2c13f43b61714;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h54235357061bd5e3148d3834ffa2600e1c853752cc672646a541d8b005dc716e28c78dc107cbcc35af19968b0a5a254ca2345f499a7f86a88c32d891c45b59ff13fee40d60ccb3eb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h835b049a81f2ce54185a5c3d50e97b90b55ff0ad6fe2bff32fb153e680af6327e5e14a6bc93d61bf8bad6daf37bb742301088479a2a85214b9e15be1049b8bcadebe833034e54e1f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h236def87278cfca1179aa5f7df5cdfe2378fb637d9ac453bc6c4a111e9e1e4f0c4e54d3e8c01513a4a72c7741dd72fcb89ae34f13ca5fe3365e40d8325770416b32b8791a08cd999;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3b0c963534b9ffb042c08a8ce76ecc9bad9acff07eeb89195761e2e614de336d73a4fffd25f3c76d86a99d7912ce43aa340d0dcc865fef18fff63dd19213d253b466464ed582b5ff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf1b14b628415984dd5afbb108a3ef5c81561119c39ed568dabddaddfdf75811d86ac90e967f75b699f64e667028815cc375843d76b00b6edac187f4036955fd57150adba1e62339;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heb5f9e0cf7ca8f7b3c011ebcb2daa01c928971a3c9b407b57a90f6761d61afa62f622d46f21c04bfc56d756bb0d17c5f5dc514aa1e39deff91d2fb19410f0b6d9c9e50ffaadef1b8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hae3b5027230603bd0297b7c3e3d570ea1b46f7cd758c0676d3582405fa2ee1aa62102894c9efbd409fc20968d024984400b0a33289cddd96d22c8f5baf423e3a1699308c3f4421eb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8c451f30f84458683b6e408c2302b323952cb1fad63861fc5eadcd09826c005755115082d30d4e7f9651da5fa9ee8231425d0dde4dca5622860d1aa7d1831e8d622f8192b6fcdd5e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99928b2c5586d8eb84d3f0756e87ef86e937b6c37a92a2974b881dbc0ed8e7505f17ec8939ed687146c32dd955262fe00ffc8b0726e17d645a0ee97bec401a11a5f99613aaca7284;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1262fe0b73c04312e5dd0e4f091b7d8e3a1cf6d65890a0bf7a9b2a8ea3f1a692fcc41be81b77e8c3fd5c2ad8e5d3f510c13f2ea16b7f428299ab6ccd1d660d1f4e0c0cb6f646397c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h44d6d994086257486c0c3663f8db9b04e508a2b9ae2f50382dea7abfc338790704fe4bbcd8106e7aca34e3f8c06de03b27812a9730fe3cb78e6b248ea80389d7e932809ac997affa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdecc1c9dba470287d527a3c408630161ff9346db6db4696f41ff0ab44d8a7437837af2de1bf7eea902bd306d5efce28ccc33345b81a95ae194f5d972cda3e1f927e016c534076601;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5eba95a3ca44ce211e5d67c72ed48c74518e2602b539b909e98ee41b17b6ca2d2a7973f1c83038f0815a5719485f44afc0ea4ca46fc6383c2b07da638e98ed2af3982ea3adad8815;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he6525030f18b924bccf1a10a79dcd77c260b192273e004746a58955b628eaf8f9867592cd2a138bbd3555d0760c6029ba513baa2f573d3e4acc0dee14933c9dbeecb79ebed5bec5d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h232154bb4ac856a3a26de1c8367de58684f1c8696327184d5ffa4eeb38244e10129de70adf08e86bd9cd02e0dbdf48d4623e34454be2625a711e53ebc5d822356104191e3f5c60d2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2ec9815131de1221e577db69ad324bc2d560226d7bb8c337c057733425ef2a68454052c1425f857c2175a9a3a93ef61087e2350407699f76f49f79b2c1cc9aeac33ef8b947ec3d59;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h76b3fb8295da13554e705c281e3dceecbbe7782639256c631a25635bf8db53a741181b2468dae591a8ccf4b9a238fb2ede558c6b0949f14bab486c9dcbc46e40f24de11c292c4806;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h20199539403669dffb31acee5160a7a6da441299a42036ba150b6641bcae431dac7031a40c3ca69c5843245405730e0534ca75a03cd1be7bc4d9b3f23ac71041a1f852155d4d0d2c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5996f1a50d77b3a60ca66a137d875f46c395d48a3432fb6bc15dfe421ac76d017378a71fed0e232811f391065606adf9abbb0d518c51f9112daf4d55289d29d8d247b3dae35b3678;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h878b609db46395a2aac4ce27c88b3c79506391b4cdaa6c1911e207ecb71ba1944d57c7d60d7a067294975df4616a02f3f07f6fc64cc2619758494f54c97e7c08ce01741fc82e967e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h17dacb847dac0cd23ada98abccc400db69a66e16356dd6a48cce8159cb260f1be95a85aa4e566303c7e89be107809fe16abcfc7a8a5db63f3ecb549a597b9ca9e56e71b25c8131fe;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1f25ff51ed99fa282bcb4ad4d8b1512b3eac94d40c825af17ef7b2d3601777f5368e425f50e2c3bd16b58d693280b932ab40b1e0dba81672a9270c91a6da8dab9cb2a38bb92c5c77;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h746f10b7cdf4068f411290835bbc34a474b60ef8094cf203606bce52f4d9b1698b6382ff121c36328d666158e49100be1c3c6637c06fd39f5e1c39ef0ffa6ba6bdf40fd4dfc4da94;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h353cb53083c6b48e99cdb713c1a69a6f592835747bbbf5fd9bdd17321f89198fc15d1dff40389d76041adcbc56f4a1a1aa7894cc8f129425b5235868eab238378a3e2add22a12c02;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9c8cdd29a079834d7d796ac8f8c34c5dae250a10869f7b400e61831c1a7f6dce561a1d49348f13615c7cf744724e5bb63feba78ae8c10ef9e73e665c45a01017465f0c9a5f766a0e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h715acc3f712ff1ed1b1d3c7fd3e6efaa09eedc4abd3772965293b4ba3a6091917543f8b5f25f5585f580ee3c8753e993b3eba4d0027086588b8a88ce58da1f424fe6bda5da3051e3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c9975c2b46fe7ddf79c41bb3b38ee9c05688141c4315a3e0b88ac943114515d485e8b63734c2297bbe3023d51508945ecbe3bc051e321089725fade5b50c6ce75ac4646597d7829;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8beaecf531c518f5adccd84bc2d55fcb19ca7c932f8e984fff2de3d642549ea7e35a461bd08ad5b0e459ee4f214c91e39b0b26f249a6a3d66378092c9c5517ef9e4dbcb06259dee4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbb7ef4140fd52ee6948b3a186257bc94d3dd2bfedc93930b0b1e98b51b20f1e44a49f8c66d27184bd3d61ff8a34be2889f1c83e5525792b96e76e61b85a8d316aab7e6b0a7ebb447;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7a3b7e5997b70a631624c931fedea9bb615cd118b450500c5502e9362e69d3801b73f9f0ca77fed426a925be8f50b635719ea7588ea7897b1dc537eba8c33a8e34d1f497f46120d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h65d275978d58ddee251b15224985e9c509c004928bc6e66b3ca67ba1b374484d62cde16098162c0535f4adbf1eab21bf695062d2c69bfef0f29f171c04f2f0ff549e2b2d74d68076;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcf7ca79ccea8444aa7c21548cabb9ed89bb8338961a69ce659340e657d3734a5e252fbf36670fc437a55e521ee4a2bf0dc25a64b4bf741aba48c63545731ce91c39c2795972713fa;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5027f7ea67c307433ca37e1a1e45e9d7a675bc740dff4a4f070e0dfc0859427abdcdcaa7e190ff3c0063f2aaa5820cb1961d344f14b5330e321527b62af3cfd76ebf5e63f5cd3b9c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h438c15167cba802f1119e0d5274bf63c5600b923984598e2d9b876c1051921ed7c457e1c46d27e567a6d48f6b0959b3170fcef64e12b6822a247c3efc2bad367c9ad57f7b74b9022;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdc989ed8afa05bd21320890e6075ff62bff492429f437ac1ed9784e41f73d586d8f17a5ead5f629f4cf9dec7f01e22f4c6fc74c2d6d973d7a4de99948d8f491cb539c479fbc8943f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2dbe20f32ba74d650dd8df7368f61431a4da047e19cce7370e0da5c1c7b5528f32ec7051316112a0506af13c7f4fbf0224644ef1f13c32a985bbab9377bc857d5ee7218d56c2f3e6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea7db6eb2493724101c53c4bdf33fd751dbade3d3731ee8e93e0c680ed6fa01d2c5d6b384f08fd4f42cb86dbe079489cf4474b7a62fe9022046c3f515bd2eea35c7b64a129d9ff1f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h46b80970e8a6b0101ed922e88b6cbf3de1ebd8855f253b876e39f8c7a4433a098a09a05569e7777e05055cf0c892241cd989099ff14a5d1198dc3c5b71c8d1068d526bd9532cb017;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6845d87ef94219200dd3c9d2689c0dd2c996b278473a52b081168a917ab40b50ebf58cdbc12479a5b40ebbffe099f28d7406cca3939e41aa878e4a31f26d7860b0b1bbc553a8c8b4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2942ce48492dedbd6d278a023f35fa59ee8b7b9014385dd96f0288f354b4b808e56788dc43c576fb9962a8e5aeaf50913d131b2d24a7c75599b524bbe6c7c8efc5f19ba14c632e9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h94708ab2171f6fc48d53bb1e846000f4d308d77c96ec80aba19225440f1e6716af98f2d5e445f951ef60fd85c8e50d215059f3a5c7d5f9e993bd6d66c9dba1686663d327ac92f49d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc6d42a73d498a25386bff215b8a110bde610934634109cce0685a1e81dc3316fe846beff46eec420ed46f6e94ed5e31537cdceb650b05056a50a65a8f415b84435bce7b03a54d3f0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3812763c35640d96f39034e66ff705bfff94b965e4eaf37a52120c6c7b38208598a2a86d9cc2fa1b3f0f5ae0c92649c6c71504abf259b61eb0126838ed1601a18bdd03210638eb09;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h290c10b6e1e33c5a24f6b0732dc3d2012444d17a9f244c4526519d7ac53413e9c9d96c3bdb847240e90397ce37c53c20ac9be51a9903d978a990c6663e05aca9feddd9669f9a9aa4;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9d41eb32cd1c7336b16ad710d525633f280a4555a2c945df087106ca66072bf3edebc315b39df0691cef1b93059bb684ae07c1b2c11235ba29118d619362460ff467225363bd438;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h948978ce6db277b801ab5f20b326b1aad2a922032f484fb61ead69355fe31310bf39df694bdd55ef97b4ec75cfab53183437cf785219cd1f87d7464be621ea67382e797c41e495cf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h859bc6aaa4c617119ab896353286ab9af7f1248a742cf1690b49325a3c3bc3087c263dd76b5374635544f589588faecad4153acf2a44dba63141758a0ce002ac8c96e43579355629;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h74f92f6ca216f200c96b15625422dacb43acf5f04db2ed8014113be557b5dc9d35e42d3b7293b593853de4401ce5832b1faf2d68577bdbe581e0be2addbbc864e0e075672130c916;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9018476e966eb450ee3ec765562e2eb7ae1954b8a9eee9e39e5748c181501c7125c1554a42594689d965dc0f4691d0dd4b843fa69ac7531190d4b9e4039fad870f40afe7f73eb7fc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h53a129e2ccffb0919a046685e0cb400bb320aa033babf9411bfc9bfab9a0e9b84be1bb8443b58d19762170beb6e718a2e1eed86c828774a56e3c76c19cff55b7201fa64255d04391;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca7adb25781d881bf351cea14a52f4ff19b4a960ac099beac4dc5d24ee78ce4b5d9eebfca4ce68e607a17e23252a5c67f9cdd3a0c24fc086768fdc038bfa1d741f51f1939690af03;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd462ef3f75d9d32e648edb1158d3359cca0d960f674466246bf64cff0bdf8e53865c1d89ab7f8896717e0fea7401395492ea90e31698c5d90c32ed44e41a59a4005dc40fe2430f86;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hebe61daa0441a3a7c244a2c6518599d544a7b107597205d768f1aeaf5464973de59d8c2d2d38e98529907f027c07107bb7e22c31ba7a09829dc66c127abeff1a602cd2026688774c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7b4a734226063992ab78c9ef1356523fbbdde2b939acd99ecc2211eb58dd9bf1bacc8308eb38f4936fe83ea5afef0bce6b0b262d0c9534bba0d2a76995e6d58cc61938a5ccf9246a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb63a9ef1bd7a9ae12315e6659db729a9a1fedb6049c45010d6ac8fd1acac338e326d65b5f44a399a102a0d62f56d26d9c5ef07e85adc3fb05e3ea72d090cdf63da8c6b508e9d4e72;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd7c133213b031bf250f96de1d507377028259f1b391c9f04855bedb962bf49a9eb1eb0e2b57302af5a77ea3c1a6a2e927742e2541f377e7b28dba672985f11863d6f4b9eb7a0302c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5d321993d34345aa07aec6205f64726ee37fd257b1f7ff161f0075fd88277d7c48c2ff921b625944833e2af7c89d3d1a0b433602c86a1a52e92a19919ef1232a614b325110c0422a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd8551428c2d1d39798dc977f36e0f276caea327176980b953843a476b6c58517c9e9d78f8398e8d417f8a0a9fca2c72309b791bbda81cee20cea99c0eabccb688fe082d66ad75061;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haf51bf4a0001c6fd424f3beabb2f7cd1fd54cb42a31ac44b76306812d7b789e465e4f0b55d57bed7e424f9d02448aa432707efbd2dc8594a213c8232bef21683accfa1ff36090f0a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5daf704a252db89fb3ca5247cff32207f9785931f54ae8a7a9900c1b3619ba91f0ace764ebc27691088d1ac6d675a8d65fe1f1470197dd3dcb21ce2c36a3be975759724db29384dd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h99833466c8d7553ff64d99a44ef9194dc66c68f0ef17dfcadbdc281b9d84770fe813f39a6296ca737cdea3fb635323766714f3e1edb9b766667a74f51f6ca6049a740cd8ecc36398;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6cf82dfc06c7f8b1c619f3eb239b24ed2e01e24a3e199bfc6bc0027ed385f6848c5d166c05f503308e9e7623255ea809280324208b6a0b30858f476d1877400bdee50922efd226bd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hea34706267fd926ba631d6514737644bc9772df50fc07071eaa78390c822ecee7951863dcaa5d117d02b430e6509697b73a8ec892096ba46eac0c5ac56be4c6cec68f26f700f2fd3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf5cc7713417df0ecb34dde9a7fc711d0e8135181f545652fcdc1e4c6f95c776f777b6b8e0b658d3098c7eb68bd5b31ec8ad4a820d52b4401b1fab5630c28e6fb59ce46818da4b57c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd064e0b10ba784381ef4de63ef934565976620398caf65a38f2a93fe400b25a99db8e31a20268920638642f465f89983e765f2a766e6180a4a4640f99ff7fed9954a67aef9e08ba2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6abaed39d1dc93acb372e16321805e906f104ed403038e37dcee6ca6018848d246be8a81121137c2ce5c77b9542b59df58a790167a79f871b857dcfa9cd404b5ccdcc05542af50d8;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd2ea3d2f15869b13d6e61886724cb555e1bc730d5efbf7a6464ef9027715ae91ff3f243dbd938653035e095a8912ea9bf3f017873dc740f4eff3712568dd724dd0b9f7d504c2bc6c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h175f8c628ec5af5f13aaeec658da31af347f3512a7e11b854306b52221e1b90e2548c7490b0b14651a4c98c669c447230519ead8a9f43df9c33e753d77e6f2afb732295e8600a2a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7cb6ab88007de1f8da8fd4f29ec0238e81cd5170dc5491f542a64f17d67aa5bfac43b9f4035ec028e7f19368b5d3ad28095a31e077c3cf711618f723b83c67b466f3963d3f9180e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6cc15b736a9b1a1310b6bb0c6eb3ce9d71e3634b75596fdba1bf56633d6149750de106cb5f87aeb7348daa0c795ab38d477952863832999233a500bb7b75fc85e655f5ea0369cea0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9958420b42d97a784ffdb079fafe2639a13bbe38beb80bd9a71eca2ef2d1459097e1f14030d9b91486bac57c0d09b687a47e0d54203d130df134108d9b654dd5394047e88819c87;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7cae7b444030c8732a951a4d35d280d9a917c1e21ef18ac7c0f0390b17ce9573c2630dc57456ebcf23ed5e7b83d0c07a782eba8688afc269886e9b8efc4461cc9660866975c50fd1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95bfbc8a9dde2814016fa4b1fbda79dedcca248a63b8fbbb3624e3adf68f2de1dcd57a3da4629001d7823a19b5559946f4d1847f65c0de3aa8d79f216b0286225ec2724191f89d79;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h953976c3ec8f0e53cbeccdbdbee925e66559aa39b148f15d4f3c0dc45c9736d5b852c823f4846fb62427266b81c34a50255b96e7ce126d092e703d86c5b30b4dccd65983559a7d86;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he2d4f8916a235de6ac71c0ad41321b05766fd68ac50fd4878bb9b2b32cfbc074f6d8585371d9e3cea8074ae5078dd4ac01e5b7423abb3bd366f1987771cc019391846d07d0764b63;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9ec5ba7757ed5d5ebf85cc830ec1c78a1f08cbe59c8bf897eda27db7b351eac2fa98c80ebec1591ae1815bde6121dee0fa208e95384e0a9db9b65f3de229fde393bcd750212802d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8818dc527d349e70a665350d479d1a6b072eb1562862c86fc77f75c0931e57e9b0e39d73739e900520fb78bf38553009c06eaaf4529e2f9e51fdb3986ca2d429ff21211fb3aa9237;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e44925d43e326c2b6696679b40e672eb5de5a1906e9247c536b3f6896bfc9cd7b2e617a83b2521060997cc61483d7801b6e6ee58e3817d86922f574a2b1758d0d9cbf2e58c8e9ba;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b65162cad493c494b9e4d2ee063b37301f36362837ed9504bd15b9acff4d1a0d1836c455197bfa55fd1bb32fdca2c0f9f22caba4ee961a14d65a456ceeb309e9251f463756b918b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3f6680f6ffc657163522f9cb98761ad5f7828d7d946f5b1d86a5e42cd5178128f68b5bd1876aeb97af8a116cc975f5ac99697f9916ede6739f1796e5fdb792591144be9a4980d962;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hde0250b8aecf65ac7b0f2c84c7e43d187997c40477f4e3c500bd447d398cf12f82dbd36efcd8e2c76e55c02638bd76b2283596af75898f486906d9d3b383c7860ed40f8e351852c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he009e64027de538796b15558e1f4d61490f6d070074365ebbbc00663a6054dc2ea17cef41c319be7f0e3e7525b646a224ff4b55447f39b5f15b4f8273e2b4897bcbcc36ba3c9dc11;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8d256145b52a7c628b67f69732fbadd379bd8502e0ce05b40c83f687f815298b3ab67b93ade1f77c444df6be794ae48524562c59b5ddebfade3e63a80996a7af189de9c3a872cfcd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h829ba12e4d7d4d8ba9080c74b87fd956b8cf68c09ddc70bd585057ea2ecdbbf8acefaafd74ec7828ee30939ff223a31127a8895e9d1a692c62bf3446855d2fd9f1993bc4817f39d3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfd964faaf11aa58a4886db41f1ea05d5a6e220fe41a5d8f96b42df9038fab61516e182a6053640f56ca83cfbb247afc7bd5a9628b40b4d7c2b82c916f91b76deec96aa1acfc2567c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h68e536f142ad02fb4762b96d512550d1e8c7803c06803e902130a013c36d66b5462434b6c6a42a76848994748bf6e60bf858c9c0b88af60fa74c7c560d981327723e5d028c6b4c15;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h3fd763c6772b504f970e106c6377841abce3a42ac61ad64f45964ad54ca105380caa352892bb8becbf1632da2b77b42b90a8ac45014367bbc8f9530ed2dcda773dd4b8df6c235a96;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h528be02ab61b47e421f061ff8ad8477b21e367ded497325644fdce2221e4b59a81dedf41baea7ec735d4be68d4550347fd80be8184e551c3dc1f297f9a0d880b6bbd70826cf3ec3e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4b043db5709fa2e169ba48620c095e5a7178e392a8ebadda2c1071a82a7396411f8a230471d2a0b7328adea2b519f5daf3bed44b996310303b69fc8dfa55666838c3bd8ff8f8fd6b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h341eebbd47fc639b59287b729e7bbbb736bcba1d306de0d0ddbb8a517ab2e18fe51cecd0578145854b5adc9e98bf169d3d5b764b73b071ddb0e2eca7a561fb7833d87b54949ec4e9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he7a848588c7f6f6de43316826ac611aa3e63dfa7bf2d044a43b6c40f201698bb17c5317e48863f2391c5cf91cc9ceb48b1427393fcec87d8a3d8c30657854ad16bdb6f774dcc38da;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4c8ac49a40a89e4ce731fa6220d09ea1186291f31718f446da96aaec198fa7ef8d1196285b4d7f49f073d5ef993bc5b566f6d2a85c23431ab365bdb0ec6d50c3562424d7e7ad8fb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b37bc3c957fbfb3d8ea96d5dc737c266774c37301d39745fd0d463350082fd9f8feded2d90a958f9990f1d6c282f3aa3bd490c2589de937f6bf201c9d32a33ab5f9d7416f6c006a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcadb027d5dd15411db919ff2473bcd42960130abd08024a1de091a8f584c0483bbc89369e3e621183e614e6c535582bbcc536eda6fe756bdc9473693781998afbaa58924d4fb1b4c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h83864ed2e7e4a21f4e22a33f0ef2a01402d8ec16b99e1c0416b12d4716f38f33cb81b59c3dc689dd9a54ad4c0e38354ba8b6e6bd980752c1cdd1ab33b4a76e328b0943933bb635e2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h56ca82ac2642e2fc01595f38c6ac204390f35a27903e8c48b863a7e89b95acc0450dfce95f1045ed8f3351fbe5ed66dbc339f88ab00c90810811c1283e0f59371f7c7626beeb519b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb1077681fc7586cbaeddb5a1295c3ae2028727c137c4102dc0064a711150e99563814360bc8f23796ef2e9408a3e1d9f2f5bb20d14bef8ca9653233216396f44d1bf167860b86cb0;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6e67d609231528b58ee151ecf0409ee0b4408a77cadc1eab3450f19ea60963324fb2eff440e20b358da1cdab801635ee2c73b2594569efe668f61219eb7572e700e1d6e59cc7aba5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5b485ecb0a07fb163d43fad494f71a97887f0e3c22b95262681769a06a388066ab2926b1fb81e756321048531c96e59d00ce2ba6942b5f945cdc4b55ddd5721fdd0a654d82e14237;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha821168941414a7d4354c540b3c10d57158c50dee5ffdcb2706255c5732b3195c9d9decf1207192d87db057b61505335d2787ac03227ea577ed398bb23a98ae728ce07a1a5751cca;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc9199377753c4029488f99c3ffc638eb42d8909c77faeff15c10bb29db83ff44d65657fc6ee9340ad1cc32a9d90e4ad3811293a96bd8aec0aec925e432169cc1cc574453755c1405;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h210ba23192d360067c48fe4522c4d728ef1665bd36424140a550d204c31b6695320a07ae8598ef68df75242c6967e766eb707efdd719afeaca58e55ba1eadce4ba2805c996b26a29;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb06f91bb996e806aa1e7a1db0b5122e300696e4a551e3b2d89bd23b14ec33f4acf7618374935ff1fb2ac88e8e53ce4af1c73e774958cda193ce054d82690d54fa08e9748bdc1997d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hee1af7205dd940a5226303623dd2218a4668e27aae255e9981eeafcc67a873bc697f140d4c076874378e19d3a5b4f40ab01665c06a980a0f9245cfca879e014c7a5b3799c3324b52;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h38ae55159b1fcf956204d1f83628f43987009be198f7f4261bd9b4ffa71e60aa89c52da0e8ed871e7aa5a1acaa49cf3fdbe526e2e60dc463fba1b429bd6f486dd884506c95695d95;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb7f14b01947cd9c8f6228124e6bc7be1a607db7602fc5e7a7d30905f48d0d341ded6a9a4b428650c4620784dac8fc5036a7a91f86f49c28d9b49eb67144b85f9cd987620a0f47b17;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hf5448c48640e2af1b27764cee9c56785810e9141f205ad1d564ed7a7851ac3df84dae96d4a1e0cd296d9cac28bc777ad3d989eea8a38327adab267578277e1c4282a65b5dd3a9aa9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he175dcfacab0041e62a85f3e6faa2974aea3afcae7144044cb7e1ffe60f374918e9ef400840b058777cdc04ee9f96c5a456d17b6547e64e290d8fe9a3ae4c8dc8e72ebad20598c26;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hb9388dacff7b5b3391c1cbf177e1ebe72c412bbd575df7158db5f520e6d1ef59d080fc05e7016229edf2e9d91510a2f09dddc92a65be2242f7eafa104df3fd27926b601c86517037;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h95db81409c639f2e0afee5169ea86634e8c0b6d9f9f1e2cb026c4743c497fdca002f99847013e817ed00e545f8de18d391f6cb64e872dd2a9dcea4a3f7cf3ef7a279c2a6786f39af;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd2790501a1ef7e2a3bd8cfcc5d7e4ec5ae66b7e2cb2fa3f58d4fc6470937ca19ef9fd82096584e982b6e44a0ba9303f7bf06d38f4738d56293d2fad03ec4e01f15d482aa2aa2c10a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8bf28c3c0b415cf06462c5725737337743765deefef0e2490f7b5ccf6222f240de2fbc2b2e777a33b165cd7e9bccf67bc966fc28eb94316822192e958692b7eadf4b2baf059b7fd7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9e3bef769fcb78855ff27b46141070d28d7be8e3b7dcbfd92ec2106e77cddc72e4d9597ff0698ed883de82d40a6106c6812ff21c1ef3b797722a44facefd082a2d0e8289374a1519;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h42b9a7553fd0abd11f316a577320dc3a26f415f46e7361cbae080603a5b61acad2ad1c0fccb44b6721c03667fe9725b74fad8192b8b37399c3963751cd7163f107adcee22615548f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed16abb009e45264604184c700ba188844eb859c46ecd7f43925f686cb4413df4478e1d474c92f682103bf28b3cfab4bd2c1627cb573222c3d9f236da2fc7a8cb9ec6bd643c197bc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5f8ee2bdc7f44ce08c97da79b9c25dcecc10b1e00a8d7f1a43e6bf96ef9a02f2c4bc0b7c75e633670a6425f40eb4248a25af2176a98c6aa32cba3081fd8f22040235f26ff8a785dc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h894de4a53840c67fa0e19f6de1cd618c806f30cb0a1585d12ba1ed08b749db2925a7b53e95ffdb640843374d2aa6127abcb6339377ce19e0f6bb4c2329c9b875aca8b8c53665e48;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6b6743f5113b714e242cba2cdcdbc46c4136b94aca9ad6f1bce5c2f13869585934346b3191f7153ac56172ede7f1f38730c02eb7a5ffcc0c4578dd694a3d099f7c8f444c87b4202e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hca1f800ae986d5ec9a1283b501be96508763bdf710f6415969958d200abe32fd654f3ea7dac991da83ffbb95c600d9034d788edf6f077a5820fab8e457e10b9eb94d1f96fe36a718;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h8518e54f3e9b0cf9adc23dda673f65629838a14942d97501cce861e048509f0f8254bab0015b0d82b25f8e1269ccecfe5d5de7f45e84066c26676288f5b61a5fcea454f77b4ec3ea;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h27ec1bb73d4f7f620845c4e66bffcc1e45d16f3cddbc9a17fe6864cd1b8fc8477abc9f0788105413ecceb73f19ede99308d82d6d5c25455cf4264dbb6bc10c98e7d969fbd37b4d83;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa1adac6acd94d04d2e8228e1ba5c9f45f36c4ea93d1152581aab70ce7ffb5b1e2fbb44379d4e83c26b3267280efdc53b8379d42aaca8e8beb37061591e70619141e1716c3fb4a3e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2681b6cf9544e799f6d8d9b3d7f324fa4632328742d87ffdeb7c425020ab66b1ddbca07e9f2b666421e1197885378006da45472fc981cc7dede8dbf58e11beaaa53bdefbfd2cec91;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcb68d35a30b3d6c318f44665132b8f2a4dafceeb84856ab6a57c5e8baa522edae5d0b586171bca33b645b74f2fabf749c76fd9b3ac649a9c2b0e4c2ecd0a882eda3d62e0d892ddbc;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hff9937f3e3584f3d8a3cd32bee0d5c287dec946114aa77095a8a59776de9d7500ccacd82c92529f8a1e3f3239af71a702b2e1993c1a98d94400644c0b4eea7bce44e08114d19bf71;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd2596fd4d46e60d521dd300726b790953c72a45030c275acae94d7cfb134fd71d848749d2ef452352f772b6d1352fff78825cc001c2c8b8078d090700255b1ca4455d7fd3aa1cff;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1ab5e51d574fc5f6bf9e557015b85da2910f5b2ec82b585b78859a8c87f4a619d89ab03e83fb881fde59021c3f6ea5f57627e068ab7c9f21fba371454464e4f89bb819ff4ab2dc99;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haa52ce17f19a43ed2a5370a64396c90cc9cc37ff9df376399136893e4befaed38bf77232ad1bacd351aa8004b6857ec30bcea89e432a5896b2c7f2d781a4a5ad909c47e4d7b95e8c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha52929bfabda93f405bffd4b4418f0f3473b1d13cc7e95cd5bfc7a2cea37c4e95cadf848a9b9fb3e85a26d54d977fc901ac647404cf802ba5f4449d6ee1c21aadc77ac449b4c446f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha5ba232181c78a45e5efc7a0a7ed7f198dc737af5ee22820423b70872b2d93c9a7c5f498ca2388b329591e2c13d9843944ce3f1c1f0ae0a01f462b5050444dc2775ce6a011609109;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h386bdcf165a073c5ce9b128e1c7ed143c7030351f91bb8126dcdb2fb092c684d8d450ca8e1d5a422a87b094146974eb0a9835e48bc916498f0880268bb7dd5c202a71048c371da66;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hed87c666b0fa535a0b92f63cf97d1269998017bbb6700efe2b43cb8fd328a98637b4dc4c218ead89f71eb6796b2518075458f5fac651c09e89b2a957beaa1826acccc623e2c22ef2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4eaa19f57cf60e100f564c3ed47152356ecbc2b207468d3eeae4d2df220ce8a4454121878ef5724c3b141e55ff83f602532fe4774e03e1268c2a7dde66098e327b769dc4f6b4b6c2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h28ac67ff9a09aae51d75e1e0d82244bf25506056e6d6656c9084873ad18c52cc5437346ab49b95ae143d55af5a2322c4fa0eb824ed17f0b195d6164e7b494060736e486950c76567;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1cad1e4450af82803643d9c4699959612f51416823adb8d8ce6768e7a9e501e0fd9de34f8f6384253a70843a3022e6c0f1350e16d9be6600b2e98e845119b3b85b6dfc80013cb108;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hd58395785da5e83246445df743cc8dbf81909d3ee502bcad8bd3adbf0f8bff2bcf94814217a511539214dfc90a2dace07d618b684d0507c38766adf4faaa7db32afa3a95eeab8ac2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h85e77d7d7bbe843ab3ab75bf4131cbd1ea98a714f5a717dc85a5eec175e50e30965bf5a509fc6a818fc84e969cb1c70d829aaa9556806a72983c2b65c15b16520ab4ae4436cb6db2;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4738fd33095f77c019f97f3cb9bf5d9b2cad45cfc1c314da8ee25128578ddacf971d7ec5aa715001900bbe7a7d6b7c305903f439584b9adc2f1b46d164a768004acdb2afc5ff0b1a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha229868199b23400ef3c63f643aaf1d72a0f61a064fe5f6fb6fe282f8ace6835d379596e34d9d5cc147588dae3720589469d9ec0bf84082953f157275b249947197eb296ea1b97b7;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5c7fec0a92a4ffe77444595289c995d2339f1c7043f7132fa138a7c46e713a49f1698fef0364385f5aafbc107829990d25d9e60444ccdcf0c8b91bb5921bf189ff341c51f9b71483;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha2facb9e8a467669057aed057e4a3f4ddc70ba902b8d96471dfb63f6bbdc1c4c4dd6617cd136b3a8723e46df646324ba0f0c0218e3e4c33aa5ef105fa5f686889ca788046956e6b5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1b94643ed61f81d1be66724a673475f92bdefe213eb3a6df396b8ccd58d0e041cec76172e30c589140e4edfc202e212af426c26e0efc8a8faaadb09a1c83f10065f96c9b69b1353b;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbad51e2436e2c06a4fb825557b318090adda940d4cb2969d701f04c36f6fe28ac775208001d88efc5c82a91aeb6345e0a3023732bb1a5b54a325dcaffb562205609e964ecd4c77eb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1591e0ce3dba4b6bc0bba109a1101bba8f47b5e149fe2ad5998c30ef93f5c6f1184f0c8fd085de17c2b441a0f702ee4a4fa25f163e5c4d091196071123ba380771d3f4edf4ef55f6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h433da03c8eef5207eef77762396bef1c361b9f3755f52d26255f68990a10c69b87504bc824a6a40f9495713a613c2c5afa138db9a5e206f36d4f1360c68bff107b4948cd5015d43a;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hdd5f1b946d27e1cc0d50bb505ecfd081f0087cdbca43f8f01de0dff05389629a3e94fa7160737c080bc61002f15d95d397327d066f32a921200403199b184c1f2c64388e41cd8514;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4facba5fcb94a2b625fd898178b449fb9708daf39b91f7212c58e50623c79a1d917dc37c04f233e16927e9d9b24cbcda51c8d47961ae3b29029837204ae567b5f70d9b354adf1654;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h87808ee8065dec6a98394e431669dd9e0fc7b3eaf760f696c1ee8333eccc95fb670b19acca59b30cac08e6c26f419dfbb943b3cbdf7b4f3625c162dd7de202028f54e6d47c061c6c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h1bdb4aa2f2a1a8fa8408f25856e33bdb7b32461f339a202a5b92543a31f51d1b92ce6d29b79fd1a1670e3c9c0f8fa76ea47143809fc929487d8bd5a656978b7a1da81ad4da8c6877;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2c1242c914c7eb807529706b4face3d34e4c3c7d52dc2decfbe8df60989ac62d557db80f6851dc76ff3c8455598b35803b3077d40e692cdc9beb0d9f2eb72382b60fab85fa86ca4e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h55a32cb0ad50b9afd062663762aed76b98eb2a841e7fe33eabd15807a6d88964f81b4d358d7c8c05b847264cd6d447ff0b7117b2641845424fdb1a1b42b03a36abbbf6c6de4b0cd3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h35ea98cc03bebe430f1d52b095cfeffae858406c851f31af8e9f7bec09d151b84bb5e962b7cf6346a9b06b0b93c112efda8f708fa5c73c5ed7cc50c6a11e33965d5082fae84a4a35;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hcab76f6160759a997ddc25394bf67d0a9c663328088c5307fcfe2d071d457395b708b4cae16573d5e84a670baf41ae43725f1bdf66b8f164411e8656f5d4702240daa620b7c0bf51;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hbf4920ca36b1a1364feec25a3dc89c6ddd1b4ae08b4767132e8e2ccb49ddc917df652f55875ea88477e412e54e7ddc488cfe2e9b6f19e23a100f2ed42f4c8ce5ce67164fc68e664;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'haee361d3c3276852a8ed22f78571630c13182bfb32a38337c874f9e78494032e604f43a8906d1641a323439c98bc01297f35397877bc3a308a9f4dfbeaa24fb00d92053f81c7455d;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h41e6d90b52cda83e6c2aaac90d713c2e54c212cd4b1c2d1fb44c1414db071fccf55f000d90016b31d29a940cd2275e99b18e001087855d4d6c10a36121529d92a18abe3e27623973;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'he887f9d3214041d8f48de759a3def59107a1b2a1ba6e321e91c86f4273b5932753da49b92aecd2f4444940f96075a62ddd993b5ad024d511617fcd1e9ee0bb7af62c5919759d6b3;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h6c31be7c9b608c3cbd8fe5dd947f467c909aea656a42f9c10ae7ea859215c280b65de2964c5696cf4ad499ffd206c823626e399bfca0aa5ab4f963733c871271a5b3e58e10c9b4a6;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha8ed4cdb1effa39b061d188a9969d4f1be8b57631dd79e0ff85a45340f32a3e13542a2cca2084be6145412e0e3a622388c252940b5012a7a017bbc302d076bcc8a9c01cc93486889;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h5ff799204a8efc6a81590f303af0d609f4116b1826c9fce2a818951ad66d67e386a87bd6bfd49a586e395dfa4020f6c2a884f871becddbb0e21254baab42d270ecebce095c395233;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h100bf720b5ae8b61f4eced996fe76bd3648654c946568433f470dee472b7223d00290333fe2395524d207d99686b8a3fb884ff981bdddc9f6bef45054454e8a0bd16a31b9f4e6caf;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'heae5f245010ee0ff14abd314a09d8583511b5e8ab2fbe21eafe832ccf8d3f277a81092452e0ebf54652a01434732759974d701e788a1b2b4b7dbdc1a9cf56c62e192298fb0ebb6cb;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h913952b5530da38bce759ac6658570ef1065ee72b407aeee31fd56b48f717ed19b68cd49c8fd687af7612f8953b6cc8e30f01dffc313caea5ab6fa06ecaf211b122ebf1eba7e7db5;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b688d84b2054e4c2cb7b04887fc8d9f4d72ea83a7fc2d727a9df02db4d8845df0b8b28eca5a6c6f30e0502d44ec1ea83a37b6a7dde5b0deaea493d81879f83a54788704c7498c3f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h9d0bc08bf069ceea74e40d37d4c425f3c522b78266b9d091a39db935f47630980da341c520af506334c61bbaff189f97250003a4d773bccd48c6f8afb4c9086ac6d01b87a029c28c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7c2b67369f1364e84f738aaec465bf660adbff16b40014d06ce514dce34afdbd9941578336ebe7e68185ebb26261045dbb1fa406449f2485c30d8f835e5a93714ac79ecdba0ad0f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2b04ce543d758340e48b7a54a0e9dd27bab5ba3fdb7ad4b010fb457ad6d5e776c9e25c7ed63362f86bb5f1a6d0e263747fe9a6f437790dce56bf631480c6f170f4b9c07a37aec12f;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hfa50f306d71dce66a126f05c5f822cdf24b8046503eeb12f316d1c2b100a69288419567bccb73648aab68a370c189e839da2c19534103f2e0869abcbd579f88a87e4c76311e5d3b1;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ddc3e46499bd2f8ce150269df734b89961b5da8802a431d69755f355a5a8df30929549ae234cc5eac29b4ac1625822a4b7744993c5b309469317f8dfc8a0a9948b1cd2f5e73bcd;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h7be534c684ba33b0f1b685e222c0ae9a32283201ca674f8e368f5ba6603c087e366035284e9b7fc05aeb2c731b9a513deff8b85de36430d25def14582038c326434c690e5a819a97;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'ha41d6221991c4a4cd11e52ee56a46c5ad130b9f094af4faf17b46c4c2097d3d6ae404e5635d2feb1c472e8a357273789d331ab92986acdef2dbc5eae7f29341974fb76f7ee36e563;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h73856de8981f7dedc1655fe945348956e6b686acd18673f9c0ed270117ca3f37939b9ee82ac3483f27026b30319bc3b9271fc9c6e0bfe50cc87546c29743b9640cd5a196e1b2004e;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'hc16956bb5478489842a459ba526ad8644cab9d3aa7e1d4b8476387edcd6d3e2a7e73fd9931fcd8881a47a6a109fca898310132142c76416d7c9228197ad541433d93cec353c3bb8c;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h4ab2dbdecd7d84ad98b210261643fa3c07cdbc52604ff145fea0bde9e2c81997754eb54e5ce32e7831d89736db3839095533a31ddf0cd6296fe82e0975a039d0267946c53f0ab4b9;
        #1
        {src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 576'h2e0dc6295f135f7d819468871b5dee0cd474602b31dead590be95f76bcae3d78139a0b57e8a8ce1ce10f7b59d5515fd6e8d8e564ca34ff3c69f0dad42f56a7a45f2010671c53d95b;
        #1
        $finish();
    end
endmodule
