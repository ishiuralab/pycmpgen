module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [23:0] src25;
    reg [22:0] src26;
    reg [21:0] src27;
    reg [20:0] src28;
    reg [19:0] src29;
    reg [18:0] src30;
    reg [17:0] src31;
    reg [16:0] src32;
    reg [15:0] src33;
    reg [14:0] src34;
    reg [13:0] src35;
    reg [12:0] src36;
    reg [11:0] src37;
    reg [10:0] src38;
    reg [9:0] src39;
    reg [8:0] src40;
    reg [7:0] src41;
    reg [6:0] src42;
    reg [5:0] src43;
    reg [4:0] src44;
    reg [3:0] src45;
    reg [2:0] src46;
    reg [1:0] src47;
    reg [0:0] src48;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [49:0] srcsum;
    wire [49:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3])<<45) + ((src46[0] + src46[1] + src46[2])<<46) + ((src47[0] + src47[1])<<47) + ((src48[0])<<48);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7069b2a9f3a50b60bb84f628b50236d18ce813889ac3b15c74362885d7cec96a327f73bf4383870c132e01a5a04d11a30b9fe7eb526077114c58a303df812ac6bd664ea9b95cf5655a484c176f9c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12c236f5b3832d05b663a912776c4eead1cae46c2601c344e783c53de11edce52695e536d619e511d9c5ff26b7d6d90421db4714aec418cfd058952b43efd05ffe8ee9167fe69bf91be47b26aeebd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb49fb8db5f4b69157eb7775b60945a8a2d6a4906abb143b057e87e2f38c147c50a2fd09850fb48c43d360e26e0c6960f72dcf8d109fd1d0677f3de5c36bb78436599087c0916f9e1cca8a8413388;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13ee6303103bd2dc5e70735b203a32513220685e3daefcc6283b8918e4b23fad1cb95be400ed6220d41a4a0dcfc113636ac58b6515dc02ac9d6e42a632895abc9de27cf31d7307b2187ef31bc75c5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1927080fba3dbe006a65040422bb83504734c356e406ed5ab4b7f0aa2c468ab4f47a30ce9018b3f3b03790e4553badc59871e62aa95415763979d99b459a57b4c7074c61709d3ad28f97bf9d14ffb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd03e54694f47732291cee8cbe33ae2d3eda6839f4c92038b70aa8c2d3e17340d49048badc2337cecdd28d351c55449f58fd0988017d790fe9fb56357b72eaf87e68a3fde6655c0a292053504fc8d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11d351cfaf2cc3113d64823606d8f469bddc10556a3f6d81cb1442b9fb9f3aa00a3198388e55c891552b789e249d6e77de323f26ec4d7e0c958a6727a855b7f0ae785c4fc06e7ce4b5a5d5cbcc7fe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h168ec3fb67b5efd86ac8f5d04009cfc97fcc7737f3541b36a0b9ed2cd473c5430ae436ce674c7cd2683b0c5c5471800c38d5295a06baef59e14e74bc73c7366cedf8e816fd5534b58fe4f34baf2f3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc349ae33d4a80a208b48ab648ca7e21334d1d799f4424b770eeb0d145956ba47ad0c31c919ba0629d39dc4361fa5d04ca13a765aa6fa2b5ed1bd495c079f9c2ce1d59c682a25e3250d84b71d17de;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f9912ce25c80a8091c46e2945774b9b73b5603cef054e2187b344eec7c6bfd4536db0e92779420c4106887f77f14e2005639afe21c33100cebf9bfedc16716cb417d4b56da0652ef4a2b600c948c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcc2f3096d655faf76fccac84465e18f8b1fde72de046e58f8636e3c4e065e57fa9d69f86d21dcc96ac966e944ccaec7096a05bcd5079ece44061d140976f443d7e9f094f22a4244205cfed196257;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a0cefcde2e1ef5464f86315f19c05c2fc4fcff8402146882eb64a662d755cd4d432f04cce945a375f98eb303be58da324145823119869c149ab9b74795c44f24eaa42022eb8ca8069094c5a464be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b6ac283415f74e113de0ac8270eae5d2e7616e97f8427abeeea44296767bfc60e2dba52f64f5313d8c3253cd18fb5225ea6ada1b7b1516589f75778d283b235919ef61f550aefd4af30191881e8f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13540f5a73b03fee1ca8d0b093138b2698237beeb97cc6e6387dc63cddee8d6f257c13e5dcf4b553bcfa600b8ab66b2f96e8387dd9f60edaeb687eb2ab77a6dc0400f59ba15ae353c4b5a95d23fa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17bfd5b19abf0b6234240937e7e23a449387a4ab98ac257d7b3439d940359d4646112b5183fd2fc5ede1eb0c0e31672bb70a28728edfffc0479520b2750c8f4e72edfd18af70cf1ea17a46f2b0a86;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14fe6f742fd780a8d648c24df4db775424eeb126797aa7079df1203dbcfa6b985144f3f0af81815c71c4f8a581c4244659ad593b316388985470c22dd90a6b671c6c75a584cf8b853b7dd783490d6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha31022b4846dbd25eafa371a4e2dd900581762bbe4892ff410ba4c6617400ccf35b8443def444b8252a13769c7090140261b92137dbca69b2a7e6ea07e5d0baa850efad47de299d8eec5258c3cc3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h43f0b97fa0e8522a65d72326e4ffc604139b908fecaddc8f28420dcfeb6250d4fc42b48998abd4c555382d5a34fa75c8caf8b211b0e90cb59f68fa9dadf94cf91b17d828e7ba5c168204ed373777;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e8b751b78b8c40a0e204344bd57c5c5113080d98599661ea59825c570bcd06207542d21f821f3e31c667952986ddbd292ea032446dbd17b072221ae0737de6281e3546d65243fa10b435141ff7b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18e7c2bda2de201f74e33cbdc8280e6edaccd13106351bd4c90f6b7b66c11e88f6e845c8d1e321516c9d9a55961b7b13b48886a9681068632deed5275f513cd1821de6e482b679c7e3da31eefd5f9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h610c90904fe7c5f0c989649aea0ab9dc7fe6df2d96ce110cf484a87c61cb77df7c0269893cf3d044b6c09cab1adb08ed9749eb30e39ee587961622edebb726036fcf4b40b897d45dd9fe1e7cfcc8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd77df80c1a6b79a57720e49dba53f91e86bab75c4ca32d7461d87b602567e5b721a97beaf8ec69588b440b536b7f97c4e4cefb2a6fec0242e1444e0cec5aaa785c2c0f16692c1d1881fb01424d5d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17ddd9f39ef4b394aa54b166b975647e777cf2ba971ffde5cd953895e43885a08f46da10218d6f5a6feecd937cd7c16ae51b08b52dc8f8be16e4e0cbb62464f023cc1b3db0c8f4a7901b69d9a0c02;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8ce68016f7c836735001e9cb906f9b25a89973d351650382cec3c43f9b6b9fc30f4c7ce4b61da7c14dbbb043df270dbc2254023441c780b39fa77ad1ba3c66c282f3813349e0c73abde5e886a6e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1167fb74f7f320d288101fdb325ad3564a609e9aa9e1476edf2f1566c57c9f8ac6a13e5aab17045c6255a3b15e9516612e5d428abf6590bdf1330519cf1a6638728438c72f7cd84f26f86f1a309d8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfe98353386fdf922f9e3e5b8cd0ba5056817922cc56e8c51c0ad0d68398e77765cd5e2330d397d7faa09160eabed7b008d8848b053900689ad653fc7732df9ab2f8e4352c9fafef8d96745016ba5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7195b31cea6bd7f8ab27fd2804b2d029c1a29b6cfaa968fb99afe8500d903b9076030ac09a957498f40a0a74ed8c949f54752b093ed8646d058a12f8bd8e17755c4ca2e50c5594e28af32514aefc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c0489f99daea78c30f82bfa9dee47c546dec10525d65ad5b1f11f463b27f5603e33ed76253b1a0766dcd645840db43c069b805686d09db49e5bde3ed4fcb8c0063a2fac8d45f8b3ee7ca7b83a09d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1269079dcd9a9d02b3ae039308b60d95cae1fb724193a78c621bdbbc1bffbabdc7e342ceb9e6fb2e0c564bf55bc69f9db65be4d130ad82c9846be8519d7ff6e09224fed936716a0ae4ab07bc6a168;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16d3ecbfc02ca9fc1796fdb1af4a0cfaf22c6795eea776f0a9b481b9f0fc6a4854adcc92e60e5f5d95cf822d6568ea865d9e311772004f00a2041300d4d66c5a6c9d56fb836850778ef83f7275bdb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d7f413d9791a359895c36e8655a844063996d3cc5ec93e223a8ca7d54d74765ffafb98d53bccc1b72754ca1f741e2af71a7c4c992ce3824ef17a123a8f20c97738fbd707f97db2c7b1023ce889e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14b102a4f11e5162e7f66fc4ae38df9c3325ddca1e3fe360da094a8841d1d08be2a741b3d7d34a8a85bea57a27f8ab2040d44e600cb5d94c70e96eeb346893d17efc81c251f8f414ee8577c3e6663;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14eafcb6ed6b7db6d1b98645458f1974671ed090cbfcd6e7d3dc832f3dc64691800a452394583ab8187124ca6432c8c6c2baa01faf17c0f76421635cc840e435f2892ec7aa561ad417ddbef8bc4e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfc750cb140cfcc85d147ee4127ec6aa982a8cf10ee40bbc4a0a8815749bbf92db33e2c5b3917c652dd6f2e9ecddbd26421c6c644231fa5682fd0529afe74eeda86ee95d65fac858bcd48557db58b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7e8e92de49dd41444db3704502cd7aaaf4bac205dd61c8459c8f06078d5454790fb1d8d964e273d6cf6fd88b668b3637361bf35f538983b47acd0e063ba36872b1ad37166444df6ca05e37974045;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h172074c87f18cf0e395f2767016c8a1f729c7f2d35bc2dd40d1fc68ef80a7050a5731820d53d675beff618f16879210c20f85afc14968e255937873033ae1886142a7a3b227e8411406ac48fc0909;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha53aad8393914b4b08eba2d2efe5acd3444c11b57c8c532fed5d13ce397cc87ba5309ce332b0b58f5693278bd9ba05634a35ccd746ca79e276ab747b863947f4a8efea72767152a44de0221ceb06;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h31f6690e65dbc77fac6723d9ac81026e8847e3555ea8eb433ac7957a2c26ee355788ca606251f4bd89a6ef318002c9d823a76224d7b1ba758b01f1ef811971464451de330fe065a7a4fb1eb88d4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc105e093e33b18bf206f8d63e0c9498b2ada3645fbdb11421afd0ef8804a281afe3ef2205321de1b4ef0dbb9c086043497b59af8ab6e06fd1e735bb30fb97aeac62ea41cbf73776589c7e9aeea1b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13ce835840fdd31acee58008e990d9c7e4c0c78a2edd74afbbeefcbb91305caf5ba7afb11acf00ec43cd6da314cd60b57fa3f31530094ca9adf2c3b22742e5ee28e026e6197fd87800a41ff76675c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbd2d953c75ee3bd30791829a4b3e51ba383c8925fc2f42d787e48b50b76deb13487b2e07816c5d752b67b0aa1d1d354bba1244687062cdd0c9aec013c2148b9926ad5fce23979d81b042a776bae2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17377d6dbc800d7c955438fb0ee9cf95a305123988c09cdb4a2481ae84073c35769dc2db0820c1242915ba932808e02760d3750a21e2d7a5f74ac52c75f24f0896f5510255297acfb509c12088867;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7644de2e99f257534641752d439a4e045172e95acc3ac506cf91e3a6c67a86b414bfa1600412ee754cb488d12d53a094c728a6e535df44a16156f4bfc5fb7191fc642273ab3775580ca242ca05fa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1908fd610e7f5c519d3a18c3fd1c6e40f23828361aa028493dadcc4227e18fc7e309e55e77d0b037f65e5f3c71b3cc5d0f116516f85a1d7f0d75f5cbc285a5e7e6c11466b99e0c71c1b0bef973209;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1728a319c51b2ed1b0cc1c70cbbc4ada620deadf93b902af4edb1aaefb6e4ec828c35c8d0d82dbb4e217c1bb805f704df6966a72a7cedffce6cd900ffef68cc81065bfcd488988986ea6836302528;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13724717ab2b9009c4bfa6d8e9d272bf11970fcbdec012d9058d89431441c316f6a5103a8523fdde049d2b177362e4d4a2883840a88eaf8df08df2c64e9b1dc998cb9c101dabe5b7ba76b52232f22;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aabe0b17d19f237cc469a3e9a2cff804c63459f175c5391cebfd74f473f33b093b98ffcda0c05a77a25f76eacd068b9497a4b30952b2e7744715a0c3d7349956ec93ab36cb2a64b084357afbfd0d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aa967515da00d8b525200c1ed2c5c82ce1008b6af826446711f02037d20a7bf23a237589f57a74e153dbb48499b9198cff9cea804326822f58371cd58a7c15dc33ba2788a598304845142b55bafa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9e0d045857251c642bd018a6e12f83a5b7ec284bb6ccf68ec291f6bb09a0639edb0afdf965cf1ccce456395865b6e7bd6e900539998c9513d9f95d1991b724972bacdad51e03eb04d451905bb8d0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11276cc1e03fb0d25d88d804b0b692ecf2b35207c67791083505f8d2012b33f11c0de9b545153fc09908871ac508828f6c400bfb7c716f992d3231341bad33221cfc11e61d665afb35920a6a7a37d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15300c2bbc42f9410b51177253d6a9b87288438a228225c506eb10113daac3bcb3592239a2b8ab7c2d4413873d83b93fdc33ac3105675c9971bde5c2905a510dfbb3531e5d2efbc9d4ab4d8c6dd17;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h676347e0ed27770b71f726a38db540f76971d7d22ebf28ded69f940b098f22ad2b7fb4deffcccc86c2318c9d7cf11d26da1a6162a3953a378c6eb87882a1cf033f0749d94064288ba47f74d8a8c0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h47242d5f317c02ba2429057087c76e80b8ec7f4d1e34c7ad82968b4bbf5c29749f42ad37a9bd44862db86db5d322907a34b4b8b66edeeebf5f76b00cecbd8dd26bedfde0672f55ca72eb04006ef7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha6a71f9572feb6c3cb81eaf7ed3e85cd8c27e85b215d9933d48e789c956498af7a92603a76f26a4eb4cd1154dc16df62014ebb422cf0b3d6f1e9be77625559609c4556a8893e182b81e9bb59cc02;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he3f2348cf3ccc374eb414e197f4e965f8ca53d2fcac9c41fcb5a62847be11f31ded1022f7bdf946e0f6ed8278ee6330451ea4241d5538d574c944573e045d498197d582d2ef85a39db31cb26bb5f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ae037bf85913e27d46115290c0e0a9ec89aeca84b07d7a9c427f9cb568aa1ec8fda7ca6101ad715157cb6483e1f54c298b3f2b79ad29ca06862c2ef96c9b57ef4705e3157198bb4e27293189edd1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h115d28a6bd93742d89c5646f0a799acdfd3ff7da15e69e16caab6d8f3abbc749f9abacf44a8774304971a34559e83015441e93c96b165b6284ea2cd6be841c285af0802022f15d49f553f53170431;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h77d8344571d0aff350f502ffb016d859fb70279e4299c7c2190ececce112929b8237743ed818d3db2ea539d83172c7099b6ebe0c24100716e448ce172430191d7aeab40a9ee169e1b340521e480c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he234e323d19d9f89e68216373e6ed1041ce9d48ab3a7d24c89ffbc2066359be7bd2aef9d9f5710bf3f20f53e069c06e49c5960ca3bb938121cf94a8635cc8d644cd617ff5671f4a19544382c74af;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h150de94bb25863e11a8fde896ea92fe671730670c4aec08c87d4e8474bc41e5c5658a3874a8646eccb7c2a5bbc2ecb643f7b1360c0983414d7a5d86a051fab653bcd5c8238569d39713f13ffc89d6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1965702566fce43632b69087614514451760ae9a41d1977779fb7ba258f3db59192cf4386c6e0b49d2e46ea40f9fc5f255e69effe43a08eed23ae90b01c249f55dfaa58bbf090fbeb93f9f87baa0a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13d96dab28c9cd40ae84b8d31f0c3607ba702e20d59e1ef16fd937502f1ef71bcdc963bb466dfa72dd593e607a9b67fd2f81cf301b84f8607747379954fa0bbc1f6099a8f2a1aecf788d108b8b9ee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b09ee72c78ea72d8f552c603303eb38af3658c267e61eac31fd974a2d3c326347c40d67710d2c41171312aa1142ed9c015f914f2965fe5eb014486673a6d9e71a8651d3ca346fa70b707b63b079a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c77ab9b10d1c50198cd913ea4edbd72f45ce2b1de8505dc6b269ea02587c15b9ed858357b2a2d7e57e79a9162b068f747accb26eb7343ca18aefa40dbb2b6d560a1c5bcb5aa24b10fe8aa5099ed0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a1dbdfa0b53593caeeff2896284c1333f7d7491df343136141ef51b510d53574e765e0fd04c757fe3caee9eef5462cfa8a308ee3915db9d628f7a9996fab35158cd917510ef53242d93250c6773a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h194d226397bd82be3575d9db43f17a131fc9d45edd718dd9a674e42d2b1d4288e84e2602e9deeaba4607e168049bf126a14f1464066437fea56cf74999f0a2ecdbb357ca467f4085fddda4e6ac27c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e5df626ed202cb149da8bc0b29b2291156897d7d5723cdd32f175a40fde5f0c5070138e174b8aa0abfbd6713bb62679b112abce2de7c981bdf097c12ea6f4f06a3b56b58dbfc6b500ec75ccab300;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcbb1c3329c63db4c177459442ca3eb6e0933d9c3cf576084043ba0db8e05c99516a9a5ccf565f47336ded5026c951f31412e14538096a210c5bd7648d0c2ce266216576a0044db19399b7a6b3c98;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hea9ed726e2b9e4b2e3f89b638678406bd01669806c4fb23cbda5f75e9112a8aa5a76c94bdbf3ba28b3a8fdb10450708ada65a699c66db22d79c4c4e0df7989d0f97617bcbe59d45f6ccc12d4c9ca;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h29a523ddc8a8d7e451b15e519a7b79eef4421f15cf6286998d18037d9a689224a0ab340cf52f4f2823ca1f1c12072c64284f74b3dc94d315f25bf4688dcdfb46c1b9640c093a93f75d7409464f34;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1461113f5e92915b7772af5b1b537eafb4598a27782da19eda8fb07d4c4f845201a42f2b1f500fadbfdd7cc615d233d2eb9936579a540b307a51c55a4511c3158f06923f20717170dc5d7b1db37ba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h175cc1add3fbf469f22f7e18d698f39a83c6375a8c978e9435525b27649552d4ca5188e75d38e12a5138b329ab3fe1e7c6adf9f3d2dbbe9a9aaa5ba166a55b09b91816250349c6facf57d40e1e8d6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ede1a60e40515e2d6a4c2e29e4d0fd0ff2b7b0d20a3c9e607139142eab830ac69ecc627dcc3dd9df9c96cefa7a454d7eed03815164d1b12c69c7e34f71829368bc1c3097af396d0835d3d1d175a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h40dc875ceb566df0c6dff9af71b4d8c8cc8a48172c9bf6fa27f2c7c8d446484790d14fa8315b7c03c33db13f64fc0a13fedcd74c8f790ac0a57d5bd54d5c1ecaa07ed07b0301f565db054a3f0661;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h164c19db623becdbb98f872ca6adff50f9c54181ab3e1b547394538efca107a8a5441a6c2ce2e48af375660c0ddd83ccb1ad83979fe7144ebbf3426be5105dd8fd9f9ad3a7d070b2502fdd7caa6f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b6722430a05c7205e45dff077545b443d568072499a3e932d9722ec1372107e2943d1f4874b109f8079a8bb1a8ddb62b1ae03b7bd649be6c2df7cd9559415fe682999eb3af1ec458a9848c1031da;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h267c0c12220f94b1054116fe0d70cbd2f868b3d5928e55248492500d33859fb299ad87a5eb64b1485d60a10093634ae94cfde5b42b0767e8d22d7abb8ad2ed800de5f471dc9566ad373936d3a4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h54d2bd0ab5a66f08f8b6f1755428f9fa969f97c5aae21f770e9c01c294134891ef07b437b8ab19a569306d0d991450355283e53ff1c3875de22c2e6ba5e65f05832c7374a41a84d221f5b1317b1d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h982582d538fbcffef97f107dae89bbf2cc917cd99f52e85f6d6db0f7b49515bc6e5492a388907cb2ebb4a715cca9ddc4da3d2cde1523d1e4ef2f788c6923c2cd74da86892a8764d89ba540943eea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8809ac2be505bc3c8486e9b43f243cb8ff86918b6b2089e003f35e57fb732793016bf8d38ce63b2e83a344246cdb4f7e3660a7cdcce596a0e95de57891c5481a0628bedd42e907f9ed0a0552cbd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2f5a11419b627c57ec622de113b23421614697bfe56fb1a61e19fcac9944d26623730cb4781734a1bbdabf32f5a26543cc4a4e20e1a345e71b27c7ac392b83627d6e6e4d5d4135582ab010063613;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a9dba3b6d2f5ca9e6fcdc3e1649f55404aeda23519df639898c84c97dce5a93fe5a6922c0833545cb0e9cfb2df1761ee89954d504f10b7c0e75aba54cfd2571c2d91bf016700ed08c8428baf66bf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10d7bc0e17bb683ade227ec605fb89832e2786176694fab451d5cb20ba2aca76df5a4163eedd9e319ecf661d39f88b3c6906ff9d94e876fb11408bce3c82aafad26aeee745b7d928d00808187c42f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10a17cd08ee8380ffe2dee005f2be89c8d356a1af661d30aca3891f92b029a45a9ca5c0e57117a7d4b43cd9438d03b7e5cc81b86471187c27c5408d91d3e5bdb7cebe0eafafe981ff451ed3da7012;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h47f58b99d792c5d1a13471e792a282e152c83f482b0fec637c5cbd20ee8457483275ce369b1566f8d06d0345ea909251b85a42bb4359f10a7d125376d4f632048960f4c022cbd5fd442cefb29c8d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1186fd298c6ac1612cb142b22847d2e30eceead26acf8e97cda862a3bc3ad94d33903698ae06ccb05d821bc48bda06f2cf48a636112da9485227c90dfaac1f1825def930f1c4ed8786ac46e5f8bf7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b8d9582ec0c23295af2a2d347f81021c17d53f57f5d78086a1e03bc104c402bbba14336038abcf5e5969f1a2929a8f4ef456793a5920b8d3f999e4d6d5e1f84279faa524b06ed7e7e3f7405964a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd6501872e13265ed8d99a5a9262da6e40c4e93b683301774bb963e78ccc8b4adf5829925f342e3cb6a4275888c77067ab7b38d2db5dd758f7692594109a0e5c2dbbe13360de203e2b85324a95801;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h50327ed385cfcd5632c0f7aaa8c5972d7abcb4d8b3d97dfe01bf362f573b674cd5f359b56e6d19f8c859ff56527307ed5e11ac7ca33865d9dea305783aece05249ef1197ea561bf03ef7e6ac9bbf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hab9001876fe36d46eb1878d6fa7f3fa816dedb4484028d870f23c1b45a0b1d5bffd85ce662d170dd26c8b1bf503399be157d240fd5c5f5119b5cca39f9077bc4ecd06aba4e5ef2fd2fd362789160;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hedb377e5c3e505fe12284d7019e975ff2c11cccab169d41a196b57aa017474213606a74f6cb2a338cde1d3ca25bf5848f6b59dcb1aa03663cf4e355251e571f9d190b7bd1f880fb93e7f68ebab5f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4b3332c3e8e1120f67b045fa188e9ddf4e21b9a13f12753e35607681aec5476d52330e169f30cf9dab86f1c20d503293f050623b00f6fc502010b4dccd0fbb4262e38dd5c0b458b0ffa3e21583dc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6335a2e8ea9947e65de2cf3fdfa61a1950086973f849e9130be782bda09b021df2e9eaa7940cd6cab4ac68eba96f68748557d017b9f18790d2503c9a3d5b49ec54237d8d5db9be6b5ace0996919;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5aea94ae7ff5dc46d64d80ea691899bdfa314df5787ccc8887940f561a9beddaff3cda46575a98282017eb728da45bbc0a505187ec63e2cecae651fb557a51c945fbc3b914f7bb801dcfcf7bd902;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16f0816224170bf714ca0bfd6da1565a5c8efbe2978cecbf547976b25c211a68206959b91994caa41fd27fb6802e1a4f42174ff45a94bc86c29c6bb2cb761f4c7a8b4a571148c5503c5587c2a1b1d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14ac52eff1932cc87473385bf2cdaef38407c6fa804727b4c8ba9ced1daa2e18d762b15e986aef9cb8312fc1ac85af91b31f6598f54fc9cb5b3382958cd75b096d41b7e222756688219a5b88bf513;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h460d92747ee702c37bf3e10772ec7aa199f14ce458d371bc68829333bd22cc20e89880d1337116fd413e76e6cd450d3f1a740fac88ff3d5cb6490842085a07a33cdbf4c3be222ecf666657007673;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f602b7188e7c94e0cae1973c5318dd336114f5ecb13ca953b89088943837c0b9a5a389d7a865d414e3fa9ddb894b57f8cbd8db4f3cff532de6c710ae4acbc6e6d8f165aa2f8becfe09ed17a61388;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc2affa12315ccd1dd9f2422ba942a9db69a7efb9514b376e63b90784dd09f1b0fdf66dae00d6f8c118b75bdd970ce787488677538038fee60c7a83f68af9239a4ea0a6e476f46eef4487f279cc64;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b772e79b0ce8270720d2f08b1a7e1f88256871f0d6e06696a10d533b572a272200dfb47f112b738ffe95f6bbca461cf32cc7faa659f109c0ca4dab8c55dce44e98ffa2d47ccf8b75b25708f18b6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c988b609f7e5b903ad223f27211f93c75b4f43696ad93bad8957944c03401f1fbf381eb08d257f902efc5cc4e827ce772a5189a4460d3252afd5d982ba06bee1732aab4498e9d8b6b5ab1173834f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9b2775292c3836112710b8d79c9a5b63fa5ad95d3f5178f0e841b90d5c4ef02c45d61a355035ec6d72b4a069d56d3291b5d5e20fc136b238600641f01c982fec1dbcde7fbede48dbe937affffde9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc876e5d187c8aac0af380e216412fd241d2574d1b58009e6a19bb0a513550ade298e8752cf7c8150933436361cf82b81333344b317d6fccf2d064e06a76633174311b0532411f91dd217f3eb457e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c9f83f1a84ef04e9121e9fd83e7f8d63a232c1c7094a47862127f7cee3a52e0f6a79614bb5e12c5542aaf0f07474a66c6d47760fab3cdcd5c0c675505d748044e3a389d1ff6745d8e4b421dcd9fb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4bc8742890462791ee0678fb11bc42fa9dc9b2b217e6fa3e404d5b1d5623b9badbfc090e1e98c8c3ebfcc6ec98879789d7a40b20b24ea624283790364ee3455c6b8ba8e7fb70f9dc49adc7aec496;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ebafb10c207ca7fd88207f0045fd85b2c2c2f5daa198d4211b550329fcdc996bb6bd3385ffdc51ad6cb6115176a9ed745b0f8f9e1ab3b95a56132e4607235cfbe3494a6fa95dd7ed528c70cfe6ac;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eef5647b96821bb14deee1a02866aadbeb87c1958da25619bee45c923b9256fcc8a5081bc7d3614d4ec725f3f39f801d46eb6b596f7488f179e52ce0f0f87450409440b87d80fe21213877760792;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fc077060f1164c44dd4954f30f7be87f3e92de688665b8d495740f39cff9702f6e88ccf7787300b3568efd771350926e8240365e17ecfd7bb1c4962753f77b186cd0afa0e087ed8b45ef415fd936;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h199e49897050ffbd248a3547eacc06337bbf33ff0b15d92c44273d64b68ebc94e9300b3c1161631967a2deb16977fb24aa9f82e071be75578963cb6c650af28cc416e0bd2fa1289989dbbb58e087f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d0572abb6a6a048348d8eb5446b8a6542f688be0ab38c10c214c36d8a282cbf6aec0d566683ec9a69dc37de0cf3cca7ef348aee22c8956832e5e5081e9e8495c612bfdae7b78efa86be3bf7ddc97;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fa344f9c907a453e3a338b7788fe3125ad65edfd88f641ecc308a862ae676530266487d5edc481f1f5936c8a94bf0b3caf7f4bf7596d3cadfecd0a176ef61cc27a9ced0c107d075770c063fb15d0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1271b0791c05a726f846aeef88017594ed5a5f8373c326d7f96e1f215c270e7fe1be357c00a5f665d06de621d45f3840bd0ccefd991e39fce83502779aebe9118aa1cce5359418a90d2db3e0c48b6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10cdfd3064a706f81070caea4fceb32ab65668bba12101b63561a3193a547f674bcc3a9326e7150cd68cb12cf95abee175440793c2a7d9c56ea0da1213e0af320564435ca17575493ed4ef54ad85e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6a81fe4321ef69db823a6fae95c15585641ba3172629b84aff7c752fe896dc0b650b804b0ddcf3f6480df83779d6b17b1632fa0c1fa7ceedf0e635b16c7aa39e40a1736c2a102636a2f48dad2457;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfeada3838cba086afb6224d54b8b3b6a554ac0b6b643532a150c6f3fbaa9bf40492762695f6f107541e1898b1ee5f7d2c30296d1640da799e1ba932be85b80e5321cc4258e761bf4eda2aaa4fc4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1999fe128f163f5d42b4f8a678d3f1694187e9ce9e6e56f9babf6e1e1961cc9db4781325ce77457f451940b1383057275caeca2ff64b65430232709103360e7cdf407180d1da7647a98604338f040;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf13123b9d76c8597ff78a83711000522a2ae076435ddfdc6258e68186fab6cc693cb620aa770982e76d7c226ed961a787f5754985679428d55ed11c90facf46a5eb96adddcce96d2b76242c8c0b8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7083e91a1bd2892df8e719005f775c0d0778e1b575441e78ff9e1c8b4e96ecb5ca7f6b66347ba954245395a6d352ab5887d87fd9670179acd65a9d5b89a6d963e32aae7417982dbcb8afca3e1914;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he3b40f2c0191614ca532a7369a857ffdf25409882e3dcf7c3660984632633681ce84525632a84f16df762d60330bc48b134e41c5bd5ea7f152886682a39a5854059fd0cc8aafe2e7febf6d4826a6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a4f69c32481f1384a98affaaab1f2d80c603940907d9720e9a817d2c5ed19d5087b9331d668bef808688061e2542ec8d83146bce6478a55a6829ff77adf08b49a53e992c3098617731a68832d1a6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5a906f011b70c92cacd9ba8784349cb734c1b298a36f3fbd07c2582e454bf80eff9bec83eec676dd48c2eb3d5e7ff1125e933a3debe171c4711d30d70b46d44d51075b4293ced734587f3bd8b731;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1afa70ee25e3322252dd112e5faa1af030f64c8e8d436591374e1df7c5f56b6c59acfdfbf5fb9f43b9dbcde8f853ebe4630386d7544a897ffee4c1c3ef84750eddea9ae50ed6839c74b56f1b4118b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h67dbb496b3628a31764b429dfb8a65ada4ba293559789e820b253fb2dd730cb769b3f1b9d85310a56d8316b46a76f8a34780e28b7882cc408bbb833c3f096c3c4b5a892c8f2fbbb773ac19ccd7d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c62e583f5518957baa48d84ae562b7518efacd7433b350fe415edac275d73052331944f73f98cc9a0d0678c09f1b20635206742bcf86e164110d6563485ebb5059e64995b8aeb1fe5651b764a6f5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3b131a380c5cebd2ae7bc81ed276ed8f2eda37b4ff75c5dbd782795bf4a901efa950287841f45aba039dc6d8e7fce7d68bd3ebe604f3e7a2a4aaa617f4f8f919591e2759d40606ff671fe67e9c30;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1797c0c8fd44a15a5ed13e88bf2370b15876246d22a2c640de03f6d586901d4c8d5abbefa04e9ea6f29ca09c5753a483c39edd2dae49002b23c5d436a01f80bcda9be6fa2f4cb5876d4cf775f6e12;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heaa944763ff57fde3b6cbda19aa35343d9b29a4bbbe6d02674ed50c9b9ff246b21956f65eb93079ad39b3e4f1e8e2071af035af98ec0085f8ff1230a4b9affb95a6c346b873259eab157904b204d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h577f4cde5be2fc1a734ca40d7dda37dbfc91048dfa861dfece52976ead9ea54125cb0d01ca853c636603d21fc1cea2a2d8db1dfaab31f2b72d04c47684c1e4f463ac29bf4cd93e812a85fc59ede6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17fb6983c60f779b2043ea0e719332125af4109fb1bec1872fb36b5e432d386ad4b0edb8bc19ffb44d9b0d0828218c986510c0216aa9c5adc2bb5ecec1de8ab6712aadab4ab64b127a2acf71ff608;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4e1cedfd37af36d33da355f3fac907a5f21d066e4ff4f9bb816912bf878915cc39176759bdaae29ba74a3937b897904e352f2be0beb8f77bcb963d3c56bdf03dac10364fac09770ae38ed7e201d8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1725df2ae53868a1f099a316e7dd45d30d7fd3b5cfa96820ce50e84d2d0018139375730ddc98da7d7b9ebaa41921e9c44df29d63c7964ae2fdc5390696da6ff11f73d9e7b9fa76801643c0c4b2c94;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'had05eeb4ee184d412d51769edf65657a7bd5615b12fd9a2a9d8db07a69df37f645ea42bf198959f51d7382fd74b5ca4713e898779d7a922178a033bd90a332d29aeb7f0ded6d44c1851b48f17d66;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19e815778bf658c4050efbad89563aae9256c1bb10926f9420dc8df69d318662b274d428a78f007ad7a9d59bb90e1ef07bd6843340f918c1df81c31f34b84391db719b38fc42a676a2cd4fbe4cd06;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4d497776b652a94dc13d48e1b19968fc29b2a907abbf4d34acc3fc709aabb95de527d4f96a6e0b312308867c6cc29d3cdba51d685a73ba23422575bf73dd0ea3a108e23a71809120d5d0c849e19e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15e59bb8fcf17fdc088bcd0425b3512e552e566452e418d069b7c7305478ccdfd2f8d29486172ba1c09159039696c22e26b6023cccf1107873915144f54274695906016e112e4d808be611418f232;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5bede2636ae7f6833e9384a306d68db3a1b2c7de73bd6a77da3fad2df49388f6a7c14eb4c4263aca5d920e2b54df16d0cb792a839fc5077979efdee4d766297aac168cecfb3ad07acd5bf05244e6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3dec1c87e47f6bf4848aa992626c18ff3fa6c7d744bc05400ad9896d56bea43a98ff0618d2283c758de96abf010c19c3a1ba1268471f2d329a2cf9d420b2cac1e5791578766cf3ed1c918ead5a00;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h72f52dd9ba86ec38e07116313fe66b0d6f540890964975958aaa484247f535bf291db9e1cb6a3479a53176dbe8d8b067c8bdbf5fcaee5eb5e9225a6dec6c54498bd91bf8c5f4c88c0ade3bac911d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h29d4382003765d30f4990e1c5fd0326f1849962ed89d8b452e8f3c15614f81e5a16ae5c68fbd2760cd23c43e9ef5fd5056907d41ccf965685c66609f931bde01111210e403b83ae9718a570d7d12;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hba671680ff0cda648fc2ce56e9ac89ce5409532d8555304dfc4ffde0a6fda2859ed7c014389baf7204e15b10dcf5018fff7dbfaaede84e6a5e613e1a78d55c876188363197d72c9e42c4931634df;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf8c78f9ef9894409f2270a74eb75ba4b8b4f6178129ab505629f749196c084ccdeeb1208009dfcd037edbaa46da278b47ae7dec28b33a543cd7e379a7dd8ad88469d6f1d3f7192d4cb985db23ab0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2d54aad29667a3e5abee7e7a6e2004cd0e04a0649cb21dea0fe238ef1e5735611c44637018ab9ff27c18611b2fb98432b4e102081759dfc8209c39278ffc406a5656477d397da6452c25c87105e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he85a549e94692e9ef649d5766615dc2753ddc72002da45d307ae6a62712379478efa2306d642087549302109c7c351068a7d3995a0c8165876c26b411d6b3f0cd65d7afd4d601cc8bf4567eb1a9c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h421b5de1720f558b256692d769856f0cfcf79253e3514dea96422602c86365d676bd0577732326d03fa8c92d23865cc189367af972e7047ceb7da7fedc1b3419e2142ff3303cc7bbf7235ea7a0cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12adc8fd88e66b41f38a33fa92fe84304e3152379868317242517ec47ee817c627462981f7591ff6e5d3e7c12d9905173ab1635e0e9c521018c5d3f7b2d2a5bb05561f425d5df534164304ff5f25f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fe06b25821462bb91adc794f1eb2fa6b9ae72423a14a84a3ef520d04798607ee18263796b1a43ef92cbb88eb79e4622d6364d74c8c2cfdc5da84fa4f4ad1487768f975e6654f9506334303ffe46b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdb8821ad822b3bb65d324c7255be6487df45cb21f2b4c1c221b07c6a5749f8efe6ba62fedaa624033371b2b514f937417b5a3ec5f54bfc65513ad5a86d2047923f55335cb0b8778f35c014c6eb60;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1383c718d5cf70e68d785b2130047d65110ef23615503d1b2e87e87fb15bc0c3112d545fb10e592a74d0177c4fefb57abefffdb423410a395a312749e1f5d144ee0822d7dc0ddd1a5d9948c1b037d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h66fc2ac935619c6cc7845a02518fb20742b4c4761fe84b49ca477402624390928a7ffc5a44461c9d864fa7e6097595f6d8e03f68fd54b45c9d34de7d443f204eaa2d7dc306d8815414a42f452771;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h369e685e378a1b24c08725ce5227573e3a37c346c2a05d341b87fe1e6bb14e8b1400752385015534f071020b77e5be74867ec784339d521b4f1efd760acecec26c3465f0387f672020b6fb275cd3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h150d56a2285e69be4276bcbf60c077315bc511eac2ced2bb7e4ad7100477fb38ebdcd4afa4ac8a8bae008f36aa3adc15389f53d4fc50c29677538bf92e8e4968105932bbda022abf815fc4b4e3f37;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc0c73c167dbf65884acb37c55faa8e62a4a0723a00d1eef2ffd327204e3df196635f6aaa25a2594075170472b66496d2f1f3f2f0ed494610105819563a1cb2e2c1947de10ea503ea126c0d8b6ec6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e13995fb8190ff937b992dca80592029705a09aeee7f077713e63968651950cc4ae6e441d963c702d2b433642c468da36e9dd73c9dd597001133a1fd32c91eb733f3bf2812643b827159722fc57e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c5655b74effab5560ba046f8e31e0b2da173dfaf7e9f3fc7de0e3907d4bb56af464290e17cafb033f6d847aa7cd893767a6a6287583c3c9f2c83c11bec913382619dbcd99e5cae744501f7a4ac15;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd620a6d8e16a265fd730a6a3083f1ff6b6002ffe8856e09f490fea62b81bed6565d1603bfaf9506680b983aa2e8277314c0dac69c8c92196bcbd059e010f53920a5c17198c561bd7ff01c4a84a8a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1688d5d64f24419dba82aecf14b75633b8b6f58308003eab189884f6dd2e08aec389b34272280d622f89d857f25836616d56266eba71d3b335d3a9c76d5ad61a49f1f2e28dbd54ab6b22e87ccddcc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he3099be1618be84d7a5184ed751184079028669642e26ed60dae60fa03f217feb7ea72dc0253bcdf8bd527b2ee052d08305280bbef85743beee08b597dca0a43142e7a9cc74f5def686b096c113f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ae1e37a100356fb2c5cf68a5ab01c5213ac29d252dabc436127e76560c654ad3baf1f04706919d42680c60252441cb9b6add546a19048c470ca9f01f2d07ce023b28796e94946608d1af57ba0e58;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11d8452f9382bf5d727c0bc821b7932172f02c2f76dcf492218b357962391f1a93ba0ca8df9a71b2c06e84bac4141fb77d75a5dbd7ed4740bac7d209021988375fd3f8c4f58155491a885ca40bb64;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h676b54adf4b70a7ecd26f5e95071409807aa2d4c1833cda3321bd0830f053f1a91d816c9e09276b52072970beb284abb01b97ec11ccc8958647d4e577a911cba46fa5c1b3ea4c91e8316731936f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1381b9a9d66a6f6a3265583f2e158265b8dc6b86e051fbfcbc044e07c0b90259e758d0b7af277d87e4fb1a273c5fc8e9310200990784ea2e8f8fb90dab6717353e30e214a5c5435455dca2bcb001c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h169f6433610e2a82017e8678a4747e2794dfa0e2d11070310d1eb1d617190477c1f0d1ea73d6a3140fa1c175c92279a2231b5792379095a69e32d313602446481fee87a39165eddf9efc55faa78e3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19d3c1c5bfaeef6200bb2d17d4c9c42c886b8139a0161286e26ece1942862c752440bc7b577cafefc500d5e76e0a44259708e2f7f5bc603ebbf991ca765db9eff00b61d380ef514085bf6d0ba0863;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a8dd9ceb8b2bbd5731d1a98474481e98b86bd8772d3e2096b8e937b90fc1fa8c1573651772de16b0a76eb4c2b26be5023839fe5b6d20ba515f088fb2eb6060f5b2801a9761c450fc81ff6f8ad4a7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h127ee97019d05f3b961a6e1cb1f4f14f8ec5edc9953f8b76c8937e5a1ad8d9f9250ccb103d0a04cc220c055aadf56ecb0aa30b796865a2be8489c8f4a27980a28e10d86be975f9f31fc0c04dc060b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18694eeae06ccaa5ff8d8234d2dfc5b31550671316d87e36064d00593ea9aa36a981fff5bcbb240e428c161fbf8e747fa8966835fe6a47a6902e9c532dea01388b614e57828259e380970e7d11958;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7381824f3dd9ec6a51cee15d3793c93b148a47be8043b678d40c567d72963a33c32ec1b335feeac69604cd614037857733f2a8fa3d1604d05128edf4dbe5c41e2c65424a7ffc3b31bed9801e333e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h415e8383b48ac49de216dd2222ed75299c5735ddda022f5b608747f0374cc2685b3e6a3f7c0eb5dba0c7a3f364efec95e220b94edd892af3d27cc12979b81cb0ca4e9c6d71e3a8d4efa809fff5fb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f6dc45d8b3c7e58fa056490dfe41e0e9ecc391deae8baf92ced668fd253e87b0609dabed8875844b77630d407d70f3162fc378068e52e0d2f34c1c47e74dd92efdb3399297f1b27b9331c6c39de;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h82aa4bdf96baa4511f9f707898d6f298555215dece388f01739bb14911257283eb7fa1575d4682a48371d5e36191e1286980350e4606e8d0bfe3598a96448598f9a0ced62affa8938d58040c6884;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18bc7a4d85956977d279e253893e61577e9c869d98e1fdb283bc59ebe73523af513f510e424078ad3fd1e18f38836c83dd33bb01baa571c5d619d52a8159f466f7ea7b0249daf25f9d036609dfe1f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15f4fdb1b65d8fca603a0d5eb774d629b08908d8db77c7a224209e9da92c4b81dad689c684be9d0e96c8f9e1b5522fd40a921ddd149dd7234c58e8bad1a9025b0419ef2b05e693b1ac8506af3a1fa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc44f4f5fd91c8e56f95ac0342759441fcdfcd2bb72ea6161f29c7a610b296118102beac6bb46192b0835a017630bf2d635145a42b17e5b3d729dfc308fe2ee643d55036737803bd7c214084aa632;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6080f1031051a6f85f7597ed3f851e35c2d98287a919ad4283ca23afa0ae5dac4dcb3872b66def6b81bbeefc058f7f581e250bb613786eebb2800aaa0ff840402d5feb00ed9bc3cfc0d2f61bc02a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19e3b36a2315d1d091de46fa654adf3b9d6ded631d14e115520ca4804cc7a267436d6ae46efdb4ada34acc87adea13945607887fd007870327a2f5335159a9e91f83cac18d01d816134be337e1a8c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h415e53473f62bd5c726604a50a9dc1633536596a11ce5335ca74fd5be6b374122bc9927cf83402aaa7a54e0fa8997d9cde1b497de7a8eff50fd89efbf1a8e12feb47e8f85ccdbc599d4ac49b4b73;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc3d17288f99eedc47f87c89705b13653afd6a36dcbcf849084d9467adb481bfb0fb341ccbab801356f0ccf6923db6477a290083cf5ba0f150cfce6c06adb9d5483f30f84a6ce8f478d1f445151e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7136200f2b1c6e16e9232ca743a9d84e7fd8f7d2974dfc0d2298f88e17ea891d0817c632ed883bc7ebce310153f2d3601f384dfde403f72a4bb6cded3b982700dd8125bf76717a3980fa6c012b80;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h192edf59a13d68bf2598b04493abd084e75a8f30de72f7df435aeba30919c141cdc2489208a3dbe164b9d7d76acc70760bab42e72dce1d96291a94f40997ef45624444c35588b42a6867f184adf2f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5011b2b67fcfebc2f0d79d39db4bf0f741139590a660409aa622908afba381e54336a167c9c78bc28fb137f7f6939de729e21813edf49f47b742a8e279c12452cb291d40a12ac0b127de65d12d77;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h142904a75207cc99c06e97500944b2c013865563f4898caf6f1317226dd998d05d4127adb70bf66b3a0a662accd4700897481808867727d4257d8806210411377f2cf5b2c80dd3425f1a0aa0425f3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h98826ad6f51471c0f97c0d43e8e50d0a504a2307b311ed635b016772da5e8534f959414401f9dbe80131feeb65b8634686bd2ec9f1f698aca56fe5802845ba5cfe0b62c6bc1008e662decefb35e0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h886ac7a13c5020ffad3db60b5b49e8cb09ec2dbefc47a4abf547d2c0c2295e560c0505d9a39bbeda13ea0a99e28e551b6d1a3b41a8e2a4925b647124aa7875e1b02ed266c3b05f802ad1199576bb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf46b8f938f74e41869d33592ba951eb7cb74eaab5bd7e76199439498851fa141c135a3b1cad65a7d1396c6150308c7f1e65cac4233840efe5a8945b74cd66b25f0e35ecf212aa08f54bfa7a9c99;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h24730a7f924612b36df79a4d0b2fee1abe2e5ffc02bc57151cf194bb727ac696dc76133590b06c310468e6146d31706e8cb504612ab8e3b336a3ceeb9d63ce68803b058c175f9ad35e9421f9449e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1def0874973b007ef6eb61599ea39050cd03b4e36d1287920feb5f704849eef498a5a79acc0553bf49dcad2df4bd53a95805dc3e14919ea1a3429f386976c58b366b98c1a06917b7b68a390342369;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h304104ce87b53770bd60a6a309ddd11935f8e6af6271de012b73729479ec20c20bcfc9c5ab72ebe480d752deb21f14d8edf1d2b9d3109becc1c5af22ab2f96771356ab9e5066ef09b27f2818ffe4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17b07d0b122ab9fbdec1192daec0db709d6db22477113edfe89dce72e0b5e9d42fc634fed8c6e9409cb049eef22b68ba365fc799e83c757bfda6c921f52098fd9446068c87e95ad76ad6de10b535a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h138c1b9f97549d60784941fc6c4674126e98e9c367c7098a9bd65d91cc35ced784b987c3cd963c8bcb67ff845c7a9f308819459d505fc958a1cf4cfccb3d714e395673899b03e40f4c9ee3be00100;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h54593c5efbd2640e9338dfe81f0482d180afb057bc1a05961c2a2558e92a3d10028b6a1f9c18de9e11d3ab6c507a2d28d0da3ffec72210901527c65cc8ab35f165648b528b72c2b6e2a7f6a58d4c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1afc04a3387b06eeeb94403476d05bf0d8189e083000affd49b4dda7ff335fb237c0b49eddda9859a9385a79b6e32e87e1f787ce99f4f7e93cfc58bb81db5072863992ea33ee357736a4eeaf55f9a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h195b3dee3f63ac2fab36b906179ba1d700015aa91002665259505e58df5e83409d844e75fc06b938c3695069db71fdda15baa5c971472949b2aa24688375cb53a35d8ed971d813db51b32c6edc95e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h188589196be67337115b16375aad351c125f579af98dd767fd39d3a7d233b474a9a452ec8f2bf128b044666b08274e93c6592493a77bc56e87f93652d6977ab8f8f35a08a3b32ad95e8558ee28e5f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf295bca39a5b299cf05f8f9f8f14378f55295a582d0ef5806a6b906b6a91fa5a19b2e185e87a33973892655e0eaab5fdfa95e196fc24ba5803c55bfc1e6c802b02c7b4cca6cf595b9c93d0cde76b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h120d8fab3340755eaf016e9c5511e5b0436e55f6c2914adc4be07161fead3f24e037e91236eff29ae584a516b4ec96bc514bd828e49c8bb8445535cb489496838b761ae17c32f7db357d53af4d728;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d3f17ee7e5ee00beb794fe5f879885c51a8282956dcbf774183f8ac06388b8ead42dc8e44432ae111b0ebaa107246dc08bca4d1da42cf854797d72dff015a1c2cbf6fc8a38567212ad8d45cb89a7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1823c0bc4bcdd73182e80c37930fc681fa557a44d2cee444236efb5c40e1444eda7b861bb0f2918da628efd012d7d1f4f86581fb4d9923010830def6d9b5313bad73cad70e04e71e863c5d3c4cacb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3a7bedc2f03bcdead0f5ff61dcd9abb5975544f77a569cecfe05f7ba1b938780d16742a64e034b9793c9dd829485ddfc4636bfdbad48aa3157c4502754700b7087219c53114b261a0be0b0bb7743;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10da35dcc5a7b2a781ace0ab1d19cdde702d6de874fb573bfd86442ec4ffd9e9231753a3a6b3f25694c604da2e00ae23e17a796a24f75f2048a9f4dcc6e6a56b5d6c267392f6609b6d32960800863;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13de0f8bb046d58043b401b62a8611de255e070d3724a43ad447d5ca247c246a024517fc3f709f866e46ce08bc4692e1ccccba53287ce4efa1e814a82ef5ea82abfd7619140a7e050e020f397fc0b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1055270f39febcdf52c8bd7480913f19b692873db2bc4aa0605ba2fa301368b950c0f28bbb1069667aca39e096abe0cb22d962dff5ea602c92349c5492da39a9bd974a2694ac298702137ab6808c8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h190c686ac7e9a1dd3d2fd45b202a23475c750f5204c7065d203ceeaae58a266f5188b923305378157baec9326fe804e8da212b8879485e98e91349ef912d00ea54a5af34a7e73f0c75aeb5445258b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2ae90a2487fa50c13d198e9af02acc37df1fa5377a24bb6607e043b50244c22c9a70c7e7bb222ae874a84e24b08115b02f25475fa5a13824f240444512bacd16c0731863fd66ad562856236586fd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he2e46917a6483988ff2a52b4700d66f44a210629c62f7ff110f589246ad9652898f2a4d15676a2fc592f1cac990b7b511b581a67cd645d6738fa8b89a337b2772a12ee4e407f5af222932f4f069e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3e507f571738733a129aafb016a7f1ff549e7f216762d9fccef703432bb0a9942f892f0c505c2806209353286fe73cebc80cbbcfa3e82870c242d51bfafcf7564b1524c408c2792b6a0d152a7461;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he882a5a233a4fc5063ceb5b7b25cbe9de6e207a9eacecfbb80e9da2c8ae9b7d13c23bd90a8fb40a16194d9e04787d1af282109e74b5f87bcea752e9327c818ad6399560ac8c4e0d358829e9bca15;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19cd5808633fb9427456ef6a9d94f0ad952aa7bec1eeb9ea8db2e7d8bf5845f0e210e8b4b0052130bbb1929b1698f77cf46042c1b6e787aeda240a53d38b94d7bf4cca46b77f6db4153e68a409f42;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h101c0318cd57c4bd52defefce478e452f818f33cd9d9973e0ec193ca7e7dba18809dc26a47c7ee762e38450a0f1e969cb6fe06d5b9ddadd41175af5cb825d70dfeacbc6b8ddbdf79ccb412ef788f1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h161a119768b2ef14478815f3981df133eb074bd3b2ac99bbf259d36044e1904cfb90a5349bdba56a0f574431becf481c49822d037008ebcede7c07737997caa28f635584358d4fe8eec8bcc09dbd8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1517a680f10da20b097203993aee43937bf4b96af4af8dba36a16728ea8aebf28404f9a3b4f399d927891061d948313054e031d67f0878f5daf36419fd180fb3b9721a343ae812decb13582ab8bd5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h910977d0a5ded76098d435f5fe5666ecf2734b41e3a9d632b404f81d003bd45579baa9e058b67850c089c220fb75ce9479d4782d78603f934d120e1b4b34bae5e475b44124ea1bebfc90725da6d1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha9d4cf172f3bc1d1654cfb1ed627d60f394d226789194c36e3c451b808292e586da51bb7e60b54415896cc8f1e3d8dccd123f332a2233b01bc3ee24a4dffb7db9929f43f7daab77b398e4fc2dc7d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1baad53942a7d3dbdc6d5abf375d0703681200d571be8dcd752fe421bc973f054b525a31c6a78c4e6a8787d87a3fedffbde39b2f593dcc6880ca2295de27dfcf7a2dce0cdd4eb3e0ad7db69a661c4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10b56584e0c8a216dd46d67b1cef38ba722f4a5719a3f763090cdf5f4f47184ed533af82b4ccaedaa906df97926a73e37c963f386393b3b03dfade66519b3d2470665bc989f07a2a7521a4f870984;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f5bcecf9dde691dd87e82bf37156eee0af78d0658282b6ac3602ef2ced6c3035f9ab79d8978588fe3e0406b4f54171a704f7ddfefeee4442e9060f5e4ed289522db464b1287f9567db37bb83c43d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h140b989582b79b83d09da6e6f308dc2567d1abe769225490a7c4d6ce60f170a84281d84a0ba9089f4b60f1fe25b8148d577355150ecf9eebb4dc86afc3eb1f419bba41938ec46fa3317a3ecb83038;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13de6ecd071c5e4a327a587571dcd0f0db61d19795307cf842b1270ec6599dc325e8fdcef772a8730dd51ea849e444122258b7d490c50bb8d4ad83c820e4c116ee5fc1f4fa2d8e2a80e622a41a157;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13105c36b87d432b41de310f77b88164ba91d21dcb6eb892d4de5536b69608aff1e207b51693bc0b5307470e580286e2c8ea6c0c775fd37e54846262a0a31e3075f41ba35eac9f9fc7ab2671fde8e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h179203226a279f3907ae65a5c22438c751e96d33c41fc9ac0487c98a220a1a26fd135f63585086818e42cb132ba71977b422f9af2f470f4d8a15b1b91ecda0a7b4ce98ddfbb8566067e3edbd36406;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h953f277bf34f84f62f1d6ce49a1cd0ce267acbcc794523587540157aad739863c6c5a2cac457df630d91a47b49d61eb2e56dcdee0fda2d8fa4440d1df92a395073d7f1db8a4b9faed4667032505a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1812c537993cf2b92917a066116a9dc94b2278a96eb78c220649cf063719a5f4f3a92e988bae9a3c166e967dc52a28fd581ce4fe878c566b9191233518a65ff999f23ed3a30c8829745eb9e2b3a76;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b408efdb21dd2a7818307b76a8009d68fc718d918878ad289ee9c87ed5fa6b8bf84d0268ab1c86b9a93ea15586d280449ab1ad0129a328a44e07bfc72aad809df0c29bdc1cfd72cb87b323f93dfb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb80ea66ab559956c9ba67680bf4ec2e2751a25a250bc8812e5aa3d0e9abcecebe8535d5218700f3540b52059046e9ca74f83f82d501c48c9926daaf653c261adb6613fe8feb95f4b60f6e44a8a48;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16160fd671610f0257b3bebe284cc3b48ff255c93f3ea149a2ffeff4899aabe925ca7550b314bacbc397c833426a4e10b5600c7e96c7d7914a1930bc20896f46e69687043ff802715ff4294226ef2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1517727fedc7aab2cd7323f6f44882fa7552d8655ee7268dda7d04bd6f6b6d7d1fd6a0472912238e3748ceb7118afe15a09bae4abb9cafd51da9378a488fd01ba3a34d326dfda63f40e456e68288e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcbbca7a94ab56c17b5bbde0fbd375454dba99fab0d2a6b22ab80cd065c98e323e534ac83bf69e43b7e313fa5dd08a24c5f82ad59ff70bba29002e03ae0d88a668cae2f30bbe30516a5c3c4d65acb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13d8da446f895f42cc2f32197fd32f3cefb2f1e84943da104e8a3ab79ad902c9a7b0f748d47c0c2ed76abf81c77b21345deae178a53c0d86c4662ec0fec3ae5c3863e239b321e840a1c90301f7d16;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12d3595715ee074637c2b596b46da8549325329799db4f81ec1f49337e9c11f18e2800e1f7829a657f4c6ed41b6d076c36488677162498d358e4a453b5553bf1fa59085a97b1460daf4bf5b57ceb5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf9c1f438969f9b59aafbe00b345de22ec81cf5700cca84187ed1da912dfe148c1dae020d3e02d4ab6af096d50b2e6dc15cfbd06cd9075972415d65cba280c9a5882624a566a13e50d7eb3bd89;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7c51f77762dd47f59e0b0c11339a15c3f655fe97637833dc117e6df13ae919c77363d33d530f016f3bbe8d2ea0e4ba249c42951fa273fe7ffb19ca9d044cb0e60f11e0ef5fb6be4388f1d4eb025f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcfd2ea08821b62b229e36ec157e430b80bdbae2c8327a289f46ba07ff99b0c3605e5eaff0f5baa8e62947d434d57398d70ab06b0335e9cf2c6fdc80ef07da9b2c105a772da9c587535b351826741;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a3247691ba7989b2e88bd4c389512a41633355e9d12e263ea31ad60d2fcc83a3d141113a59b8ec9fbff5534311271ddf203dc5d94b718f65cf7c646402575aae689f21646b886ddcdd9c38145079;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8225384a193c3abfb3d97ca34fffa439b6650b38e0ef23cc7f0dbd65dcd0d7e725f5d22eac0cd3207b26a58eb64221bfbfb0262c06d54f98d0f4fbdd6d1ef7832216b112a64c2bb40d4a2629fa1b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h92e6da7b95765db2b73881e42824c7253dfde61da1a6daf37ce2a25d0c552d1616290af71d567adfa3cbee255c61aa776b33fbc772cb7d20827659b7afa946c405d1d4f3ad779643099f30f55d76;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1638a399c45b6f2a2b72833d90f01d1d7f6f5fd14ab5d48649995cb2be2bb0f3ff94146e1f64aff1dc7911fef0a142e3259811f3d4250fbe1e6caeb8c6e3e538289a18dc612ce6a0aa58e4122f389;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc28b3a83d8dd3912fc97c427b72832208851e40758b2d6e95f7381e0b2d165fea3f187768956ea8cd4a5e1f496df7d58af38cfe8daa4f3ad74d6dfcaebca1d714a16cc62ef283be274e9f5ba75c1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e6a5d76e29373f149c86380ada1f7c768a723bdda7e2a888a561ced2045eefc74e037c18ee5f84cb27b91d9c6e1711950153a7888425cf0b6208fce98c7b39231661da073e1bbc10b438696302b8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heb3141a6d079c456ec557bfc43008eb74377ddab7822f2d4d2e1d9da152ca734aca7052cbea4bdfa3cc769b7365dfdd8ce002c760dd1ee041136635e89f970196bbed86c91aef3b3b3b36e3e7bb6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19f54da681726ea49f085824b4f4eacb135426ec589ee5b36d725c3b311b55f8d66c0f4c09b7be937ac4deb7f914a13e7fd50d1a11986352eb7c9a9e3878406ee92d0600b9bf09ccf8413ee96ca53;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1163004686ab400110a4d70a5e089b5d1c3e871d9007a569ac23b6655b5ec93b390569c4749b959d023df58da7a5d9378b846e923f108155e66a3486cab983a93fb011b46a4d0981a584977fb7ea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13dd21158490b40d8981722de1d2ae876cfa45ad18c65bcaffdbc67623cc700ae8a1902991b3a1de939fe1744ff7f995d68d9482e15d329fecd4b0edcd63873811302883018d828b828b826b1ccfb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f71fb40c1391dd453973cb303fb63d7de47b6a17d250dbb3f24b8744ad066e35f3daf3c659eb9c209444a26ca5bf19ba9782b19ce056a4a8e37d3c81ce233b789aeedbc127761a59434e97a87f9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h110df273c310f8cfa5c2f9d14c63ddeffab245bd5edc8619360d8165316b3adc1ac6e80bc5c224107a60bdf9e3cffbba388fb5159ac2d866f840e87478a9b069f6f1b3289a4ce86297dcd8ee8ab12;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdb3ed97baa6cc7f473d1228df8589f2b3c75ac600d0d0b647b498a513c7ed1c4f4b96cdcf3829080d430d2f118c364ec53dc2be9e96b4d3d8dc1b9b3bda113bebc1af2b44b9eeb03e482dba60053;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e4e1ccb989ba736a70e8c8cd904428736e29d9da13fcce63a420ff4e88d6681b3864f50fae6cfc845fb3b80c5d4c2403e88084234989cc41ceac14f123e19b5cd43dfd20315a0f441445d0b85a97;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b29b6df8788397b809c73cba2977094a821092998935ceaae00dda9fe3f6f267767742ab0992eb9f10f50fe6c8a4a0eb6a528bda31986abc5fcfd3992b9fefd3f016dbc07533ee4d99ab826bbb9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h83de55a72502a397d8f1e084c81401ab67bffc46c54d12122435019cfb85f73ab154e085d8b2764f329911917d2ab3a180bdcc259eec8e7e6b18c8f8cbf9ff6ff4a1736fa2b1deb39a3b0d7c53b2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16a1d31699a24733b217b8c3bb839b0c0a9b0010ea8b272b00ad362238a884affbb8f97519c6754d8c829d5a060be7da017e311f33b91175cfcb04901fd33231012539d1d1238f229f96fd5a165d2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h52a95328d0d9baa74ed82904eae35ee4f2e819ac574474bf28d47572999e1e8bf1911a24ac76eb9758b21113c91d2a2384838240e087f60cc6c07849da7dfbee97c88d2763573d021eb39f62d2b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h106012f98bf76386d87b7e4182f90adb9df852443b1d3dd5c7335aec41a7e991531b068af637089c73f1bd62016c6327787823d5a04198d5603fd0a2e7d89d9e928b3b6d691e12212cdbbff236638;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10ab739e9473859f0480adecb2c641c05afd5cb5528da0c07f14b5b8deadeb02a6746aaeb2692531ccb59b8a4c9633390afbdb111897bc94901f383948b1f3ac361e9f3ed114e72afab1f966be2aa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d0d714fd6f2148c4df973b1a257717c0deaa2eebf4ad88f4f93ef9d090e1c72372e67f06af725d28d13338c27097d1ac96741e90e18c111acee363d6f5c40cbd184c51493c5906c7bb364e492ab0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fb022535193a6609a562c0708a63a8155ad73ddc86332b0fb41d28d601466857208546ed369095e57cb30bb54b55dcd3b325ec3221514b46ec47b51562e084017d8fc2612fb89426fe86b12b4ee7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h138e16f64198e5da3246e8731f11553c55fce18e5ffbc653bc3f3d1ea20e3e11958e37e389af019b9b87c3317ff05ffa6ce3acf8272f2593e6a68ff757dd352316be1b29936c16523cd3743e7a332;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5d6b29f26e1e7e4f3237bf23d5f266579c5b456a1ee5330e54e9def843e768bc00528074049753a682d1c37b9618945a7f274732b601beb7b3574adb7a98f3b2685824fef2c27674d8e80c1e204b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9b6adf4293449ac81bc54125bb4598cfda7a5df10dc44319be98f6a3f083ab5a20204459e8c3a5015b5b9b10965dc2e554c4b8668f59d5ab62fc2b37963fecd376e27397b94f8df45eed96a5779d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cfda99a58521928905bda610fe0eff568c3945a3b6e6d648337c3edfa7dd769e1714834f87b56155171bdda54c623d38de900766dd3fe70c3fbcf7adde55ebd25d203627bde9273812427a5a7bb3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b84dd8ebad3ca6b2cbe8a10f4391c6916fa83f668a413de23be07bc13bad1eb3e5f2414d05764481b19357d8b0e7dac66d36f8387e164908ebc58333d6e50a169e1802ca4a1ea8135898371910bb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13dd23c4e30eda6c1a5105605ba26b654bc6d5955a89137668bb46a688091c3fb20e568b41ab6aa72d6a590cab88e2df61a5eb92904b70893e87805536cbcf48c931d0b2881641f9403f9e090bfbb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h66338d7899b4c9a4bc495dea283ac8cf6c9c8a4c8fe1b354d7dcb371e750c896844a6a8e783370df0d4c0244f2ed249d43805e6d622e7aab2d26ec53c40ce87cee8e7b34ecf912a9991decdbde4d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h106c033ee995747449a4121acddacdd0ebd183628e0465e8fc3fd5e1281927de71ea5acc5236e06abc5496b4c21d46167190accbcae332ab3b80edcd0745aa3de3c985677a340c089f5d909bb8ce8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19a06336093865a9b476bc2a1310fb46ed02e974bfb18315ba7f95ef49185c3abc9117ddd5ed6126d3cfb2aa1bc884c9860a5bb1fec3eca47c88f3bfa9853b98b11512ec619ac3d5cc261cc3352cf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h74d4cae61acaebd100e36dc7f789aa1c988c22e141fea380641f5190cc1d4b8f7b7f7bf7a8e5de7d4149b062e7aeebb4d4b109068f61e18337b42e8b80607d6e41e288ee2a2f3f6b8447a6108e38;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15a894e5e62061d47dd111eeb2f719c20bde3011c7d8105f318282f3adeef103e76ee1c8e559656632efbb81d20d0aa10bbf193fa60403c64d7784f7e4d30108ad48fdf6d0eb7b5097001f23932ca;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb76e75ac797e0e941cca6dca91807460b01bf89210a1f0113a8ea2618f502d35d8fd29be60ae0540f9c70cb1b087e9994f95c42effcc9cf9bbbef83206add06b848e82c7e4879fe1a1677b77167f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h112822589b705423465ac6f68b03d0d26f4a5bf87b69f8dd96de2e1877d9f2bf72ad6ee3e0153aeb84a11da6febeb801230d991083e86a500a3eff481caab5d14ad3bbeee51583ead5bb6c89d51e2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14fc9074c0654108a686e209e60d94027796026c6095c8c3ae1eaa0d8706ee875a6e64028823c558095be5db0030492bcf590f606e487555eeaa86d9d13b8f52a89e793ff65b4ad64512a89f82a1e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6a50c515d3bd1a4eba752e8f8c54459ecd917fc999ee924742919372c419aef9468d8fc846af731d6065284822d6ef5417b60a5c1582331af03c3182df462b1789264bac12b22fb33bf09aff09e1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1132d8c450a8e16ff4c2b63b3c06309b75dce9f9e6e0f286f1dcb60dd3824af4ebb5af643f175b81869c690447467b424e47e223acb736ae88f8d5dd58c7a7243840f25a3291ecbe8b7109f96bd4d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3aa665eba55cf747c9abd3afef8e352f9200798cc6c3c7e8ea8476ab2af54d83b2c4c56aa183357914795baf1f3b7fda6371d7c6020be092d81ca10e3035133d4454d5b75f2d8f45bfd0b7eaf0d5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bba815d458b31daf18d1f5e93fb9703377bb7c90b7d23a0b4f8989939391d78ec95e8afa623220b65e8a0dfd069cca2311a49b7a3de308627c8ace19b4c2bd17022fdc698a25bc6d5d8201f74e73;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b4ab5461eae834c3c738c2bd80b148b53ba30f09431e08d9a9c1b86218ff432521f475cb7ad264ef2fa168b900eff58eba97b2e99e9ed224b133471626bb09c2f1bc2f841388c7112b0608c63973;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h143a894c578d72755f9462675ced675e9d6424a53f13483284d76c19212791d6f6830fefb6bf4e32aee5741994d33364c4c753e29819464bca74b5da94c16091905039f6d66d8bd3e50256ed3f771;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h160d12a1c62ad8d53ffa02859e8e750e84060611a792df32f9c1c06bd5e5a91a0160e183dc46b31c0a488995a5a8d3c622e859adc3873c06716c8fa02cf995a83d749ddb322998cd4db3a641645de;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he0a3d50536d43be2f591ba8dad984c11a1c5bc240e451afd4bb7622c4b372d8c93fb0c2f44baf50b8ef75f0b8f208c0636dff1becb375432798b8618e8baecb894f3d65f1f00d388c5baa854c2db;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19c506dabb106ed0c1e4c664d89be0ca3aea5eee273a849fa1d9ebe7b4152591ea69b435ef14f1201cffdcb2f256d71c5b13122dbd1441f2391cfe87bc69b251acb6125749a2c761cdb847ee15a3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6adc9c1b13f4b15ff0735d1bd2dda84299a18e651bdd18511173e7060bc746f2df5282e13b2b9318219ecdcf67ee5e1fdca089144e42c2368a5a77d7528580bd91432e47fd6b19f7809d25f0a2fb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c75cc2bac0638df5a28c34816eb663b617f4fd5a1cf20cd8abc6745cc69618e554560de35959728c9a12bb5ebf16a335812bde353bfec6c3240549359661b261c01e1cca5ff2929336c372a6d428;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11c2255ea90436539d127fdbcc2724055a638a3e70ea9f6494c7bc396df3451f55af838b3973789558aed65ab0c6dadbe6e5498f215a24e4cceb8dea87e4b3e6542df4db883441fec02a825a5e34c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf5e17ca6db83fede65995611794c0318ee75e336a92fdd250efd597ca37daf87f5efc6291854a03b92cce7901067592f431b8bbc3a061403e9f797788d5ffc4834bbd5b43dd8e3ab513cb54392a2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4bf97cf066b30398e35d12fa8a5c5c57a18d78ce26057cb2113c66dcd372bd328ad7aebbdf66b6113b5280255a252a56f6e61fd34e9653f2f245c718b21e21f56181f755bfaa999d3c4e25e384e5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e707c25350a36f8e1d364d0f6a1a926c01934e8d2708ba87dde08e78b08230d568eb501ce1fae2425cee179a30da15a0b4e72dac6c6b146d0d39a6270583c686cdccfc0257fe6acc46a07bf04e32;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8ae97d9b0c92e5d97fcff9c9ec4828cec8073ae0938ceb858f3c8c4f58fa42e5a19742eb7593f222587ecc1367f8a288754e432f24cbbda7e983eede9aa3ce30c93464135ec8b4cb3a5f2b0478ca;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h729e8298ce1f165ea93d3bfceaf2a0cffd3a8f03df0bfd2395fa6f3c0d4692f31b4dcafa0e39a69239c582d1b5ac7a9ccc2ecaea0eee113cf11fca36c1ed7a35318e3ad2295f6e7d1b7770426707;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f64c879d9f94c34350f77bc2383c8fa686a1463dd2da9b61159a8d7fff2e85e986ad2be85d97f57c67224cda24103e3eab7562b74e1105f6da6ee529fc292f7cd72d772d574a2d281082a604f368;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9624e420167ff0761f8c011cb0172e9ec638a4a1a43cd64a83d07283362a1860334d75e68840969e3cc5e7d09bda772b499df458bfdaf8edc89d99ebd2340878a48adf80986650fa8234179ad55d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h125acd2817d032cf12eb708872b87dbff59db8d40b26a0cbb422435cf47b947b784bd94c71c01eee3e20f92e121a5944c4a8e43a68397af84d92e5490a61d32d83583801dec796dce77832d686027;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a521b9f1a03d93310bc078fd4ef3e8200668c60e52dce84685548783752dc7f4e1f813c9f73124590094c84c9cd079e2362ff166e3547e6ff0dbfa1a72464a5e95157d7986da0c009c9a697580b9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb7e6d6294626fc673304a18b353026c1254dd318670bc83b012b6049896bc7c29b849856ecb83c0a325f7c4338381cab939ac17fc840f9552768e401a436c82c2d0954fa4951bd9a5ba02156fa8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d3817d5bd13b5fae4b2b6f839acebece2a11023b7929332381c8c1438474da9e0b49f5a3efe60e9706cd0d621339823b602ac10504e9259bf9daf576172472f1f54b3a152e6e7c46c2669936d33f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11c1dbb34aa8f9eab8fca502f584b48e46dfaf3f6249eb58609641d52dc25fd73a0756591e1b6e8dd31bd23b8533392403236e864a9eae5311525044383733897cc031d6f65e6f15ee42a95cbe22d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfe2e54df0d750bfb29fb52dfc7832a1a8bbe94be38c659f28696a0f5d5b8410da62ca623ef101f530977a0ac12bfdcf3bdb89766db9775569677bdbad759819ef97c50d6f6a4a75081fa8b1b3017;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h106ad1c77c90ba3846f3c546273889bc07706d86c761ed1dfc8fe56afdb2caef4ed38e3c585efe98c061bd3bb7ecd97ea01e2d5662e33667b42eb6fc127dfd7df6262061f6933909dc8ecde8fb2ba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3b810986761a6577e11ba38782841c9825ab86843837bbdb88a613abf605980cfd2eb7390268f969c2b4d3f48807aa3a9d9083fe938721c7e0fbf715e524faaf9af886d3ba8fa03882f7fc944aa9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd234a5fa548f3360afda852e9271f8c4ade4607a87ab52e7231f06611a28b2ad8dd00e95ecc83b0240f9c7b1d93c9b559042125516ece5631b7780e05a098b16b67c195e23c4cd3b6f576cabcb11;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h82fdc9bd1ae32b7d5ac1049f9404a6c609cc24ec9471558a693784c7e25dc2ea915da7a8497c3832eacc13971b526c51edaa4d332dea82b9511abef8a7b45fe101d041718ff6c070affc963566cb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c9e1493e23b69345393b7c78e54e4af18e396cef3653bf075d5d24f6c8b5347e0e346b9c26693d0cac83c41fd788157d96002aee36407d310d72cf94ae4ee863cd06aaaed67eeae4be3c062cec84;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a70d5984f017ad09b5164101446f0dbeaf1dcf309988701d1d3a01deff2693305eaa862c3d0b89158c7a4e458a9e0c38708bf03a45ff6954fd83b6e1a0ba09bd54039b07699931fa8b81493212de;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hff50ac10a5c928f2d83bd0dec2236f05123198869db4bae7b41fa6af1d73e57e40d06dea65388d8b730530a0d575d74e70d2d80376641d66f4465b93f31335e4ddaec4b6d40214b565c3f762902f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h194df31d6064e50d8007eaf7760f57ad43cfdbb229289150ef3f7e541432ca7d49eb053452ad8820889584c9d1e5a98483d6eaf8da33e278df91f7ae5b74768d1f475a962996e998edef9b3b6b8ff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1749d259a3f61228e83c645afb0855392180641a6f59af3990abb4ba2c2ce9822438afd17bee6a7668f5e8a969503d6bb971cb5e9b9a82d6749bba10652c5d98d60295ff914da503d3174e2e0a186;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fec54b9eac6d1859476875046f66509f81c3d960b4d2b39daa035b9b86e7919815b24dd235f2240c83c32b00aa754e0e9e8a3e306983e04f50abe8a5d109e6efa9d922d36723c73b7dc828bf7371;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15c62b62506aad86c6d61df752ac4342919b9c68e04a565ad384e63f78c70742bcec5a2bf5783378b99623bd2bfbc829e4251a6b5703580714a91ca6ba4255a3a2da4d0bcd76741e40e830fff0666;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e63b744b65d026885481887a9049bec3b18ed01614e24ec738b664723bfd90d22e6c7ae1f360566609d62d7050a3395141fec717eb604a055331bde34f761cff5d12558e0183d0bae0a1228aa625;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1731437da3e6d16cf56fd7f9d2197ec37ebd1794bd40d70d9b1fd907acb8bb23753b88c18b932fec456b9fd68e47abf2323c465e2303fcf1fe3f26a031a184f182374056fe36ecc887a9f9b7dbe31;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2a3c8909f82a5140856f5bb92ed3a03df4b7cd0d66ab9e8ab005f7ce6f8a91654abb609491cee02bea2485e04ebd237754c297d7776a772a157a5f1a9c3e77d0f0aae55befb80c27348c9b056d4c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1145bec515f283e18a0a9be0f7df244eda760f8936c1ae8a6ce9cac4ceae79881c87ff96824b98ce54b80400b4f3805198334fd23276dcd28c50c9aacdfe192e8f3957dd17310ec2bb9c7fb60a332;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f14782eccbc9f560a9ff9de04c1d92f79b6ae11ba841e99a67dd720112983ff2c2c72e573b820d797ac67d5356a2dd04006614b5199ab0a82e693b367abbb9f872cbb6b6f93fc477af750e02f6fb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h182cd8276fadcbbf53a8b51eb0809677fbdb36f36a567abcdc40f0a66b7749d734067e13f7bbe4820a5ceb80cb6eb9afb74df4bc0d2fba818539dce1ed177ba97513564a9c108413c425fe6939335;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4a5c25a023b7422e1fce1e416e07c457b656985c6f82c03217dc52cc30cfc7ccbc9fdb9f3cff4b156891f64aec8afbb6a311600a68612a2a591eaed50855a07ea1029cbe6d3f8992f24f03fd9f62;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cf958e476c90eff329821067c737ec4c932e826a317d90c439af730ecedcdd2bb49d711780c0bed9676538fbc6fc8a38cbfd56b8b7a64d86156a1a34a1e7a78a2dcac0e59a63bb207e7b5a19ccf5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h48dda6732f58b18b4247b347406b4319f4bba139505ae915f2e5c646ffb0778a45a6cd8258461dc67d3658fbcfa065b0e6303323b6235451196bacc2526aa8f651c2d1713f9dbbec90de25d96343;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h82da04007fe417a9e54a93fde4b00bec8d89d8526edd7538b182e34222de8f291f864920e1196a971cbe7b9928efd20a5e765af10068bcd268bbee4af4a9956995a5b76c26cfb58705b5cb2ee9ae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ceedca06f95b934784120f0a00815fb72b350934361bb44050484f537f5dbc8be778a84764867f6d063906e24f431b07ffe09d88612752dd4d9f255b1225469f380e353ffd7221958e39eeca41b6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h154fc2a75424ede4c6fb914f01bf610032a0dffbae5d0000ca55bbf9c9bcfc83da3127ab3f99af8398c0614f1622d8d3a36109c911391456233ec89746147978a74804d085e3ec347eb4b62e5988d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6e33b8d149be49b20618a096477623af407888799b6f28250b04d46f2c63bb5947d2dc4bb820d0f4afdf9078f98dd5db485da4d400bebc03875dc848c4dd23a0e4b859837120840aacd912156ddc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc3388ba2ab2d2c4b7717ee8bdd42d54ad7e45e89fe58fe20acca180eadfa05cffca656649e77183a4926b0ea4669fcfbc45ff8d90c418bea934aa38a1f505db7f5647a56ca1b73ea6c799f1ad65c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7e06a4352f7a1e531d27227f21a3f4d31458d55cbec38c8642af3a79fcd93e612b779627eb729e5dad860ca37dad2f513012acb1f5963c1bf0ee05efd607b4feb010aca2b7e4e1e31f5623062072;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19e24b89629f3384cfe784bafb594cd326fdb1d1b39e7b037b97354826b46c950a3baec4924d70925cc26cde6196c5cb7fd6add2246692ca0f3e530790b165cc7ac6ef5459c937858490b2131e768;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha3e52431d86a08d3e32263da0a9ae2db656c0446bf11bd3860bf388bbfbfc66c68e9f569c65b225b8d871006f2edca3527807030dd0e093dac1332ffa7730dfb6ddc1eef2279aff08fa17ecb7c13;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc883eda32a48e92e77531cba405cc64ea6ec5921c5ed21802ca82b51d409eb8dd7fd7488fda6208c3aa0abada87d6ab705914f7841a0a787a8d11caa85d9c0cd7b1d5960de39489eab44091f4150;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5c177e06b06d3bb4c7e2bc7fe630a1d92ef45754878311d2b8d0a5878c1f4f71b7dc58946fd799a095fd4e1c51ec7cc58347484c3edb84a3e3cd66dc1979d0878a44c284b2ed7cc40fe5963d71a0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd1503529e2d796c5f180f5a48a101d95c4b9c217f589748717758dc9b426189e2d055b952307abff857318013fdd887a58914ab421413057e74aae37612c399fe482f4a1dde306b82eef3c1b2a40;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd47f0d959a1435b1f5409aadf84084732b25bb00267038a718d2c165a2e7330470b6116e830c09bbc9b25410b7bd7e4ef68787a5416a044a6feec5c726f31e9a628c710d5b6fc4e5d6159f893786;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc527584045a2de702fe430a1c054fa8501c87cf8afc168b5a2704f4c0b8903b26146f22cd952d0ccec3710737b593422dbd08616af1e4959c6d6a7e1e9c9b45135e7152336d71fc20420d5af798b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hafbcefd8e8af3b82c96bc8ff007a959785cccbb5f8f4bace527a8b3881178f268437f0b7f595bc455c01076b412f348d4939dea8e32af8d44d94e8927021597840625359b7ecb77b079f25a94be4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1211348892912c350f76ae5b6334f3b9dcdde234922ab6063d78e2a4228bf35e8944d82ad12a69ba26bd8bf2d7a98a9b9e0ddfe24e9237b91f19ea428c0b78108d89f9661bfa6f3bd8a5972730d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h69e63b786109f80944c0fcc42f2a4ca84cc1e06962a8235ca99b58be03092fc0372a479b98212f3752cfe1bd8ac3063f7a8ae211146d423d3ebf0d21f3e041c676f1c5ddd21afc3f2fe57b0b6274;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2a48e30dd3933cf4b9772d9f3bec8fe5922dff105096c448531290dff17184cd745913f987bbf994fcfde9c79b13c2c55b2d5acb123211217884fb94dc236c01e1adbabcc18fe48083f2fde9b7d3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h334f3822749b44b7c8d0bc439072b7195e040d2a8ffd28355c370051a61029aaa4565ef30735f466b0ec0ac5b62fbef3bd488a48965295d94934548e7f14df4f2f15dce9921bb6441563d2ea3a21;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10332fa81d551af73b24ded442c9577e0fbb1d82cbd0d8050dba0ca41b95039a692b1fd8c5b136cf8122fb09196c6d24aed465c9c192b6a5d0a561e955790a2fec5e7806641a82a13e61105faddf2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h93b4d4ca18839af5c82523ae3a49b711ea2aa6ab316b08cb9c7601d8aeadea2bc94049657151e1cd7f2113b8fddfd8b47764102feff04f9a37d7512600d3d1d0ffda7de1ecb5d8ee887a8e512090;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2d237c13aa424952cac07037dce24d006920a4c7600ff02c1a8d8d019b71707108f62da3adab2f4e14e5ffd74c1f4161424fff7ae198648ad694e7200dc429f871beba7fcaae05b9306e2b932a31;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h51100a3e6be6371bb9e2fcb45830e204443d826666f18fa1c6c336bdaff8c12c1f87906d3cfa903f8a3edbef23e5de2461644b55aeb80b4e277949d67556ca532e87243833b02e0a8164bd53f5ee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h328f9e7219903c708fed3cd1990f2f5992f23cd7fab68ead343005c06825e1f5ec1b0631b20d0dafe7a92fe434687e85307e31f86f7858e1eeb378fbc15f6d3c26b8f91bfe959e5365198f897b11;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h199514a162bb5f7f55633aadb7f05650e01d5055f27ac2176f88037ed1c1e38abca3633e8aa65b381dd27e8d59360ccaf61eb9e3df5b23d269468e307d719e5aa336b5e70b5a04a91341f7bd5233;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7c64ca5873429d772a135f01ebbee16c2f63a523ffe9725cc59f4511dc3a0a13ff6a467b4ce4461d456affeafbb4e7ef7158f9650cd608eb6c4847ff227e68696c8f977018e25430f9cd881e1feb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cfe66829e9146c0d2d369e23d1d0473f7a88d5cfea78e278c074ccdf9183f205132680f2d1d9d02d46feb51dd607f84fd29ea34074d1505e397456e01c14d97f7523ec961ef1a36cfe0d2402ceba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd26962c199cd45371ef0219946ef3465a95fd85409c8348e06da1d04b772e7edef1bcb1b07f0f0ab4fac0a34a3fa87c0d15059464186bb007b3a4be1029a079df3b0fb54535afcfe563407cbe2bd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1afa0b8ffc6ce7e245f18c75eeccc92118a17d8261a67c8212383683287bdbb3aea3eacbe4666edda4279821422f520883117a0941a2d361b5f9f4ee50a52b8cfab47d9b2cc392da6f2adc0239d61;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hac9f3ca250bad9b63f879b0da6c1307c8b420aeeb5bc9bf45418d33563f753a7027793fd8ea80ec565f2c5b793fd791926b7d57b5f6ba5397cc7b6468fdb92c1fb1962563a32891f5a63b36327d8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b71a8ec5ec8c369f828db2452995ab1c814f149989dd5353f395cad68ca6b36da305595a1de8379e2629815f19eb653d08170ab4a41d600d3702a4fa1044b9e206cb31c9ceabfabf0d64552b8957;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a3db22de5eddfc9c681374eb2f746c2d51e0f566a4da060661ba8b8d2fa2529008cbc64527ecfa7c6033085f16e8db8412ea45778fd8187efa8682e0e4b98ff32038b2092e3ca87ebb34216f13a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17863274499f29a40f074b57d9a96ebad3b6cb81083f99865f730d52f4e22cb1f769b8a2c8c8b0e47c52360710f5f07473ebbe5f512f17093024b029fbf3259e298a1b62d9d0bac88e4a393d5aca8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11a72730bd3f2d87e873c9075e610b3fcaf37cc7d1edf305421750364e908f77f919ac5234448e0b735a36bee2d44b53e131dd44281ffca6ded5ccf6430e862a8bd115a9cbf842f3e75301b7aae2e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h29edc0d7cb1ff6814253accb91816674389212b606dd6a2a28a9418d2348a7f9497cae4074f97e96cec2c0ccf5a445401b15ac4e74cba6f5648f46b47298ff4294efaee16f9ccc63c1f507a6c442;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h159c1df0c2d5b8d50b04e0988b8949039e8e39e152323e243fd48832e145a898b2c647bdc38fd812ea25f27d0aab30935b8a363a6d1a744aeeec9fc49cccbc4bd20bf99520a9740c2abf0d7e2352b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e21a130d3efe9511f1be9cd5838fbd793dd989bbdf36ce2f5090b71ef0121593958cd753c2178a56f99902ada1893299e9e5fae9dd0c027c3d50bfc6abcd0763db0c7a4d39043bcb2b9eb14cb142;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13cd33b7e0b0c9208f96784c0faaf55cca2ec9a59beafab68399d9fdf0d5026cb7f79a34bfda50d3598eac9bf6713cfaa6991713488adbffb7ec64759990a01dda857cac0c5a0cef88e62607483bc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h612b95d1993c0ea3238be326ae2f34b1e2fa0624978127f3b7163f2e48ac9a94fe61d15fee5012757a7f33c6173ee9c6a3263350849b5b4a8abb52a5d53f2a6fd93b3ca3f043f4ba43e60f549089;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd8fa90a55dba39e7322dcd48978cf1987eed8e5567207a119365071224342741a053bbd5dcdb40cc063b6ca436a07d72af4dbe29ab880c627e8b528dfb6b1d2f1f52a01d5ed3d92c49d0ce84e0d3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h131cb6f705338eb1024a097aa14eb51fa3a6a5fc594af1c774e4cf2f14556b54e7ab8e37ca72d83af280b0719bac9f752b58296a7f234c4d2f867f21965d036af078386bf3de49e70e683cb9926a6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17192969b2af21f2a3ffcb5bf5310402d227b5d24a29fe314f2ab0f0b65f8e6e6a8ffd4a90561b42e859c0f91c3c72f78c04e443a7c439c371cfe9d59bb377e7d4d32a632435e0533b200c4acff49;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h69b2131c832256798d364caff5d513d26656342219ecff9c486457be5ced6c4e6741c4d523b511662170a21efa774dc5d7202c09a3d5671b71381e361da57c8202a36a80ef099759f0d1bc55561f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11b25767aab7c2c575b8e21efdc9a84feb0feacd1d79931e0ea28063213c20efba528c9bbc3b90e8784f2e58620212ff1d5f11ca73612baee3fb74268672eb8e3db494610bde50fcf8a11a6de74b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbda69ee16e9845651ba51be3d9753d67ad6f61f270c7552e545443cc51c612991711555415a4d539572cdc160a959dea78440637085a7adfba7181cf85e7e291ec2aa0b08a0bf2b08f68f349dcae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1de3f463f2e805647fdd5d61938c73b47f724b8042552ab4458291cb4c36620639c8a4ff78fe6de9ef98a373d9c4eea32b4b06ac470aaa75f5320c76dababb334709061b1635e19d8503d9be8d43;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e421b66a5adca8ff483512ce431d72eeeb579379573e34811321bb18198fc32ddaf80ac80d5b9b6cec8ffddeae96d9358df5020429d6c45453877d08c87220eef3c360ed37cff9087b2c07d9a360;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha81dd246ee00163bb040dbcb4ceddccabe7bc2970e5680d4df42a1bb44a1b2783f982ab9792308b9b808d2f5e51cfd33eb0e6a1fa6d45d07fa39443a722a1a7c0a81e5c07d83071fdd0e5c4d041e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10c96f09f12ce3725fc03c78ebfcc49a04ea4b65c2a98f54924dc2f139b21ad1ffb7d191b9e94a05af17bccb1be55e1ccfcc92816a5bf57f2340b1b050cad9b07f7c39c540bce86d6fc192c944532;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10442bbb31a71393783ea1edbdf5b96498d70e267a4e3c17620bf300c87daaeb43a63a4b2a680f91f15850948ba3f7e0c3860d46bad21915299f7f7a94fff2285a6ff47de33d61ed39bb403898d5e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12f20d7ee86395c8221d1d36b371a55300845271afbab20bb869cb160094515db20addf62a29d9ecebc092deb92dd7dcac211f7de9091026d10903bb4d778265995b9e9a4457c8fac99fbb2aa664f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c08048e02b414c551e02821c0c4d4cc6dc98c4a2b6a0f72647561c35ae7f63a35baf8fb5cb04977f8142478aca5aebea51124fb0454c5291702af48d558c91246ea95670fa894bac19a873d4e986;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf4a4290f4ee162512d059c34f817aa64c9e8b9266ada9a8ba4579fb38928fdf13db83b85332d188110e35fa25fed716321cc058790942291cb78f750f49ecc8daef28689d5fcb6cd9ae2ca1a28bc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h239ab2aca3846e81f1554ae864c3edca1cad7b46c113f77bb78ab2bd11ef2705001d1058d77c36c289cdd4ffdeba07775f05c247aa87461baadbba2d5f0db53ed823977207b09d9d17ae0423a378;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a517b0b081781b883d461ec2ae8ac125461a317ee2838fcc9b3e78d2023e6c58d54bdf3db39b962dcbe73310ee84800eda5ae14b009351df91f16a231d452cec6b0a3bdf159cddf5b469d70f899c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15fd7d5080509c83ac7f1418a705940ea13e6c0ee83d93b6fb33edbab55048646d0498480f3365ea2f7082514ef4c0dcd092b1c72709e0f278899fabe25939110edb5dc8bfab9b53ce915db14a6ca;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c8f9d978a1862dd78006d8ff707f7872547bbdab67db3f7cb124b88bf3e48d1d79ea4e46ff3c561fed503167ddb065eb555aa152f5347536973551629cb0771f5f0af56e09ca7cdcae0d49028988;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f9c270c1bcd33e3a60e94ea021ecb1ba0a540fc712f8264dd959fa2aaa43148bc12f7e745733793226bfcdc69d11dda35eb4572e354737f9e0ce5f53c29f72cce3729afc387069532a7a694e43f6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1abc8a7f46844263ea6eefaf720f9aedcf100954b02714677baf134e0f74f44f42ae4436e5cc0f58aaedfbf54867684bd3ea8bcf4b4cecfb6b2bbb74f9061e213c741ea95eb55fb47cb5f587e5c7f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h149dcfda24131d060f417e8ce36dc5448847538d01a4fa7b2fdc6eaa84bbde9d9fd7486540205cb91974775c01c6e1d059c3d7f9c2971daeeb5008e2b44e065df07b23a718a4c5144bc52cf91dc26;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd1f6437ea5ea68d9919d66a492e2e669b12c0b35982af912c93738f3af970f0f63249146d9c48a6d4d92aad02703b911c1f1026936a66f398c3c9e8c59e9bb394798dd31002dae884624f85851;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h94e1c09fe0ad19644f1932f83bfa04f13a20190167dff9b34e1ec049c5b2922f8828ee2eabd6755e63f6e9d3e594cc651bb5e32e98ef12b126ed2de67f6c9fc7e04ef97b23f26560ec46bb3190f3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h97943ef19e163c711d407dd0d2269bbfec9ccf05c4088fd2e19fa97e3ac3cba661e70694815fd7ffc0582e413e98910eb973ea75402a439a1d207f3d0744ee4e9cf515f0d3af05950ded5f57cefc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5b722e0f2f3cee1915dad1ca9fc1745c658602cefba92baf69f10ba743007d21180644b1a0348748cb7f8ecc4e4fe4683a05440b1ee1bd858d2ff24d816b4aad2224528e77847672659da6168761;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d0a6a55cb5cc09b4939df27cc3b335bfea8c1e8031fbfc4197d9aa485ac5977e846d84746f299213431e140ae2f603401ccfa2b6f926c3ba19cb3cd71b411c17f004eb8a6dd87ff8eb20e8626429;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h56fce6ceaca840fb52de98156855324c17961fd9837403ec8e09d8ccf11305e6c553d5a9b9e4b92f06730003e30f647fee236c8e6540cc3c496a72ab31a16ebd33ba8a0738a7fd350067a6ae6229;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h136ac1dccb772b827c31bfc55783cefd79da8c03a94fd96bf50c956c43c30f0899663837eb0721eb5a06d54d99a69a9ed1f3da197e0178a5dde734c10e0df462a05540c0e5b07515ce1d1637ecbe8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h40b728578513bbf3dd1125fe109f581a04ad404d340e94185eb530d6725a5a16b747b900187ba3aabe0d473107247ed4d55a275d19a840714635f7fd5ac2675ed2fce97901bb260ddf7818c35e72;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h546c68ac0e7ac6889ff668f1d2623503c3067608b2386b27b2044d8b257b3140b1751157344ee7e79ff68b204330ccade6f4a1c3b45ce9058c05d10ff5cae4f22cbb7b31585a4b06f808af25ed4a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4e446f88549a6de5a7b7aac2a8ad394168efdba8c3e4152fcc6c67d400a3d47afb2e6cbb3e5435259a667ddac947dbc50e14b939d7596ed76972b589cd8e1aa7a771ee0c515c96849d94f6cbc1c7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce74a3909d38b60d55ead1db4b53b444f86ace9e10ee73510c38dfbd1efb3851b2ff4a54c7a547bfade46196577be737709fbd541b74f589ca70cbe94a32d81c816ceb7408dcb3402e90ffa27ba2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd91d4954027a98181c7496f3f7cfb923aaaa13f664c526e1867c1a26c756296a00837dc9d8b58b3cb286302ce3c0003f4811e5a648187d1deef7fb45488418f07c25b6b7a0810085b92ab861150d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h148b581b411787696121bcc40b853d6432c67be999b01d4d6ed58640a1563708b0ffa5f080441df450753e7766332e443a0ba3ec928441197f66f4e714057d1c4ad58caac5ab15857b2c3867ec895;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbfe50ac26cb85d4da5dcfee9cea0cd984746a838d339d3f78d08817d40353e8ddcc60051cafb557ba7a33c53fa71f554e3625c32ad279eae84b54cbcee468d4f7d9987ab63cd1d75df427ce41bf2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6661a7b0791659c50bd7c02b5aa43e41bf7f341ffacb8e1de36d541e2f23f290b0360502471122c87ae11e0779d93037ea2bbaece7120b88d09d3c430e582da99e5f155dae75e14e8222f75d37e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1734bb927a9ddde8eb0710bdb3738d4485ef9884b2bf800e48f11f5fecb64fab4f19fcfd338a84bcbbf6624671b1fade68ddbc91705038ee31d9efb3dbaeba0f1d12203fb037de9e5fe37bc796abe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h236fd4008d84b9e97c7148082aedecfd3b5de2af7375e907f41687b745de8924a1d98d2dae664dd9f12365b664ba8147767243e6fdac40f3f73eaeb2bc4f109976e5111694201e6b694b8ff1b892;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h593cb6a327dfd5f0db8d61253f91022ec808e39c907e26107a685c9781bc02ee2530cb89e6ee9f95b92f35a4727303dd1d7fd92eb3dab5109906d2fc44ce6f84aafdc249002e25f462c1f6d80e06;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbbedc9b1d953e92fdbf75d5436be3df720e7dc5404d1b66fa6454a412b2cb1f719f32a35cbac024a6694918efa6650812b12db709033ac7f868fb2c387ba1251612fab5c5542336d07ddb3da1bb4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11ca46dc118055cda359f578735f41dae50e07a3f47aceee4bbcbd26c3882b62be47f5b80de249ee6020a75d8f1a1328400fedbcfb16b5e8aa8830ee48bc92ccac7901817f2aac4ddecf7c6eab220;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4684f597d2f4e1f5606c5b41fdd6e37181bd94d3098ff49c8a943502aae14a557712626269c5c6a1d6ee11b4d89223650e22ac04c5e070ab6550ad9ca20fc17c8264a7a77f1aa5535f1a3e4fdf40;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16c291ef5ff16fe97592d1cf9fe1868a0f62033ae4438e13bcde7372792085103b3e56568362e0b4abd11ea1ea321d7b0946472754fa26211ba282f66a48cf430a60c45e7f8aac94b804e59699c83;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fdb189a5cd7358914ac899166a7d9d1380f1c8e11375681aa9676604337b8f2eae3beb56ab7e3e6bbd7e41a9d7f696ab2be162ce2cbd186f5e985b133b0bb16497a494326cd07eaf5b2706808ccf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb1dabb60c2a4378acfbd7c2ca4da4b6d832ebad494c49507b58254b5c069b588ede9554fe5193bd3bff3b1e0fb423479e0a391fecea73be55860ed94a776a4164d3f1ffb9ecef0b14b81255b188c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a21b6bd45fbe9fb7b25e0060985902081ace5482cfe65b98a8f1f45c5e46402ebd3f0f54767f6de8f742f1481ae9693e2c5e062e8ae80d98fcf56171b209d1e171bbe860bc6cc18387b04968e533;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1df1d0ca2ab1f37aa61c838f0feec23ea02448a015f7eb0e5c600c614e08b209cc4e5b2479b089d2512eaee1314eeefc4601c76e0cfa9cfe4710054e471a36f287147875824e59d89994e1284a8a0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haa6798774cc5932e08113705325fc9a72ad27006097dbf1ebaf5becb11b3819f694c43acf77d2bf3d1d99f9070efd6bd2841922da969b73595a3d05e2e7ac1c9766f27853ae55ff43b82dafc1be4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1745efb80d9b618f5b7893e2b4e8d95b22eda721f86ce1c3f55bfdab8f26e8b1bb1cd2f2abab76b5bccd38055404db1769a26ae10a554cddbce80c1fc36272dcd9f771961cd4ccf6c4ae57bf7e3e7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h46a5407541c7c5baaa0f2cb09f51ec9c8dd26cbb7657286d16c68cc0c27fefdec174976a65c3118e6deb58fc09c007590bbf255dd3868bb2ec735fc2e76d4a8f4c44611e9198ed26a8c92bfff1b8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h191280a1bf0a9d05601517d89e8ccccb5b44a94728d99128a8d45cee6171345108d665a885b3307f12ee7b8ab3c05c946d350298e6e0f616593caeb392e3e82893b6df019ae0d760ddd8977bafee2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf80cb31ce5d66218d30e457ff1dcb9f4b8ab0fc738b9e130c03d79c5cbbe00ba7066e7dc0104547d80f0c4d745c1b0ad1ea007d690c50a6111d63542fd5a19baf175194812ca34eca96baaec7b78;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h98aa97dc91a36b234847541d4489aae575a15e91872342ee01d06732be073f8f8a66bcd185c0cf8eff3373b40d75473e64a94964346f5b6ba2f24548fc53f670ed739418ebe91a44865d942e28f8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4799e455e16b42f1455aed87b9d841a543be1a469d55c4d969aad162655be6670f9a3f26207a0f7c3d5a68a3589b004763b4b6a422e98f039727e12fed60bc9ff736f508bbbe010c2238fd6f27cb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18087c00c88331cfd575f3770fd63ef4606fe2c5f9f2fb6f6ecfba6be67f4539e184f2c79d055b2b10a140851da3ffa44e09f089637dd49e8795c0eba96ecc66038341270208bdda0275331d1996c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11b90d06f690325c018c7f44f6b0501e51f7725524c5d9596d105d7e629a1c825563dff1f57f4dd659a0018b06e20397f0901cf62fdebacf07546a581d2864ad22d49458a1d70126203da2ef79de4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1ca764c50377b6026615a3d951b7a1606b1331e72462f2c7fb2da98f599003a8cce51ed2b4d638da8135492e1707c92406015095ac1b52e29e44a898348a0a115b2093a1899b66178d6be926e7b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b423f16a59c7b08118fa73ea9306d95c01bf5cabf426cad7f7799bb364be8783db070942c8eb23072ef8c7c5d4dc988cd2922e51b8039901b7e5241b301497e090e982a4324a7e3028969147d005;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h148f13309f499d5ad0512761ed4e9cf0f26485f143234f7f57f229051fcd961e391553333d071bbbfb1201aaf00793510732c8333b6c977c6277702eb809b07dec4390e5a7847977086cb05bdb189;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb4601f86da64c3f6cdb35fd189581266138d44d0b64c223defd90df7a662dbc06516e5c4d93e8c3c0ae62445ed068b41c7d4cd317250a5476b6e0f22d128a73bfc3c40f984291d42fbf6c9634be9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb82506bbc83ee47f5c42756c3e98edf48f9f946670c5d50cd4856af413e5e6991367d1870b2223140beddc9b9885e9a1d58dd9f9281f762d862a8422e90b92e40b2629d228088b9463c4b9a4580;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10cafe006fdc64dfb94d6100a58711373991fce63234573547b78b1223d7207e55e6f03fce3523d9516038ea5ddd268c9ba09aa273c50a8fd1637e110d2937c76a78a2427a37457c784277e47eb30;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h46e16823bfe20aefeb7e883a1edde39986a212f98f947e34133d552ba2567df55f87b161bdf2250a502734c42ac966b1c9c16858135179a1ba43eb1b1413daef9fea2c14f21153bc625fe5397d86;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h177dca48cc2bff2ad9a5eb745a0ae88ba8bf63e6a070926733e9a747298491a5692a371150122bb2ff46d00b09a2c7de3181e08e1749a89a19f77b0bbe64295551d8d3f448dae57058f16b24f0287;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc2b85cd05f53b4cce126bd48462eac1903ee03049a6fd6d1baf1620630e370a4f6e16f024f17aaba090eb35e798387904be4aac6890489d3293685ab194de222ac42fed04a667a58400c71adf82;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17ad2a4ee1286d5792875f91047bcbd8e4c5d51ab8d62c18e81c8d443bd6db3838f65a97c985008efe54470f7b6a9cf0e8817ef644b5a98867ef09f4466b7a6135ae7018847f287c1e4fcbd7a156e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h63f8e5d7b71d9efcd821d476a48329c3a6c424888ef37cdba633f40b68a5b04bed2827f1e5de322fb2ec8f9abfb0b4f88ec4fc3361a3ec5122f7fc6a3edd1452c29200990cc8cb6db388855273d8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h30ee746bfdd97fe887f9f82538619e99ea99e61bf262c76498fd0f9c43384a17eece3c41077fca428e5111fcaf54246ee814a04d2c9904b332985c34e98953b8e921b3acf16b8d6010c1c5b86812;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h130be30d183c6662922268c356a78fbfb6856de31aa5bedd4d8325d3769afb68bff4c99d54861bd005b7a09897eeb738db038f1589b6e9780b1f503392e1ee33ac274ab7583c4c2c1059f98cd9501;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1014b6e774dffaf1073f39f4c3206d054005b16132c9a19c8b8817ac4ceaf3e183f35c55829f7b4ce23ee235eb345f2f2d4ab4f0005d3b374cf21a933628d77a9d20e9e29a638b989a30f20d6acf5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b0903a6391acaf9bddc72360f63ed2fab9b54266be0af96da582a946b444ed2b510f6a6590400aec42d3de75fdc27863cc013cb402c7992e6cbdfdabae58f253e8dd9cd1434b8244a95cdc45a0bc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b4e685a2407c5086d4c46b408b0cce07aaef37cc496dfd83e08c349d2875ad5bf1a9ed91762a2c40074d7524e0aceffdabb33115c84098992a16bfa9702a46a5d0855f955a1208f70e8280acdbb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aa8a7716505e78674a90fc6e160ff07574d7052ffffd27d1d73d4881615bb41e936ffe00fb1c223d7ff13e517f90bb10392aed42b06e7184500347107549168feb1174a0b5abff59b434ad3a223a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19b414766b8f92ff1e332250cc70c6d6cc52b543f9c2d2b444dd9a7dc5b2b5f2305cf8a645ce6a885eeae2b2f907fb40b00cfc1019a751c444773f396eb767d231d47d9b14d74b0b471d2227fe238;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc8313e2c5025b05b77b24633aaf4fe8edd7663ed18eef28ec270571353176be9f605271e577f8847e768d081329f41927d48cbeb20c35ecb9803c30108b52d4ae8c41878aa3cc664da500f058fb2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11a6ea638fb432c44770ef91adb62d088304e51370d087fb26258e924d1146c6dc571509aba1b92edfa76ede5b79540d06ef6aa58bd1b5b54ba3402ed9a8cb58d5778802487b3a8fe4288589f74ff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17968c53a2da7eef4176de2732e96fbfc585a0e8a1063d4110ae5f49bde9629edc4e4fddfc6abf7b50a641ee7012b2f463c900bf5d343a9ff1d7c7486034a77eae4fecc2ddf4b74a4539c7c95d378;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h79bcd9cc7a2279dfb446f62623f7e00f5a2e2df6ecb758761c8f60f7603c0169444df8b87286facc4ad7e89b3dface810a80bdbd9bad57de551a5dec9eb3eb53a5de81d8460d9198533de3ce4be6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ed63b5115c3f8935bd130ed74d8d705caa04e6e2daa8cb4e45baa60e4a746817fe3309ae93192b2b777ac516eedb11ac29d930e17d359eccdf0e7a5d0f4e7d643918043f26812a27a48203d611;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbb42cdbe0a31340da8315fe3d1293ec9fa6725557a3c2e7f06f399667fe0779070f9b81c89f62ae8642ecb864484326842be9d1d9ce8b33cc1194cb048bb982c9f819de03e4c3df9032acec6d3cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc3aa27717db1a4a6a30dfd2529d1e862b73a03c56f804cdbae5faf072ccd692c1c66668a056dc91fa5cfb0d64e5dbcf7ce196bf59b4e5cc9408bb0c5447469ac37ccb0cd98754ffdd190cd33b6fa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h458bc59250bbf5adcbefd65d8bc63f93a2d6f16a82fc50721d46e2a86045754159509fe3ae6dd34ecde32d167601137769bd70538656a110196c7f700ff15ea4b3a47491bd5ac75ee1ce7595e495;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcdc3191ccd8659a84712f63216da440c2bff2a57dcb260bae1e9735043e93f9da5f1f23adc897e04ce0eb5077b1a2fec0e97240a46ba11933d80b3b791c2826c03610b59a53d9003e7ce1b01418b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c1f4a3875cfa92a1fe61cb67a7ff0c5a9deda951f602959c98e4a694e7d75bb00f49bf164b005b70d89fb8c389736600ebd8fd3171fa8d6683cbe7b251ccb10d7510cd68581c0822ee0c9c5172c1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9f1c705aad2eb46dca624ae597adfd11fbc1d0e0b3ab11fd7a5dbd1489e845320ce3dd5660b60695b401b0d1676453f8861c20e3d6f9f6d9c3b5baf5b42a8bf1f6da0bb0eb803dcb38d6bceb47b0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7a89ae880c018165b98ab09414d7cd3896ac984c1a281194e43057ed44967d78ecf18a3d77310cdda6ac4a19b8fae85b5fa8d1dd34e9ddc8298bc042d6df954a50e81dd865069a144522c024f35f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h162d6df1cf093b323eb3f44cde860036ffa6e7964768732ae24e320cc0f864d1968268cb390c54d8679caf23c5695213f52d7fc5c4007db465b8c149c246fa945c7761ad62680b9c59ce38259c1dd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h182e0d92f2552f36c0e1b75e239c185b72703f368a45655e1ed7c265c210a6b943791ad3f6db03f9b4a494f2d8076bfdae668c7b552ecc245285ec1527926c3a6ecd88bbdc80cbecbff245d5deadb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h34d35a854fbb59c7a5ff6dbc534ccb8cdbbb4af293b2da3ea81b6662cd016d75a3d47bf1f04aee79e200967bfeab8538e21c46e2ee9cd37b91e2c711b1dfe3816981f42fbf32c5176c8cee1c5c7b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16800c7f8b169ba572273c7f822a80fd2a5e6bb8c36d7ed37ec65c9dbcf08054a07c7c77b568bf46fa73165f197231c33eb5304fb433f2d0a6a766b7d1bd1706b81572a7aeb97113e87549d5a8220;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7295233b9ff4d29a608acd122fc211d268e7ca43daa97f95938415897d7281cd52071adbabe9c028490cc2b967841265bde330ca55fe3fde76c5134db8a4bf68edd19ee54a56c15d10fce8b0cad7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf289134990e9f75ed79e683b625cd86a14912096b0324ba3315fdebc8176981ba0874d7e95982969af30d0ea7de9f1c0eace444e45c42abca458828c986b450d0da7bbf5be82c7999e13ecee1665;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd48208b1333ad63d187bcfab3c91f1fb34de35c59516136fc2b6182cfa1638329528ed1805329e26607875200a2f10aa46e3802c1fcc986d3a7664dd7a58795751f88ec808dea91f75ea4927c65c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc6cca235073630cd1efd3cd159519cc0f4b488a0084165c5d674317152be1bbbe2532c9d5b39940c75ab87cba5ae3e9f43533f2552d4b3fdd1375c6ff05464fcd3151259866cb244bdba19e1c62e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e8d5688ed6f0ee46e10e7b6ab2352ce0a69984a828120c505b49482ae7edaa4782583bf55e1c18f0ba25db217ee3b2a19ac12f3295a83a0b3a5928a01bd88a73a4ead83e478dfa6c4c0450a6c87;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2e9e94beedbc9ab1269882e92de2a227252c6906e5b8a8b0357cce42c4a6f09588f3ca010c81a0fd546b1125f1b6635b8339048cae8bff2d78d6003c2adaa3b24892ce13916b667b9a77cc1ee69a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha6a28f2daae6999a2c659a1b89ae185f7ff80c7abc554e90571206e278dfb1ebde330afb4781f5739ef45ffa011f87843090b6820ac7697214f7dcb66c78afabdf5cc5b1fa38727a9df4beced30e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ac16947bcef083e4129b547650bade83f4b383db82ac880fbb72b8896f55a7dfdf03bedc96654f44f449f68ecf31a49c92765db4869096a74b54d7b4a8e13b982ff1456cab1bcfa157e3aea912c9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h68fa4ed868b81452bd2b51c0d130322e472fe573a2e0e03897554f3bbbb8ae814c64935cee98d02b9e92af132c038bf95ed907a284cbc82bafce049c2ff604d6084b0d4d064f568568b424757991;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h66c465221ef71c36855356a0f291c340ee9a527aca34d2e9cfdff731a69f2b191c2187589a0d19ba7bb43add951444dc19ea0a3ead4c81cde99a6661c6beb5a3639ff72c42fb4655c2766ebaf5ae;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b7730a6716de545be1f1f3327384930b1d29fc5e6590b2f63c3a100166e4b099b456058243d1b461e5a9795de5d45b50f2073ff1ef09275adf23b8b4d5cc8522e413799809b20d9b08a6775e5268;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ae6baac9f4967fe9688bc4292dd5e7a1971dade74c3b315173db285b2f5016197ff621e159bee14e6402bcaf4ba86af092e65cf1fb794f27e1bee0c172f53953e376f3e057695e786405cbe9114;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18def6483fbb2a1c8d75a69765ea79a8cd3b7f0ed880185c81ae436d69bf47804e4f5d8847d76608a1bd206d0f6d5915d31fac89ffad12f8f61752de8f73247326d251ce29dbaf238e61bbb079f6b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f2df6e2379dd6443720d6b7a25ae09044db5ddf8f1cdfe616dd700dac5a61bbca2e790bef35703b264a9df84ca2b0b457ca09f33d4214abeef3e3da4665df0d2e26bbdf62834670a118a279a93f7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c0cd28a4b081e4312a67033bc98dbd766c7732fa15d6a3a43f8f8e37918cfa084c1227d5f2e115a58a17686075969c3c45f0986230b504b68f41cb233bef83b6316d470ff22bd3f6b58b505564bb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha51186867fac6aa8037bf37a39a8c66f83905aa127cde603eead99fb48b69aa218075080398a76a380b841344544b762b50c5cc7a20be14d3514c339152bacd61b17679e764f6361c9b290c80524;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fe3946b1ff121a182b20eb023d737cf3ba3a458ae83cecd3ea837655390a02528b0294783ee8e1d4bda67855df13ca997cea0de98ecf11f4b5b819c747ee7a41530996f3bc0056baaac640b1b8b4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h92fcc06dc22ddace509088d4724e3995bbbcd31dde74488c775a9d3e98c4c93fcc6056daf225b2777dd16053992c33d13f3915bdebc738dc42288aac8d89c450ac3b60d43e1672c383cf2e34db8f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14d3d47ba5b426ac04e0873f3bf3b45bd29c3e73441faa6352167604cfd6b7d1a83fa878ead8f29eb3709f774d83afd9d0770ff9318a81785eafe30d02c4f27af165937110fd0e0f220c1879cde56;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfe7884684ea6760121092dddf2c7d74511bf2d23d2dea99cc5157bd3772fbb9c2c75a7fc4853bb364784d2b4046d01656166068deca529f3a56cfd3835a526f57ecf5eb58114b1db93b41e9bbbaf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd755e6e5b83317b270e302bf0058b2bd14febc348e73b057cb9016ef03c9358827516b1196c56d9eef2c4f373006fc7f490e12370e56bba666863af54763b9728ba68e67b73588f83b6cf0f28fed;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h121ea0492fd6b720130b93fd2d17ff641c57a031be9ac800b7d9b6eed0146854b54633b6c09f55bcdc868ada66d5ea3cdb05938935dc31de6aa30f5efa793e0fa0219e1c92b0ec48648c164346503;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7b497748cd452590b30a52c6fe15709e319c60c2c2e3582e88f98d3734be0776c89fa5de281dbc103bf41c46b5b4cf414e5783ab637a75c670dc172a9b7afc6dea4308bef3d933d6c118914d4174;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1537fa0f9ee016a95ee056c8f9b982ddae10533cb6c24484c3a25b3497ce5cfe96a1a7219ff9c067dd2ec91a40a179705f1082fbd9f835d3677db0dd487abb85c6b1849281e2f1b831698bcb1c024;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3b1395da94b57fb52b88bf7d40c0c5210415a56012fe72147c07642328c448bbdd95cb884df10a5a528c02e588cf2554502eed11e81c09e61669891fcd9ae4be807b4285a27579b394b8c0d2952a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14c57a0dbecd3c4f447cf7fc9c8e0981f7b07d393b400655cee1d9cc51e07a8d3ec6dfee6c5113d98766384bbfd56a67f65721c082fca3fb0abc4087ee7fe74f519d4b6e9bd101e330a8a512cdcb6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14e310de73e61bd714d24ec3aff45526f5f3bff601e9d9480984d1d9d00c6de703e87b6ed4c167035534f2ef324b58c5df13ac0c46cab20ad957a9b98cb50b42d552cc6a3a5aa063db7556bed1bd4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e1b19e6e327163aefb2166d307a4e8182f5c215005d36293e32fb32c5c2edcb8bc0d7d1bfaec77484aae74cc34e03a351b23c97e1d06ff2c0d3d82991105b2b63543a8874fa6b39c3d8134adc34;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ad99eed12ffcd5135635757dd413029930a70e27dd832808db0baaa49de854de64646b8a06baab39c911563119de81e116b00893ed2175ddcf52aa720fea359dbd48d8f7f56a73fd9925266f69b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h426a87bfe882189b55bce75eb57f1f926ddaea726a374346fbbc84c4c30e432b092c6c910dbcd2c6f092f7e9cf65e676a8c03a7615e9a1714908c3c0f9723e12b2bf9dec670badca89e09e228ee1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9ca76f562f9c331258437119a93489b218154e9dfeff3e580af62ad98d8d30cf118ecba0a6f62c71975bc057d2798fa52da491fbfe188857b1e68e5a02525e35666a7692313b4a538eaa61d461d0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12a9bb4268d2c81cff7d2fe4abb7e356c71087828091db987c4583d5e300065d10227d4eddc17e73076fdafe119aa69043efbdf3767408b74a32b9974df93eeb33bf6ab31f43ee15356540a48ccbe;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h79dcd31a54f623a34c1abbed2f889c0b4ed9957d162c39f0aca39ad57721789a2348d82e8dfe41fb10ee4803d05b0a9166dfdb5ee28614417a4ed18cfce5c86cc2e5a247f3ec230b665238a9abfd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h166a1d0d4b426144303de83b329bbcf63ad66ba16976a41dc9d8d5a8971ea2bb29b4731356bcbd3122ff44b57c33895a5ddd2d34c6519fa0da6f627d9b890b92ae33127411f7a75a0d11fc8ec6977;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4eec32b68b1aafaa66971ce8d3cde731dc8977291930ade295a22d90badaa0829c43747378d441775b0be18b583ebc46e466ffd10e600be1fdcc7df50eb9fba3817ba1cffaee7c84451ad123bc51;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13cf08d4e4d1697404dd0697521682b28147137d4be08986456c1e86c699719652614b5e3860564e7aa69dae6cedbfbe5ef7894e50df1190c9e70d102c7c619617febf9730e6ca8b42aba742fbbb7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf3bcf90c109299ce877ec07b3eed123392e02ba7cf20e3c3d9c38908d24e59ca546ea05adaa8ed96fe2f18339894c1368bfa4a7150b0463604c68e4e13b872af2fa1ce031a44d5950acf766323d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d364cf99ec89b348b6b5473eb2d3af4a5f3532f01b32818464a02ef2fbf78c691511bce219603b61477ccaeebe73f0cf97cfe32c8a616999f2ac23b9e89b7b9109213e8676a9ac4c7e94d3ce9358;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9a58f247dfff24d4da6656dc3085527fad41496dbc8249e857ab7fe32f1fc5368a8e9bd2759c9f8eb56476032816ca7693264fd26124a72ab28fd7d3999604405f6b27991c2538741e6ce56b84cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9f8142a39e4ca4871eec5df690eaf0f0c43869fe52e49887a8b95e8eca0a053a5839dedb4117a4c0d68239a8091d8154ac7ceeb9f113443178136b416609990402f98280702347b5d7cdd4945e42;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h187887b9fe7488b7213b66ce16dcb92794c064160a112a67f4b65e1100b2ba06dfb860fab5245bae3523349ac6b3835ea0f3894c60633ee4c9cbfa00b16d87c1ae031b7f84a16ed99ceb9194391b5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he8d6ae5da04870f45ffee5dcab8b4f74140a9cfd65df829fe46cad19ebb2aced553cbc33d6ed2bfe6824e41345f57bb71d0dca5e9065636f20d822c2205419227cc82374868bf6860aea07a382d3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha23f7af8b905503233cb6043a9e0ad35fc25ba7f65301bad322a1fcd0c994f63686bea70dc83eb6d4abda8af6d58fc3b6f10ce969462d41e540002221321540f76dd9c2e9da2a11039ee437e1d2a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8a73317300f0fdbea82d319c804b35d1bd130cd3d69cbda6c68a95ff34713aa43767bce2bdc9713ad8ea47ac9f2d8c41f35c227a88e5a9f4503eef7db4194e5743fcb40f2411334cc36b0a322168;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6246fa8158fa1143baf0a93ed5aafdf646712af62bf446c65cdff78f1d21f532690c80b922c4d0de642d1a33032203d16c00b4bfb50ab0c1b083d32c5da0147d3118da3f62d22642c376c5d0038e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d9ca436fdbdf040a314fd0906f59f2428e531613b2c209160d98949ba062b577310af81d0166b86b967657f95ac9fbc0b24ea3bddbbca71a6da34f5a1ebf5c5179d4c3a59ce15b95700569999307;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e5f0f9fefaf87744b75e1d95ce8f432352b575be2c158628cd3fa51f4d1228a5c8eea0fc12295fb407e88330ea4a2fa307239d051f4c4a52175e730e51eb4410e74d44e60bb23a156543034c1a5c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d9c438e4c37f755f0a2750cf0b234288fc2a26fad314c3eea1d150bb314d8b9f27d17125f05ce458392991b861c488c97f1a441f0ae9eca8bc8971cc4fb7c2ea6c7abe53667d2fb848c2a9b7bffb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h162ca126f9c03c43282a2dbfb351affbfc767275b922bbde6c03da34920a7d3e9d4230729e4108fbac49b876052139abec302fbc033462b50418f562338409a24208a5700e259d84e0686e2f983c6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b5e52d04af524eae4eb62e08a2b8be40d7c109127e7a49db0827d6881f7d7f015489426698d331041feec9ff1eae4218c55d42a03bb4b08b74040dcff7b064cbe5d8291fd2daffa6ca1beb01f77f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdd772ec0071a8708564a501841443feb4cf6e8507826807d759709bddc64ae0fa4e1a0c423ec520443fb193323dba4bf4f08dcfca54d7ee3fdb488199689485224cf52c59fbb1142e3e4d24d768b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h127e314cc6909c1df7b87af91b03749196dd67bbd8a64a73769da9af3b1d6d334912bb0d980a747e62d28243bcd15b5d6c9d37ae29230a859ef9972fcf9e4645b9a55cfdc5b480e3378c4df019865;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f094885168e8626a4c4f50d312fc00fbaf1f11ee3f7dac241abead769f132a0aa2c5900287f2947074def552e92efc524f978309c96b3fdd540efe1064c322a6e93b408701d3a58716edb107d406;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1016067a0e47d45c936953609f9dbcd2751fab5c062c9a0f9da549ed24226382056a3ab5a0fb3e086d5b293388d5c7d2e8161bf8c9d8933f5c513c16003281811531a359fb89e9ca9f177e4d86800;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h87a6e45e237613944b557242e2db0619a332ea9119c1af78b1a33cbe79671b377780911d6210a6ff0292489ec17558f3d8c5db53774ecc29025f1df20a98a043e5a83a977c61edddd93a355434c7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e0d60b7635b2e7de7291575ba598cc704b372cde0684d846b9f06e8d0b06b4acf3ead7a300565e5ac2634188d972530a17ccf58b7eb11568fbdcf21f4577cd0d6565bfef9363acd1650ce2c05756;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e8501d4cf53305cd2a2349d9a6402f71dd969fed10a7d3bec0c469523e4840070fbc215d8591dd19811bc91504beb7d3c5c047588adfee34b71f7a44a89cf209d9cb1d1e366f685f1b5776dd1a8f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4bceb09149503efc36b1eba46296e4f4bde0d01f4560459fa80c25762454cc890da47f3c9fd4f28d09fc0a5224fbd8f73f83f4bfc203041c46599691fd034aa7001034335d40d29a88e6649f8609;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c3fa23cb803016faa23f0b07f991ab127b492e0047c2ee4b2a6367515cc3f7a172b8c5f5c5c99e6424e03b7bb7d6bf745d10e5a4cc921990ee3ca2565cd900fa524716b1dff51017ff08a23fdf73;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16136e9becd63abb610e8424da6ad5c14051ea62d9253018260ef587d69f6420add580a9ec348466db18e62824a52a9faa95265907dc5040f873d9561c5dcfe83922a4c3f49d90b61a643f3c5dea3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h985be5c49a36f64868c852eabe7893289872330335ee52383be1054c061136604a76e35530c0e303610a73f7905c7e1c3c14728e0f47295b5a1021e1ce7253decf4159e96b61ca0c6bf9b847af4d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha3d03cf8e2b5131e55e3684bf45662d8f42af16210ba18c7b17f86968e84a3c95de5b1197389aebadc48c0112910a72e7f763efc4e9b72d8e1ca715ce0882024d529de3d999e46cabbac27e2a400;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha7a028f263a3284563a9c1eb86beff0d81e4f9a5ece3998debb8d73fef0a6d127fb836eecdded0af0003de3557f3b038065d642f0ef928ac8e7a2eec4799f003a3ba105f17b072ddc48040394954;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1093e562ceed9b80378c6255d5e221665488fe4cdf2e54ff4703debd7a8fccdb811f3ab5564a8e7cc30f61935fd2fb7a1b98ca44cff39c39f5d9bf56d16f249f65962c9edb387875e0d7dfd62c730;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he6e2dcef2e2f7ad57a9d73eccadecd61b5689d7e9a8983110675bce9eabdf17dd70fe28c8c4e4b4d3cfdd60bc59e27f0a6e2d474c34c0bbffeb5da73aaa9890d8a480f7f7748e8e285d023650132;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h6bdbe28c766b1d2e1e4cc048f4ef944ed033535c04177270b4e49da4046ccc152632cfc17cd322a0cdd4f3399e741b4dcad70f545a67d10cdfea669f18ab1ba4baf355e97b54b5d627f68144fb00;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8e78ff9f175cae73d64e85e5b3c970b5f0152a19d024c9a3cb3d8da0f96f52d0928fe0394fe8cd382a22bb63df6470363fe6b4f7ff93789ce69b58041f13b6804f558b69b3f49d577f5725024626;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bd6c67edb4d739b3fe4081697d2d59c4fae4d3c165803dc3a820bb7b87925a72c0010e69e69497b411cea95f25217d1dbec2e8f4ff071dd8cbcdbe6e8079262b2a2d7061ffdf30521a6b3c11b4fb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15302e5c7793aeab73762c83cf77b600d87719289e3b3b9f76a1be0fb8c9cb327e4a2b235d2f793b7fc7c9e55d753f0e84754642bc448b571814468a1b9fe4258a0ff17469b0e82940a8ebbbcdc50;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3c3ae05465e771d6aada4ac4a061424e5c47bf260ccade399884f391356fab017bbb10ad325d069570bc9585c53bec84f04b6ebd9b0b508b0700346e70550ac7ffcb6de88b65d625dc2b86898fa9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h75a266d786b1458334814a572f6cacb08607515471ed85789c86279583d901a71b89ce14ea461043c4595f70734811416cc910bde54442b9ff8d83a34277ed4d3dc571760f855a68c1d341074316;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a3e75c3dfce2a79b516a3363aacc8c232ca93698f6d534133fe3c7e9184b9769f2b62d73593d575c8fd921ceaee52d9eb6e7a8d7f1b79338c7f7026df4dbde88cdfa9cb6c908f51b3a895e537257;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16ec82e4a30498cad77ef2b004820a682495d7676c64ecb3e09574622c106d071b2adc9fa777e7ce8899994924d6e265fa8805c3f31e20c7d191be198267e40675a06cb8bbad95c9e23c9d18e4cf9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h28c5785f284b0587adac0e024d32c9b93446684010a999a9347c0924b7ac6aa791959c9a7892d1266f1622ff784c499aeda6339f22f9e8446514c6cd9c0944468a2c8681fd30064c348baf968fb7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e0ed1d393fb3a460fc86e38348084060370952d5f93e134a532ca7a547375571f496f9d33e61bd6e9979764441566fa44b8dd939b28036b99489dd1fa64e0339960dd08a3ca563753372aa701c6b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19126916ec73f6e1c6ba81d73f692c07cb33f9c8a5dd6b923f61438b214450699a3897286c7e8c98e1bab9e8a3e74d7b6b7f8cc9d13358cace632c1bd85044ecd9183c875d6431f8e0548815b4995;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h407bb0531ae4c00347e163f9a248d5a058785d673179a3218024c704836124259c0c3ad3245f0bd2e90f2cb5368dcbc83a34282610d03315f1a7293eb930240be417c9cd29f97f35fae840b1d8a0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc172e25e4108463105112e1112cede9c8a1ff4ef1be69b86b0c2a212149b4829d29b2f41473e2dca87d282a36167a4b3167331461f8f8838b1bf3c878d2ab938c9db205f54b599f875c9a77c5516;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h75e85972edc7ab24d4fea4c2000ae0fe12b23724fc057e76d865ce54342569af766caea6af653f94480a4fcb07b96a611a7ceef2e7d68d858f2f248b8392f7f152aed5046bce3a84967941032dab;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h57a767fb61b859eff11f865307976b4d6c83158b9103ad8d103664a9ca18ffd4970199078baa25249ed9635f45128cdd58dcf4a9197fc0cfed395c6e077521636479b6649d4e4a2d368adeaf0f08;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd3778a984464bd26f03c00c4041d536ed6bdb8d8ff7143c5651146981da4ea848979aad86c7a4336e9fa752903da84821b3531aa28009f1196473e94a9a4308aae2d950fd467c05ca7ac646a48e7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a88bb255c159e45351aa6c48a7631e19453700826d6d21b34479b78e402756186b3ab9e20f0c696bf3fc43e3cf7d17f3d5501a575f36639cb01f2d3df155fc80cd28a0337bc9ae03de888fe3f56;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5419883d122d941aa9cf1b54688d582f5db2da27f2e665cab03d770c638841f5a038f962c31b4c15df48f7cf857d9a6f58ac0b6bf2c83c116daa0c7ad87e303c1dc3f43a4369230b3986896de7f4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e6014ce528e9554f08857b6c7a4fefcc014b1b0af9931d526c24f5bc64a87e1b060b937d8e53f9d1315f27165b1f11781f4a169c075c294a78bea1983dde6c7f241fbf5e54014a145c35a15d76e5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14f6240e1caaa63e4257494c9dcd2a0946a917bd7ba1949fd4916acd701b69ea77b5b1d788cf45a0785b040ffb3e0f5345a4226fc52b309c856923bf78324a41592668c4600916c3f445fddd9bc8e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h927fb00bd2c6bfcf3dc173ff6ffa2ad9562e1cdacd994681eb1649b951bb8912b705afae7c72a6f62823c5cefd952958c210d1c8140d438c0740ee6ed067dabfd751ce27434fd11d80a6068d7ae0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'heaa377b7da80e65d2c5f177e20cf923b2b4b9a0fa9cd6d90b11c5b892973ff016f590cebd8ca24e19164bb2741d8991bf52d239b4c10038617cf93f112e25293ca7a640ba92cf12f9414cbe76e6a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf5314ee1b4254b997c4090d4abd4fbe8b0cb9b7b5190318535151065341bf32e8d3c9dd30f27d2c00853b3694532562ee12d633594240ffceeb18e193ed891cf8bb1ec30cd9a6019f59836ebaba9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbdc4c5c201e483fa7a06a08150e031070b1a1350c89d983cc06fb12dd17e61fef553de9e74411a6b523d903233978fbbbc58fa0da6a4ca7bc8f417af02e78b7b0a2fa6b7fbe89d36f40c9457c8b4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18885448b3a1849402fff2a4fcfdd944a0422eaccddd94c88ed64b208feba9eae95d18ed6a9e4051c04691010fe07a979dc2b605c8edd8ddcc86d4f96d22412a6b3cf583be468b9af937c0d312033;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd327629b513ee04c6ff0184f2bea110dfdd19df2c2a49721185394f1567b1adc9420884e72eee52ddd04d9f8511a3ab402d21905b3f19831ce787ccb2b2a679e0426af598b575bfbe6656a884e84;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h143a3234860f0a875be5d494f52409bf959ac0c439161794e112058a46255c880cc88a904cae10f5f69e18b1d414499bd500f3e0f2e7819606d89ae91d65f4947093c5dc38e9130dc3546892b7a5c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a6c8b1f58f48b78df056637dd1c4e7eca817cc2036b9f064992fe57714cbe62abd43fb6545dad145583e585ed49bbb9801f5e4e58c88fa483bc24c5c7d59f7e9ba601eca3adec5eee14d753cc78b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbc35ff1d053dadd21c3c4864931c2e67e322e5ed798e0d93d4b7efbe11468de3967cba79de8e634e5780d4624efa86974a9f4864e011253a0a4fec87de3d0ee60c23060577e80bf46934a2d699ba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h97df4f452f4cd108f7131d0acd1a3db9245751cd4210a16c8c9df505109edaa355bed73eb7fd3402957c1e0f0fa148d4c7cce439c8ad91054f1b55d236bb62aa0499ba13e6571e2db5589189dda;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf21c718aac783a5d6f59fb840f6ce0fafb421e61285fe26c7168d5897adc19efac1b4504e957b5d0c3f75ad125a881f91783fef68f9bf2f5fe3ecb69bf8c76434b2e5aaafc506163828a6d755aa4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h729ea57a8f2249da448886a33b7a120e9158036d616dd10904a77c678e34b5ab564e69a7147de3b0bc3f4499bedfcceaf91df76cf20f4897ac2106384d3260930d132b905a8a09aa883b3f1f672d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2c23d2f1dc4a72ac6b6f15fc09dadbd0f489fbde8ebb9cdbc9fac52023bd71dfd7cd568aed566b87c8431e665907e0e1a8e0c7850546e46b8ac299d97cd0e565bdcfaedbe8897aa3c0cfc7759d40;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h117dcdefc09158e1a4f20f81cf62887cc4cfffe54dba289239d8fbbe2f348b7bb9b69682b155482aa3f50fc318a866670472eefe79c37821863f6585c9da8ec8ff16c6b98dab091abbacc8f5844ea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17f660435e6c9634c579f1efe2d512d523a280832d872f1cb4f9f7979d568360edbfa72b89ae4f17230aae4ec9d1ca45338b13f3ce9ea2d4eee43c02f23be265572cddcb986085109db50e46efbf5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hff0de9e5d05d1358df1d38777a22edda539e65b448fd7679938ba93572e410a5c2b14d91d62d0a83079072eedbe0967f299621b8b077ecca9cea88f61e2d723bcb1b8e3a1f24e3015cdd6bca4d8c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h117fee032cd691fba936fddd7092dd230f33a555fcd030f9ddc4d4773b6108bda251aad940878e11bff4377c5c432135a9898be60e8c01fa43f71a499b77629aab4011dbbac6e2d311b7528365ab3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d32c798266aff5dc700d6bc90254ace48a01725e7abcf600b6e5c6c85698a125b73d69614b538a2f385768a0d26e153526611901f6b34c667294473d91ee4a8989a602f8e11a87efc05e16d81c95;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h126fccc46d739b7af2e350c1e8fb15100f17b52599405c8f209b4ac4b192b5b6fc005b782362ef5f2f377ad6ff2f7860956449ecbf09884d552d7f48da7b364dd32ee94762f03c10f0bf5bc310a6f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcbfb5729549bd604acc9f59663ecf7cb299631904a059f3c30b351c8b06d8e8726589c26c9d1bebc0148a0b958bb7322f815a9d0acf6e5718c6b3dacb67f5b7d340e7edfb15d0194ec9397426ccf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1be7ec0797d8104d11871d71c942c8e0fa9306b40b6bb5affba82f2da4a693cd3691191f02c5c83c476fad242ff9e62bcc50ad719907b0d4f5191aa94708456be4a0fb1827adf39a0e2cd63e008;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15b5b051301445142287f1408df8981507ffe494b6eb8a79480e816fc51e422a1916813506766f124a54c5ffb5539e53d671bf1177a37a4f06bc7ba1ddb893508da544af0c996f50e9e3929f3e693;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h388ae331ba6400220dae794b8bf457448eeab48e21dfd36d476d79a84b742864c50cdb243ca3dd2fa868e65ffd5d7e82cb6e17717678d7093f55e17858de25254440b8984df0532c973e507fb462;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb3e9ad1ab4e3d0e111c9687ad25f9ff4365da7ee2c775c6d303481cc0e4516e32413bdafaaff54baddbf0e892fe8b3483729d528076d3d36534584fa11bb1f9239dea20974606ca8e37033495660;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h84dedc6a7ff15a5a4ac48f843819107e66becc23d18f11a22f02180fc0cdeb6e981091d396010dd91b1d45c73988dfe31ee93cc07868580729e9601aae20971ab106185c34704b419b57e5c6645;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f6d8d6ace1cba0442eb3d89bb9aee2bbbb5c4261df1d1f8141b36bbae0da0d1cfa92a87cd9a1a3101523e529e9a6dee3f4b989813d925404ca42b89fb156b030f39b4c0eca259d5c038c517283ce;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h547c87f651cabd0b8ad33e64eea517508d4c3d609c3cf175d6ed67422caa50efe8f2ee4eff7256f54a4de7bbae5cf520428c6cab1b47555b3a6686f4fc4481c60965d057a6a866483eeef6d48fa0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19c1fdba7e7d1a1f7ff4c678a07f3a8d54f29a153dd411bba2209fc95631bcbad0c9ef824ea9ac5be951a0753896a95448e727ad5c7eb498223d79c216a4f4a6544e72a0b106ffa621eff8cdb4b5c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8b0213957e2e4731986fd3090075d3eeaccb028a6754f521097d07429ed21cec90fc5cdda5c37dec57cfeecfde1ce0eccf6f6bbf874bc07fd93acaa375be1edefddfeb2e7d2ba69c75bf6d551fd7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12be3f540068872b5dd29a9fb311248a31b3d089caf600c81852aacffb070ea481cb79502826c8d97555fa14aec39f33dbca76dfb8f8b835f6f65293288c3155026e0e030b936b2ae850e439db85b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1609e272d2e10ca5e0f5c7679c53be59b0c32d974336f2eebaa5069e062c3034c610b948053935ecc67ebb0a433199129983ea752cdd2d162036f417b4a561a13ced8908969bcf2637ac5f69d0eb9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc2541b6cf17b09cbcd34d585ade6b3f00a1e116ee88b692d0b50d722bc11cb9ddf4aaef6a55560d7e6611a7f8237d0ea6149efef6fedfa835745b9fae73438c55e15779dd688434f550c2a20aa38;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5f7a814eac9c7c80d83186e67d06601d0f87bd6c425e008a8a9fce8254fb376107339dd7f1876a393a3adcc6c2b52bb995a6a518acd46f9fc3dd80c7dd479bd1520817c1b91b461ee7a6acb41c0f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h87fc21d0eefa7b993fd2e523a2481bca2c8fff6c5d5cd8c4c40de281050cae951fa7e659fab787bdf7b301f638e24521bb1ed6286841ab2e528adbaf77c45f2c0092f00cacfed486fd8ae8942f36;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbc6575b37d32ed5d52422e0c2b07d4db869248da4ce22066df80b6fdb9f7b35313516f5c5f4d7080fedbfe6b21644dfb7701b2e1feac6de6e5e75a4bda8194579e99e5dfaf7675995a0dd8e3cd15;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h143e8ccbbb1d829c89ba7ed84f0001c0d457ade35bd0ecbc25d841e6c424d7ae0c62514bb47b174c3d0e9d30d8c584390776c4bbb28783e5a444cfa087d90d96945d7614333df6193b482763e5268;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h402675903d61ad2f99228159ea9cb9f2f3da3cd198909b50a92259a7fb0cebec392ce306724ed08d1d0f8233e2ad3830c079824030edecf459e0723653817332773da91c9d593ff840d04d77af6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb383a9862b69e1ce2d0608ab8825ae0d2e284f2fa2e3f687ab24c43eb379bae2275cabd9b397cad39ab045f5ac6d42deefe2a71ee6d6b28880c92031ff8bb9eb0272d2784bccf73f23b171c07bd8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4591fde9ef7995d1c83fac18fea3e7f3f6fa76b6602489df0651d762faf7280750adf653c53f63e3a0fb027a13d343d677c3a4822eb61cd1913dcb48c116b7213a2acb3bc04d1ec151eed2f6a404;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h53a6fb993f389b8d7c996c1bd8e2615f91d9c9d30755afd58bad48b5fe404a2de52d274ce25762ff72d8932aa35ff6d79fcc5f87dc2f7f7f7533d84d2666aa728942c4b77991fbabf97fabdb632a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h336bcb83f800917dfdc3872e98425648ef4aca77489af5d44872109bb47c117082ee603461a3e348426cadbce4034b4cfbe7122dd13e50c223bcca0509304aa9624b4f6232dbb0e616009e03c60d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb1eea2e6a053090ea251d59545b4eb562a56612ad106e79afc40488f19da2e67418a07490e5094db190e3207089e954048f210f8cedf16605ee7f13aea9beeaa03b3c6202ab52ffb2f5f2bb4949a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19a0d55560fe12b646940adf1f16cb63131c0de7e9fc34bf9f1124a9758bf3a6993005ef5fbbc8877774ce8ca24f7817a56ecf06960a177469750cb479d213e7f71d16ff1aa11a4725d3f8ed0b17a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7fc5562d1738cb072a2c192d500fe01dfee2006ce2ae244df4de5143e1bfc83ee5aa239262840205d996a434253264dfc758f27cd8c9aee5267a80c6b29052ca2e088c18d6f280daaacf2c2290a4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h152cbda7d9079a491be048d45c41539b7f105c1d53f7c1f10925dfdb2faaf5c4b178632ad042f2ddf3cdc249d12a072f590e82f0507d64a5d02aa8f1f421296f1edd1b524258b527bf3de731eab95;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1419d01cad4c61c2614c7fb4e970d68ea4b54a720f55aba46f12fffc43e2150e1fdaecb8baeda1ec1a621ae7af99eb46cbb940bb86fadaf64236c70e2844f174c85aadb2908943d1247968a4b3233;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a1b29193d2b2e6e6cbca3808d5d66b9429d94e47793bfc46d92aeb37f81f268f7cf08c32bfd984f679790d6531f5dc79927bf0c18a87a6c747dc1942b8430877427d654accca5b23a62085577fc1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h64aeeefde2f52de9fc776d6f2060e85a71e189312fdfaaa261ca0b67681d57bd891c78f7bf6536aba169f46252f6985541e29a19ae9b4a14eac6f7352922248b8d261b88379e81cab23ca14c3b8f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2a4435ef6c99e1e7a0da78861b1dd98ff799e70a3ebf728e7c7fe6b488f8389532a4ae1345e4489d73d84f9e0fbd99b38c3e8fe6c9a3bf3af68131fbbf4b00b04fbed4bab99acd9c228948c1d66b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10520cad0214f90b6a9613de3e21f84c52893b1093ada97179f9bd0ae6d57ca33226a11f9d4fd44fd896b9cfcffbbf3e17768c2c66fb98413041aaeba50773dd4051098c366e943c2364b1b6e5ba1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14fd5b50c06fa4b09a2d4fd2750b18fbaa8e266c9c0819ef2fae72f5255c14229a8f341d1a80f8bcc1e757346845ca72d4d5de6b3ab3ef258cf695caaed66475aa061871d41e2058e50f19edcce1a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1370670d34ad271c82dbe5a6170599d9014319400ea4c8a58cb32b6d600f469e9941dddd46cd2fca90d9edcf4cb86df059e1e2e130ff79bf1bb036e29ae0ffbc8bef204d21705f9ab6b16947d9cfd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fe8aa704d646ba60baeeb226f95d9d92a6a4f99daa77e7592efe8a9b382a7b468299934f7b6cf4dad07a83a99a0492b1abf4d849c41e647543e8ce1ce2f74f0d51357dfb9989397a434927d0356c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b740611bf4846b6771d5c70d34e72578808cc7d446c08ae3683ee6f1b4831bec6af677645f52569031fd957f88c1898bde5516c5f39df863cd2201a483805a01f1950c61641e6b68d7eae2fd73d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19e3bd52a69906791850aff8e5d702d7ec14ca3a366bb7939a76f63ea22a7a0e718766dd1f5c4deb9e140c6cfa865eae680f75017918f939aa6cca36c53042d5c2c8debaadd7eca8fae2856884db8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10d7d98c012f82188812025fc43648d172948d2e955803f6024108d3901dfc5b44c4b99d617dc6d8f8354cd8f1ce6623dfb4a86eca8523aaab261581eb4afb2162623a60c39092edb4d72fb0fbae7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10828fe507aae81dae4b94a86e3c1a558c2cf6a6513400ce1d057a401e7de55f83e56447b6703f331086955360e462fb628f535a2d7900b5077d48ae981a2a02923facca85ef38553d2b182ac4d4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h878e0ba55b6d23897689150710e370c00eb309142fec71814006ee80d3d04e820d4c1f4ad4c8f0ed8b169d0f0068441341ef6b4f71b5d6e98d1608518e8bee4e1f3b11afd7737f9df37372617500;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1293caf5570cb16874ce265feb0b163091f44c4f230538f2aea6e4bb58cdfde3b7b2480f28ac967b388b9a66f23d28dc9db0388b01a18fd750d0f574ff48e64ea60f977e433df956c651496b4124;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1f4857fe0a1ae80bab8d106f973329e20a01423d9c6068f74594de48d63e3e23509d3e6bf85937323931a20e3eb6d2bfceec2ddd903f66f0f4505a1db3dfe0bfccdf3135249d718a44a0e5cc537;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h109cbd5d038f639117118bff17812a96611feef8fe8c5f28bc4340c4f77aa7fea2037cedede77a0b807b859cf3d28d327ebc087f77a63d18608bebbaca17510e03226b451684fe7cf4e6c3289ff4a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1030e2f49ef65e34b41d940ddab0094f7929c68bd9baef8a4430875f7c8004d21d955670573907f234affbf377b0d820e9ad6525f8eb66601e00999c5dc5995a95e37b70c69306985a04468a5ee60;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cfaf2d0b617fddf77ab8c02624384dd6a0b2d14ff0667925b692db7d66fd5accba0b746089f56f13c61e2fb705fffcfeb0d97d4fde09a2e6ca9c429afdb64eb613e7ff2fb0f4bc82e89d10270bdc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19b726b833d1923d1e799a0616315d619deaf61695c761427ae853837d41bd61c218b72d53ffea703a85ca2005b2f4425975dc08094ad5e533443502402e0445cbb48d7120ba3c9af017fbc4812fc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5da3ddc4dcd95892707939706c777e9ba8a416c88990ba6a278deee3eb361d36f63469034dda6dd3a432b46ffa0d716423d09a29306f8097b566d4b4d74dcf814157a20bec817f06387286777dce;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18dfb6e56b597e52ac57f9e2cdd469d9b34ba4682c0354a551bd0bbd22e0abeaa44958c614086965cb0656782fde0ff44fc9cd818bb48ee6df2ef67510997df0f066c6cea7fffa3d0c5305dba7d29;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ab7d505a288a9fb0389b2d810861d25a38eba971c5f990776673b3ae9ec4eeab30a8731ee9a47a8d1a9d666617f1be5f6baaf00b632f424f6f8fc58b14ad8464d3b46cc545662d0f59128862e4ab;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f9faa4b70fe3296b619db32350f56007440625e3fa2524f69032d8e5c469306290695777b5e59d9419a5f0410eaa9cd0149d8a1517fd5e3f12666561837be65e888d94a38354726a4b237d76f709;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1365ef47e6a91ad3fe2c85eac6e2ca915584ac3299432684f9788be015aee2bdb233313b36114037af65a8eada4a6c8efdb0a89d16761fd386370b6952f8749437a58e9631b927a2352f141583;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd94a1dd40f8b4cdfae8e2e0e66f4350f96595ce83a8627934d63d0d637cb2469e7c15cb1b7c4115b97ddcb826eb15e27b4418b33abe056a00c93ea8fd1ca78fb6e1b06191a7208ce995f13378e1b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h95045d02b005aa7e35c7ba76e51666c2269779d000511f5250ef42a2bb68c80e93314031bdf13733db879564d2383fe817e388fb7a89f5d4117d51c9861d57967f9ec267138e4698984813a92893;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bb24a792e71581c544ed97c8605ede011893c6e2522265e63de166405929a7085a5ab9f6051ef7ab4f7e667e27a71f403a4b7210f264dd565ac60f397de322d77df39c43eeddb6b84e6dbab0f569;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1612e1419f96e9240f20e7586cd0f589800951c4834d5a1632434299d0719942863b827420758adab20cab76fabfe549f055019f36dcb4acac8ca958b6521d20568f29bf8bf95e7cdc3971dd73bf5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13a7833d93b65ef5c53567847ce2aaa2ab49411ee4621241d6720621c2b577d343b2ac5c5f9b89aac8866b135935f7459a1a69b2bbfccfd73522d002e8fe995df7c39b1746c4d45aa9230e93661fa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15415348627e1de8d001ef0923b4d7cbcdd94e32a8cd789c05607550ff5f83b2e74df5439b83c456112edf8b470b01a3fe5318dacd3fe22001eb6d31a9d8ca6294179fe4f4cb5e66a38b04422ac56;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15a957a1bdc785177a21e02c19bed415622414184994f96fd6de90cdc71aa20c1ed7c42c761af28d08edf8d49bc465098d5dd8163f47c56fe0d2336484248971334d50a836b8e345d0c43f0bbf823;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd44e803a8f1ca1eb3c8164287da92a971480fcf76e68c550098b76918af61c846e513a7d13da429ff480900fe3f0888d0ca27072336a7d5228a329ce81375e594433252469b027d2440253d72fa4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfee4247af885e5a8d792e1b6cd7d16983adf0d273013055fbeea632f45dddb95c51aed349d986c847fd2d6846fe1e7e0fda2c3ba5a87a81492c7ccd796c7db899747c55a42cb153184bc104e95bd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h163276035dbdf1a45fe38b23361b50950b9c0aec4f048770498a6eae70e074cc65efa66de04fe7893a4de9ea608d850f48973bb08033e6523e1a4485d6fc55caea95ea3850064847d8f128b2b37a4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h85fd2c3b9b5a5aa33fd79def2eb6dcbe6b60395009840f2389392ddd419a07f067c611bdf5d94197eaeda65fbdfa3ba0f7de7f8fd1060e3790e92a1fa3d3848ca57f3a11591dc6bc2276b84ee9bc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2f0b82014a0f3593f094b3c750145e90b0d1e9885ca848e3cf498a0e157f451ceb404ac4877d6985b5f3a3eaf31a6de6efece659b119ff72db22e893bf4c8c964566e2aea29cbf2f75d16d471d5d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hab57a639ddd711a0a765fa1964512529ae8345bdd40f6f16c459be013e219320687f76387b5ba01bd96efb90214e3e448e7d4d00892c0b5a1c9da760fa1e8b3794a6f5e23306c6081ee768a796ee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d3adcbe1b1f5908e481db828fd5404cf8e0083f537866231fe6111a6b6855e6ccbbf9fac0b7bbc0871ec07119c2c0c36859b85f59c0a653c60d9b06687dc36ebd440063ea7704bdb1ae086599309;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16b6d484f583afdf65d4a42a468b1b4815a3de24d846e7b161c4c24149a16ead5a17182ccd10c95a3a5a1edd5beb8ec2f92ee1f4d8b9f9f6b47b0923e5c8e9bf2b8cf882fc239063770e18de88306;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ea5001d68fcd782d3e080857572a044abc2a993d42d15b481e926f71e12b43adcba18618180a7823b0fd9ba905c49dab024064a32833b14d8b81bb2fc0c3e9edbde5830d97ec23991d4e9897715;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha0cea371ac8c23d3c4bdef462a3e4fb7009d9bcf8269e2677ba8e464e6d3f32d645218e84e151bf31b8645d86decc2b5215a867aba40797669ed03fd40bb5a2b53cbebc411fe998d203fea4e1224;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1375188ae6d0821ad394fa7cf9e980ac1d89ced1100d72ef14679d4ad626a2feb2e02c0fd0ff4ee72943c3825f8aba49ec25a6dc571f76bcf4f156662bb0df1e9e6ed172373cd7f5d48f77b95dccb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h477d6a0e55d65b1c3f522e3a3a648dd60264470ce8e620982e0c0c35eb37da8ffff08efd1f7d99ebd8af91cc8b54ff0045db5ffa750e6080b6ae2874793495e4eeb28dad5538399bc420e5192fc0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e58851875fe5c4cd30f390171584f5a0464d4eb5db88cb388aa8fbe316201f2d2cc265a981c8546d7f0af0e77a69d156f47ec1f672e52176dbd11e511499753aed3802418d3d9913ba58884a6bb8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9b464965c95813d8fcba329fd5340ad18324b94f26bd9522382065718d8bca8ce1ffca9b4ccd87adcba0b92698a3f843ff93710a456ead9c7d644c8c0fe6a29738108ac9598422d3145c0c9625e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf5d569280757c395a83af8b03f68b3e4ee3ab902152f6e0adfff633e50da9b308ec29dbc89a564f8c4e57061a673e237a8ac09d357fe0bc9817ed7f6343e85eb652a5221395d350682bdf0f0ea3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h80376fdf514b9cb28ddb05bfc4c4451f5ef71cc5b7725cd8e9de6d30b6f6debb4ebc832bbb4a7c2c9f831c19386195099ba847ef94d40366b211bbee1b30a96a701997664efde18315747b09825e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha584691bccf2386145323d6bfdfe5a1105954b3b820140f632df8bc1513a65ea99250dd42cec04665c3197297f3eea2678ecc309cceb5e00550ed02ac8187d6889ff815bfddd73254c7bfd3a6346;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aab5612c024c45f2976bedfc2998b7e60bd30220b7272e4aa62c19f406d29d9d179ebf4021948a7b5f8be44a61388dfdc9c2b99620a836a4b426c1ebc9f474ec74f692f6bdb25bb432e2a916e510;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14fcf5bd39d2d30bd32c7d3ef8a635b4bf838cab1a53c442a739c83def1c974a2bf454636d5d98314627a06c8d7d0f79c73446046f317277f9f5df0ad1b57cbb3e2913dc9c5f2b2de5f89974a5257;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f80f2c13d0006fc6c4d0035e5f4ef18f7baf3adc9a45dfe4490059d091c07c6c4abbdf41f60a44d3f96d8eed7f8b2fb23593f005e39273ca9a4db08daca539cd464d70d0a62971f8a90d082c9ba4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha319ddc7c31c41edf8e632bc94c52787de62513d223dec1660fc074fc7b53f24d79693f56291024a24eeee397066915b09d329000b358fb7eccbd0197dfc076d4fd2983f019aec34b03f182e6368;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14bf7220e4a7eaff169d497318d38041d7cac8ce75349cf7a9501f95f005407b30ec3ab6a519e3c93e713e0380ce1ff37fcfb48cc99b599172856e0d9651cf345b2b312c1a3a22ab9762859210208;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ab0a9ae01e243d64ce08c970f9070f5b610db894efe77b31c91acb8ca0467fac4de70a032676716b285ace721d2a5bd2d7be4dfc771f3b04d9c511c5c95269c811092c97df3ca2e2d3dd16239a6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h158d258b27b093192e60199d2a95a332aa4c93a1596ff5c291ffcccdc288aa456bec8ecb581b96e127ba75547ee53f87e66f20862bb69ca397ced2fb51fca238bb622c7ea49e251a365358912d108;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h454b27bd557f127d310ea4465afaf1d386ed932e36db937d13cff4d38bfbd6eddb53870f1e042f3047234ba1175ce7b7042fdf41743a754c165c7517334a51d7c82ae422cb8a3a6598c2363ce7a9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hafad0769734f3702557e110785cdd5f8f21934e7da7884434469d03756e11b9275c0516916e247ebadf8557945b66a9c9a7b1747faf6cd795a16cbbb96d580c59052df720fd5bf5184a4dfef496a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c41d5d4b942515e0b312c6da5c0ce2eb6fddff3f7e76d5ff9d050fd775a4a4c33b11b9471aa020f3600f6002572a48198647083b1ef1bf4893caf19e59126a42236481684816f6d4d08ef38f6d01;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18a69777b103956cea51256fdfc1bddd6b6b1d56c659b1fa0de033c881239d60cb3fd5d5a8c648b4ae861af23f722a85e2b1f5701c2ae9a355c876b0553cebc9e69253fab8604d83be2903040ea0b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h269d22a1319ec1d1127bcd556fb7c126340b15f4ef9565cb2811918cbf8a7ed151fe037c809682d7387ec420fdcdd649b92ff95e2e54cd813e960dd07785b8826e43cc8ca835a086b810782f5410;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aa846f9281c4deaa1dbff2346bf7ae5203f4b61e802c66d221f6aa26cbacfb15fbd0b619e814d97bc9a45676f5014e0ea871619c89ba37b73a68c83bf98145b8e1cad6fb7cb7fff664cfd5dc00de;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h171511750cb11874bfdf0a086b0addaf796c9bb19b839ff2e977738a965feaf643c9086d1ed5f74fd66a2737b040c32768774a37806ece2f0bb31ae148994a35c9d260d2cf4f19aa666533c43bcc3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15e69f3634eb6abb5e4c998cb044ecd03da68708dbe470e2d46c55ff04e7ea5697f1de1ed68328f54410c3e0845cafa5f608e4d1368c0ac6577cf09d4369e9130548760b549de0f7ba7eb19718282;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4fa5b834e85690c840addc24bb09d09a7141c6f04de2510cb93fea3b3a305bd4e7e4e73f8d2a21a432a54747d549cec8609afd76dd82af1676b7454b8ad2b41bba5779ec4295b01be573d2b4f614;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h48dc09e5c94b1917f7dc2993d6ffcd1412bf1594e3c534d3a97f080b138417c3da926368f0d22b2e137dd56e5e0afd4446b019ace61f9e08c3d372060d313ec742aa4865a0b4bc8c5e5a5f4e9072;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fe86d4c8eca73a88d05eb390b96f437fd4d36c9c14f225db316672d591bb5eeb913e3abd434036d33961042889bedaeacd67a3ec4eae2f8569cfc1b6fcf61c1842966c4a1df5bc89919a58b8c379;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h50b42215b244293caa3eb88429da7e1a0b75c81169628af252eb329c0878bf4b0d53e37b8c419fe976804947e1bd1114bb1718bf6beda029f6c688665f6d2d0d3c048229ff990fd4b9c94f22ddbf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b608a2f09ad9b04ef1bb9727daa43e64bf03cfc96210661b470b5257c203b86f5bc22b8c29c73750e44544551212f15a29da3e0329157afd166fdbe401dc9a1ae86dfd0e412221ffd874fb4240b1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h115fef68a48b99e95069d17b3f4d3e4ea19fadf55879bb93d3969ebcbbfff2ea13cf45b5eca075c1fb7fe452e16b7cf4f5118e7d59050c9d05f89743e57313c47fceecdf45da60563df26d178d8b5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h411ee3ac3e85697bff5ee3032bb79259502979a77db59457de0bbd7c21f0597c3d7cffe69c83dcad5cf38beee28ca8161b63f89f05e459df74f9952ede61bb71e0a607965eba1b751d217133fc4e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hade20ec0ee71a726507abf9eb1ffa4a8685cb29eb96fab4cc0fab8d9d5d8f07b39040c87a02db8c7120feff7959538c998460325fabbc65913a9b79955c79cda40a55e7c6db200646cf1e856959f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15724055755a26396b996cbc2ce98c24f374f1c1b5d8b067434b90ca52c977dfa69b94eb379154e2f539ab903caf4296d45bfc613b4400a31da3ea6defa969240f7a30c2bfb4ff85da89c6912352b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c902fde6a2af420709a54d2bf5af6a079b27409feb02d0605c4d1fdd4ce95fcd0f524dd8e1576086a3e190b9de4e9b60346de9f72c3172d10a024581b886a94e5f7d9febacdb38c4bd9f44d4bfd9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbdfb18138f404a7894f0b4d50efb68c4093816e45ae7382be0fa313cfa62bc904e60b3145982a97c241f48858034a19d8e47d61621888348a54b3fdbcd6fe6a4f6856b14e06ab1abac76517bbba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7be252c95b5cd4969a70924ed0768fe142ea27afccd582b09edd0710346fe8eb900aee118b2442fcc433c97ed7915b85040ff4970fc570c2e73325736e514d8fa5e6cce28e139e07566b38c47ace;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h111be52415136e8dba126747337716fc0a71d14129bcd4633947b29a1640da1d12550c2217122bd954404ced71452513bf2245145845dc0c66ea28f1c5de877fa4fb66724ffa4f622f9b1bcc368ad;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf24ee59125ea6e8601a81a0c87dd8acdfe64ef3f5ceac503e63928dbeed32461f22f54be7078a838c0a046f5e857eee049b3da88bcba6c0405f5f0ff1bd0ece12b933103368c81d13bcad79f4b5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e0a76ea47443610568c89ec93513115fc4063b45a93fcb2db3d4836dbd3fbf6f559d4f5b8ec6123af202a1155f08867c72fd59dc56d26fc55b5c176d568bf64c3af59434dc21093d2b2cefe25d01;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b643a2d40b7b5a9deb63dde5cec5228b3682e713d40d90c0784552b28ab543585538789b7d9f8f9e8c0bbcc06422eb0f4653ae85c1b25d8cff8a61e6830314a0a873f48881fc12e67c9670e202e8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h25988bd6648da7cdab577ab9f0ccc4a2959776a85fbeed6b42da9af0f1bcfc8be3315cef96b59008c8af383233808db74c6f7241b5128040b630d48b108f66b106375da072348810e61e8b54746c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1db359d4d82d6c3fc23ed7e6494aa476ce4822d19a46ca50369bf5603af009eeb8bfcd4c4641b038b1a0d72e9f5dc3a367748d57683ca9daf8c6a14f6bef2ec32dd9c30d7e14a7e78e81bc0274201;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdf2543048713b34baccb1a8912b574307e5965cca4657d11c356850ff864ed08a655fecb47edd4406fc39f99e3e71bb3c9e03f2f23e93e444d473ccc5ce632cff4e78e2813f8a2eb7800ebb69815;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfc2857c990b2362b930f2c2bc6d34c90b32d1e847a99d36c48937b44361a4b0dc6359ac189b7c46aa1b3a298b8afdd286f0516bdb7b8a18058fae4027e4496c060a53a87031030ed614d4f16da2e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d93ca7303c2acbba2b66c6e586b6c9ac75ef6292d1d214076bff8edc8d2f6832372608f2a7cef6817fe9e1e9551d62a00adf6276ebb7885a19b49da939a419268f51c04d194af2e9c65c28893e16;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he3f0c4c69138020b15dec5a009e6568bc8216473f20e5a85ee734691aa647172098893b3ea2409452862370d6f025ac7ed7b6d716db6220c53d4eaa6f73a420b5201a3b44609c4dabe0d3e68aadf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he905c5a91f7d6791bc808760c69ac7b2848049420d722c9d0e20673fcf70a4df5d7c6373266eb40075dafb6acf70b11e923c58cf08abe269bb21c94200196e4758f490deab8662ef8e0dd02e1cce;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hed7f89ee87828b626a04e5b56d8d363025c27ced961128c6399883bc444b76081236c668942ffa9cd7a6d5966b0dda7824f0a130a178a4f9d2df0139baaae4a399644ee495279eb99fa82d5eea1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd26fb28733f6e5892a1b29d7171e5654ca9c4f98433896a26eaab06c28ede026f1ead4195778f2562195fcc2098caa005a02c93ffb41c254992cc152a601307daad4b202c1d4d2c4f9932d335542;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13a838c798441910fd315ec7f7a71de273ca5afcee03540ac47483a3e781105ab3e340206e13261488d485f09b4e167be16ddbe1336c118e282dbe66addd483b773adcdbc582664d556a293f96aed;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17960a43268c03c5dbb58aa1aefe301d45b387e9ecd30cafdd1b7d0ee4b667fd3f5e86c33ca5d0f0ce9482310d7da82900c3f579d9349b241affb013e1b6495cfee2f9f89b4e7b84e8e465aa061fd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb0fc00219286271e694a34eba77505f5feadad4f3f1acdf8608a9031fb8a4267dfc9541a82b39dbe42b3a6ef0af9ed42c3e4926f4c64edb27e941dbe629548301b6f10ee732800e8d8748a600079;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h114741bed61a24826e1d264c4c55c087a907f45fa3577ae3d15cbd5f3ea75ed10230e20536eb8e379d52fe0988ba29ce87e3ee459b8cc9cb6a0c16fd4accd044107ad68d3d34760cfccdfe40cced8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc1e131c1609e1ad2c31f9ef21498000a321bb85c5c27c3b39ae8dd7e0bbbefb910b6c6aa8a8608bec6f935ff09d9a7a30544038c7c7b093fff9c5323ccd2c6c16081ec7874c523fcabe16421ed78;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b618510057179e394d89893c47c8bc88ae7c03e56cee7180e70a1a7e9d29e21c0ac9320ffb6eaf2a3dd49b43716d819f4fb630e337f38f59af3b440e90a3baa92f0b414fff16e0cb2f0522a358e1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8f7f6ad61387b534c26e0cfe1dddf6572358102fd7cd78410bd55bcaaca8379241b370b5745454991e805f86d95339d415d38ef7a31cc4b6cd0787eeb9a102667963718b9a7cbeb0425051cb2fd5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd8addb3e02336e016a6838ec20c641443ba64868383ccc14012574e1d4648a297dc6789a492d5727e26906db8a1271a515d9af63281bf6e4dea062e8fe08eed5d24f2d8ed51b0aff4415e8c6dc70;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10c6db3bc81fe2f83194f805aa5ac698b03ac5cbbf1dbbe86879017d95e09e0091b1418453c51d2dca5096dc79b07254da5e5d41ae281a07f88cdb8116053585ccf992c6625dfa10dac844529b736;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he1ce55a473dfc3bcba67a7b64bdb9a35213b70c05470bb31f80abfdaba7480bd242e74b70e87ca00f10044f0e5661f4969fab54a245f3ba629b2f0fc07e5f13560bc27dfd85993ac96fe0f93dea7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1692915bf2cabec886e4a4bbc3206e000ee0524035b05a781dacb777f55506a589c033443137aaf15acec6d07c90c540be7acc3a4343c28b22bf6f990ac3c10eb4e7df42570ec3ef0c39f3ad88940;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h32d1f147c6953d7bbd591d1fec8fb65ed28c31dcd1f5953c63281d16ba1718811c372cce031d2519a18d91fe88eb0491240da0755b1b76fdc4779fac79770cb7e26d306c0e239b42d6c7ff45b6de;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf99759df8a30ed8e5c967929956360ab3dd19b2a7bc521f3674e743914051aaea49fc099a0e72d0db9cba5af4d3b368ed47690f2b1782f13eb6b5a71bc6af6b798504c8ebdbd276dfaf14320cd36;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h125c50cee051d13114fbed4f0c32e24c549d55549b15b1acd4b1bf2aa586c789d6247997cf368c6c84aee994c39a465ff05d6eba55a84b6eeada46e49442f316b41c435b42643f881d67eff2476e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h141eddba906fb728d561ade4f79a90ec8d01b455f3005c0a6625ab861b3761def5bce9c5071b8b837ea08466a26c13bc7de95907ae43b50bdb71eaf99a41a444bbb74828e6aee3ba46fe4eda0a51f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12ca4e93017ab6cb6a74298cac2466c84f47ffa662f2c9509993e86e1c75b45d7e9a9d623948d765d7190bc26e0cb818fda811bd136af74c29210bbe8a4d457746eb281768526b637f30e6cfd68d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h26e6e3b586ae309c5344f91282d91315133a00b724b81b8d720374e132620fac2a0b3607c263cbafb68545c3c47332dcbeea7e20b6cde4d6551971e6ad1643077771b1425f3b3e92df8089c146b3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13b1e16369f47ceb562559845f58e61f097744f78406e25aa5b5c3087b86deaa77d78866e84678031f51fec84dce4c359f6898a8cb6c2869db69e3a9752a890222e83546cba872e18a630af84cef3;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb02e391bac3516e720f39a43f88572be91a767ba86d613f9d702a02ffcab942fc1789a6e7e58e95a6c06e8d878f06fd482b753cfc6c0b46e04f406b0ff882ea88f9bd2f7f61398cb722bc8f02673;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h129c215840775d267d85122ee98446939a356b0424fdc0afac4010058318031b197f893f20a89184ee5e1da46dc293b040b8289d712361259143ee9d168bbe696d87017bb8237d486a17c410cdeed;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd038e56898297888e7c19157feb9983ec227119fec78d6e85a8998c33701696141959bc2d50fec0c5b9f1ae3f6c9c70ce4ac2edbdbc99bfc157ac84939a3254894ca9f085ea4288916fe5d987413;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13124d63fdfc48dfe430cf35a91db1acc97a9d20115349cab8def29b6123389ede8d3c0beb7348da17568214292822f362ca8ba343d9dc74defa59b186d278612bbfdc5f281d268a9dfee56d4640;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h69121e62ab46a1bad9808128890e13ac7faad00069dbb00d5998bc052b14c761978f6d67d27c2105d03c720ba32af1b6f9c81510559de9c7f4ebed0aca88f475b7351f9c934c0fe01de203a647d6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h43fb1017d0b9488d094d0b97aa98a4d539faf7f9f652d978707b5ca1350d75f142822705bb89a17577328f5befba009cdb2b9bb9bc6aba36a363ad9c5cf829179f60e77ec488867d405d0020c3bc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc92eda9e45bcca1b22457c941a897b673c300330f7628d68801438d7f7d711f00f79fc725a8628a99c4a77eda710b500d0706104b917d81e4f7d22652811a00ee8bb0c12a97b296aa204f8369df6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13569b535edad1f21da5c5c24bae02883c8271faab304c64b7f372a1c7f0bb28e0f4196f6bc6735c52764268c66f756dd84dd26a3fd112f20432a35d3336b0c984d9517cbe62506d620cf786904cd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16e5b36c8131c6e3824f7a192e2be16eed376ebecf84688074ea76225e082634e2e6e6fae01d19da315281e69da6b699c6f3246b2877f8487cfd53a47c4e219f5f80b7c5aa992cfe8fbf0976ea9ac;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2296c80646aa779664f55d8a5ddfe20d56583469583c9c798fc57239d44d679569cb8498172ebb08192953cd1a39912b0cf808cc050367ac6fb77996c9213eb73998dcdb54980500eb6300f0e83c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fd24b710f304744eb8662b0c7b8a31286982197b629391b4f8d845d84843ea5bded219982eab56dd58b968a9dd94d3b2aa0ec1a83265ed4ebe4dca94e33f170f17a12e6cd69ceaae9806d99f0c17;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcd7d43ad2fff7eded67c316b6c351d20e21c137f1aa5594fc894567d2951154412bab8cd6cacba2c7691445c04271d0f6217bca43cc3754f5ccf202823ac7c6bb3d3f522fe1de9bbe2fd8c5be317;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c4c0d2e4dc80e08c22d3438b59b81e7a57c6161b8a4351497f406d5cfa9d9905bbc2d3420a20dac1784c47ba792e8719fbfe24e13a5dbe2206090bbf80c9891811536c21ae4e757d80f41fe754d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18160e86297c0b39e1db62c5219afa0b741df89661896ec85646a0135d0c5c95e728eceaf01d3e806ebae93743d0be92e1acc5027794a63288c5666403208502a27afa96c5554ff89925fb3eef237;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd5b3bb18cdf4bb3ecc9a6148cd9fa1c9ff6cc955509046b97667c8230ed5298354ce2e6fa767abcf22a6c326b462404746ab981bf2119f1e935cc9813a6d486ce9d06346738c4765a5222cae8e1f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1264003d7c14143fb26230b3172c312922c5ad346f9c6b0a3943a09a132b8dc8e9b67a94746dec278cc4f14cf5172c1f93ac5649e7aafce1fb2003bb75f6a1add527dd67145f43b4c828d876f7812;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18a6eaab3e90e611cfb96b44cf19dd1ffe383d3c6e4a1e08ec7e05394800e925f26233d9a525ce951ae928b636ac63ed3cf2d84b879ba7c967231d0d23ab25302bb3ca663ab8a5e8071b0b58ae446;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5983a05186c5d15ee2e1ed0016b8c0e939aab96819af2a86ab1f9ccf29dab9efd1b6d79529861bcafa7d7010cdd58acb20520dffb986378b4bc672d26d572c42737dec78cec05cdab8cf2513451c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h53bffcb334ecf7b7d7b892beeb4a4e682e9375d6fcf7bd2b0aec648630f82c6525f5211843a7ee44d25f58e70ae78c11c1ed9203469b382377fc939c5083d9383739fc97841a1860c1f2092b4a34;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdebf32e69196533c52b77d26be032147b6312057cb336a2dd5ad7d6c2439013f909d9cca7442e48c5bef9b0cbf0b2dbcbecdce961ad4b78f4f3eab7e44a00b3d1e704e47dd9aebd3132bb80303de;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h883e2f0f5e9c52dcd797694a5017489135d96ac1cc4cec33e4cc85034731e1ecea97e51a9e942e6f924e7e3d08d2dd0470d25d56d80f05e3a52112695902aeaa3d9ef289af88caf05b62ab3f97c5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14207215ae9f2d3aef700740a1fdef74f1b91343ce15f8e11189741ba4097f820d85bc19f4f3f95cd6937e2fea265aeb5af48f5159ade8b629062eca47fab8abd07525ab3a0b93287abd580450220;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18f256a2fb00fde05ef1b7eac24b892e6c9606fad6d61327dc8f3ac7b9a15a6a5e777f33686485cf11322d62995b0b6c84c2248d971bd7f4116d6cf34d4ab5c167cf126cd1c36203f73be3d286366;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18d08e45b9e02c6cbc160f5d952e5c86aae59cb61d4ea577f0a4e657ad5ed4d029531927a7ee9787f47a6a84cf1a58c55486a6d36dddf45740cdd914a07e2eece3eae390549592a4d5a8826e8d079;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1025dca8b3c5e4b57240141a67345587728e97a8b985db94e7d5ad81b9b2a99770f5f3d7947b86a076eeb9594906142a6597a039a3f55f1f45050bf5430b9885950766eb9624303db2f37b0d25099;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17c5b04c548ae62310bcebba6f37f26d877e899e96419fba81e9a272ec1a2b83ef3fc9902c7fde652d4cd745dd47f5b9c2d5cc622b38edfa60a216a00aa978b02202e5ff6d16a51c934314226b9b8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e73ac55944325219b3928fbdeaefe81f9503d5df153eac485e89b96a0821b3722dd3d17eb87e7e479d766423795adc133642b422cc4b91c54e57e876c8025ed5e35f5f5c8e86e78460d84ddbbce;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h155edff810259d280037fe028f1bb265b61a8231f36b5cb43a12de433950fb06547d25e40c488b7ebbb0cfc8af61d80de6cae42c4b5f2833a3afff8abd16df704d55ba3ca6755ed66488b5f77265f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfa592c42b32a71c490ae568bd1119af0a76edd53e7538795596a15ad4f58573f9005cf75e0f02b38859a85fc74e0ba52781abad8ad9e76d62446ce44adab3940788c2d4f07a3cb39373f4bca12ea;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1603dc4ccee2fd14757ad657d380f2dd591386606174e05a91f9e2e306d4e03d4532c3aede7837ccea256f97a28f4b5f64470cdb3023ac03af9521e005c2be057b34049ee0147475655cacfbf5a42;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9e8b1f363118ecf2d93f7cf6fa2e393b9907490f49898427cbf99a0748d6aa307a459370f3d2fa97d4a731610fc1729a6ded630db17fa991577a2b1da203a30f132168c77be7dd1aec2573b84fa2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h48036948399ef2faa6a5613deb481da4a5454225dc3db8cc230b3b12f402e4e03b437364d744485f14bfc1e924e6b0b654c4b8a9e59de963421331b65f78ffb7a0f1cd682e928e66fb6af7d1748a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc44eda377b2d2115d3f9d36ce6bbc662294fb6019474a199579017112e172480e006a8d97f879155c70f7d9c891c2a2a55dabe756fec130c2bbe70eac115bb8d2b27c4d87b861a4ffdbc9ed78177;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h96f218bb3eb28368146b9d88266a53b56b436042a299c25828dcc8af81d69c2ebabbf7c84996b471ba90d59ce13b19a9eb9ce4ea3a9a84f62672063c2c2c2c024314658098d34e7500b23ef731e9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2cb6abce3509210c2eb9e16c3024f29708ca2d8611fcd3b8507822045d7089b0fc0b510bab046151da97307344da672c5dd5b939a2a7b46e93ec1a70c6b27aa6f896bd0f826a47cdb688e3d1922c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha1ba5f96ab6b35dbb0e08e755257093c3637c85a486c5f96bf56ee64b180bfb2eb86c8791df03a3d81a28e7a1113827b71e6cfab36f177f4fef2e4e16a5d37744ec498d0e7129828b3197fdeabaa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h126de5e083813ed53343c225fee1b1d93327ec0b98f42e2cc108865602bc4f13587c9f6ad5ae96ab5d9c495ad9d4a9e099a645d8f517b3648e001b7a08e363dfa0bc61e615cf90321aa68f4611d5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h116e5e09950656849bc932433be70808bcaa6fc9ce9f726489c0da2ada69a2139e601b307199d9986160d09c197fe57927b7976e1fc7f74a1b704f27f6bee794af013db6455cc598d5bd50bd5b5ce;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h754a7696d1fdd262c236202cf3bb898709d32eff7769118ff5577de32a310fd2b2fb0d5d6b259de494fed28213d0ece2999245534901da02bddebddcbb27d0250dd92bc06be15bb0161ba2469eb1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h594e51e7db1610f84f7a3b027046496e9fe71b11c2ee53074b4d65453189d78b7bae05aeb06bd45743bd1595d443ee131ecdd78fb064b8ab85e9fd467814e66b1788c15c69410d5f6162d6486f68;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7ed4131a6efb7982e1d4783f9e70b15147d81a7e9b0da37c8f8e1c35ec2260d816fd0d67789729a75f072bbc7ba660e32f175d0a437ab52644de5ad81fe459f0ac91a264e1243f9bcd9d541d66f0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h462afc24ebecb57b88a8571664010bc82e3dc36bfb6935292eaaa1a9dce469d188bef10683375acbe8b9aed8e7eb284a8e3cf05f109dc5fee595fd824effc66607b08965981d103db7b12de31005;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he4fe37b63836748d85ecd37d32ed4c34a4f825e4e2a492af4bf40a162e958f98ed6f2c2a77f05a04594c3083e6ce3547fc3880689144d2c35fa40a99b7242e650b59907f186898a26f1363793961;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7e22567fd2ff6378ee6c826da28de42e7a2d54d3d34c80a1797302ea582dc93246e8f0a552e7dd709962ffb096bd1e3000eb36123abd7088467f4c960fd7ce3ed6752812c25d3af0d39ed45faf82;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19a69ae29c7b7e29a7bc5c1382dd73a0647057525beb5bfc9c1218e954cf0fb2cb83bd6df0d5549db32cf0ab352950db858573e96b9f1709ab950b9d14321fe0999338175dd6129d43d83e2d5d6cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e3fdb89daab861a8332dd109555938eb7b9395d5785c79111c1dc88824e16d0910ad7cec768e76bd817a2f1c8cfaeacd8bc37753f4e12610a9fc349f14fb205b6e6b537928aa29119c10fee30a27;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bd76e42b6fd7ac7a9b8a86cf3e41b5fe10d50bcf082117af715dd1b1f6af3919a85a3a864531a7f09d133777960a83d4ca81b6b8cab521f66cbf091d39ba28b58d94615789cd4b00986cee402069;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8bbd6658a2736d6f1f5069fac251d4696727541efb69e943d97ea752c160bdec4c71727adc1d36017df72b98b85d0ce5f3426051d2f5a3b8d6d7e272285f03e0b72393aad7d2cde3ce0c7268074f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12110250a23657ee730166c85183d7810859fbea7d9e308cd91321e9e16c9fd5f9f784af42343d0654d4be4775034bcf2cab7df3572041248f4b425d49655328a78a86a4fb4c0da9d3c19678269b6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h40eec4aa536e0aca699b06b7f6b41d5369e57a69f6c840684ef832ccdb231c4313c12e58cec6c9e9dc21340755e01b00201a3875e5c5ca2edbbc70e411081b45d17a8bef50f76a04dfa043150d1d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbcb80d83a1930e06304b241ebb9cab62073760b93d917170dd1e4da9e3f13c6d6cc7e5a557e8badf8f3e805a8f5315bc14a2863646ec7132258e23ee7063d881ba38925c12c58069a322cff7c94d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e74bad9b26b5d8177e0dbb2f3fce31873f596eecd07e8d8bf169da3538230094d4b6b66d6a132fe704893e8a89b12092ed494610ae6035aac5f9d820dc8a1db11917c9f1bc31dcaad44f94c9104e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8fb7e48974898c359abc1dd2c7cb1223cfe70bc23b5711c67fe3cfada9008f82e32bf245a725756ea413acc24621d3ddd035b1dfb3feceb8db61f899b967e07aeaa7f010e41ff0dba481daf688a8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8f92b7c950447b1730f01eb0342ead9e9d6e6321ef182d4aee1aa4bbcdb3f37cd7d498b30929c532f36d8a90c5dcc94d9e742f66cbed0b4a4f82cf3e754f061de9ce47efcc2564e8b6688ac9b72e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf5012a38303e9eb74805c16661163d4dc12edcdc6bac8bdd5bf12cd1a425fe1a63f9b30dd7b8315040ca87c9d73c01355bbc8ecb2d1e0dc7817e59a736a09e528ee7ab160a2b94e77abbbf6e567e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb0f6bce190a55a6d7d05f5b4eaac643ad1ac46b3b3e582cef48ea68db0c1f67ba2d859a0fc9f0ad74ac85ccbcf2bcdb7e7daacd421c1f86c791626f547ea509ec1510e260359196f6ae840d3489f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h108c2e36641cd522a3b30da4b235f9a03f2f1bdc38ded450e88d17dc87d81a94227199cd77295bb7aca1ecfee08d07408f98d6e25bcdb59c4ad64389ddfcdac60030d2071142bd22bbc6f7319752b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1930306d063d4f110155c0fe6e20b6e9106a2bb90d7e8327ceef93516ac9bec414aa345f9ca954fe213883f4830c02435e2334a5acb889065994d04b059518e6a9c96bc5edb0f1fef29d389249dc8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h93a9d19f96e6a5f8840787a37e48edc4e6ca54066492e9b744403d8a7f83721e86e4507ab64ecc1f7eff91e64489fe90306165d91dc4704090010698067d6123f45b48a7f2e2532e2466268f3cc1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha2a35093da4159e60ce0024fde98f662d86d85012d7bf4ed3b51556a3128e8a0fe3408cd19484ee972303a0bb0aa28041e6e060c9142a09f42fbe2b57114adc6b234c6327ee077eb0f4c964f547b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2fd27e9a61a540371683e40ee41182c4c018e10e041bd50e58ccd5b5fe46581aaec5720541a969c1fa391bdd2199154fad49565a829cc216e8171818a2d82c21beac17b58dbc21ef86bf6883698f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h479714e24db3accf0724f5c03a197ea3e669e81d74b9bd27f9a3481ae04694d7a5cadab25f653a9f5cba4c8b94fcb66152d6493d663a976c29d829fa079b3f67c62d1f670c24b2f095e43dc3af79;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h176439d5c401df8589e296e5d0143a00e5121cedf1596f17fa6c0d1daf1f7dbeafd83fcc061bbd79b5adcb33ef32590dc917368bf289b5d2824648175c3db6eae1a9d903c28d834f874fdb21c392d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1806223dbda59f67f82d4f74f7f315fc0d9437194215531b794bbb84305baf3c4fca78bbff5d960f92e221efc2b7686128bf206fa944387391170ce700e863cdcffc4aa6b0af9c7df3a825b7631ff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h54c8b9fd55c0810cb67d8b6c5e3172b5eec261efbb891dc9150e681d8d2aeec7826f6f400c7ce8ad6f17a159ed03e84a058c67245d374e573c519e9b6f7a8c66baf79f6971fec3549002af9bcd5b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18abd1493e94032278ff2444b81f43fe5a0fab058242ca0a3a0d99679a47450b9c340fd6c9430c0cc4409764655668d709030036dd17a438d0717c327503fa33c97ed934e8ecf7d652b028894cceb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h88e579ead04bcd3f4eb229079bba18df653ae9d8b2591b496a52fdac6433b32621ea2753726dbd6b478a9da8d0a6423fe90a7b2629720fbd998d8bd55c253c1ce2e67025ab2ea33483f127e34594;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7b727ae291f31734685715bb89b6049ccdc71f24fc1aedc6f1f795dab11e474c31ba1dec3c1ed0a2d884a81a2d8fd3703e3d21272c523b885ef9d60b2f05cfa1bc809426ed875c0887d77620e923;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fccdee6130e65bc61772b4fd5fcb411035b6f07dfd168756fa4c49f2987773af2a511dec1ed108aabe4ed4af087f43e2f293805624642fb480bf6d856cbb375b047de072b6d73e772f6b8b373216;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbc25a2cd532fcdc4514dabe1e4cdb68c984cb60aad09df10fb3a12a19a31856450a5975fae1f8137ba566802fffc00abedd60dd8b30cb41021c58111b229b0c47ee6e5e88a02cfb7c7ae4cb21e18;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd55152423d825df6f6797a2528065b924783a84f9c281ce6c8e0c2277e7246bfbc3bfb01412178073e489008b453040b103ade14e174d5cdbfceb8876912f9b99b1b2483dbfc15ffacd5bd78ac75;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a8fd29301492b0d7d54a4531134fea078d61f7c0d0e1f8c681acda56773c4405c0f56258f6df29c2797905d7266ccf62c5ae1b83034852580c02fb6efcf9cee0b6b90fd72bc76545e89dc71c6806;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bffd15afccfb8f4ea8b9ffb4b37a0bc80aaa6358d61f6313e3a282b2b49e0ba7f0032e324e4abdece32d44a8371a009878e43f317effa097176630293e1fd67f079847b01649556050daa2f6aa80;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he999ce67abf73e2d4a3a39fd08d81be9a1cbc1f6e96720f153c6e05417b947516c4ecbe33ddc899aa5baab4251f54c76e136f0e8072ca8f3bc00fe9ea23fdfec0a61943bb647bfce4e18685986c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4f69b897c17cc1e40bfd2775a16ef8a9897971296054496873faecef8df0f4f7e10cd31e2d8166c03e6a1f5c64f581dad05cb5d836a7dabfecc818c7abc1d657ab6655b3776b17b0330bca76b49;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1222ce5f2ecc7c3bb3d0cc00a510c6231f91a7e0ac20912ddad65916fb2444349bcb8c76e3265ab3ed62f9ae6dfa52c6b128c436e7c3e686065d99fc48a7489866ce14802273c6eae206ef3a17a3e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b5748b99dad20865cd573000f1a0759266c6b1a144a81f28186aba52dee2da03f45a78a067a23096b2a9dc95e222303a9ed6bc3b30e0372dc1e8cb475774ab9467ed217ba5071906249425e320d1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ac6d7044f2d39de8e3b0fbf893ef10b3260d3b44d67a17e21592287b66c5811c6fd7af56a9a9adb013434149da703c957ff4367e5f5fff7429cddbf341bcc20f705415283b62a575932b44f571cd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a992d1138c6e2c2ad9921179656038a8e9e4682877140c85b70691864942c00ee0da99f42c0e65e30112acf8b13f3e9a1de356f90a90616391d2aa125b94a6440b8a034234dbb66c2b3cceff6ddf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h153e712bad04fb296993ffdda046d5a97ae22d2f57d2651883765e738596075f6c57418e2f57fcf9159d80bf0c7c23fef001c5ceffc443b77cccda25dde2a9b1d8b653f952c6e4dc6555518058f47;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hde8886d37b4c0ca9aeecc35125c6925a242765b3ed6e98f1afbecf1d312ef78df014cda31310829ff74000a52cf96072cee810b8152bf1219099eb1025d0ce066e47f6af96b174631235c9932336;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb8cf78140b501fed97b27722403bfb583e9ce16abdd46117ed1deed07a8fd5cfcfd48d408cd601fd5c3ceefd975346613339ac633640ee1e8cc0fd1761275d88821f3ff433d384c017e5134f51ce;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h72863cbe45abf186db4bf4028b35ef84fc9967c20c40494f9c7c5ece629fe9882e922a7b097af0ccbf6e4c5268906839aa3a6948d81ee55b7aa12f0a91c3de108381ed15079b9c54a1d7930b382c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb866ecafdf28eea5ebdf4d0f8679b899f366aec6b723ae363f50c809bb1afb1f289c9f62d7f10c579463a90285e8445e67a87d1b3c914b24b92d83674172733290775166bdd0a406f352f90bd44;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd523db63dbc392dba8fe5728202705b621a9442f19db857a916ae22a5b26a839638fd60f45772b89a40535237a6c158095054ee5e4cdd8788e4fac205ee6deb621651d11d56a8ebda9437fdc521a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h107dea32f1655e3e20f617105160a872c8e95a6becae549076a689556c3570193a4ca378ba575e608caf1fde044daffc8292744eb88cb83f6178f66d614506bfefe038385247399e0026a12c2e96e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h108e93fa4fd84e52c13da02d1d279c9e6cecb3c0ad831757b5c6153b321e65e28d8f4746cf08677242da13150fe8c5194130507369492a9cc107c022fd74cd5fbd03d7c1f988768335e52ad291db4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h62520925a63ac3f4e56669beb9f570c9e8cddac536a1799174e5ba298d4da1a3c8e5523511a61962cc9d33d4038c80ba4d7c8d5a0336913cec8e0bce1b70ee09ea7399d14bba0c06c352d415b555;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e84b47343594c7880ec33a953c4cd96e3d73bfa00d2ba22ec960f52f7e95d9d8551db488dbb3f18df19820d22cadaa83ce79821bae886711075383a03463e13f570d086741792ef4dac7be8326e2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e581d30d1e59aa013492c807b62b54d4c5bc10e8bda580abb2e4bb7fac77d32fe6a01d6beba0ee02eb8b315bd8a5f8974877dc3257c3b085b2e37c7e302bbda7d71d6279089c0a75b3c81c77ea0a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4cdb3c06364df69923a6a31f90bbe0d19c7cdfa010475b8c47aed5c699f8aa46f8ac7fef96cf69ec0f3c9b229186b1878b796482e4c70a33914cfd5d03da034a1d949aef01692bb4b1b8b255dd49;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1da30c77d93c405d5a690f046c1607f6b8a7f7a52dd3dfd70e012cec59c1625383640ef4793fe6912616b13df87a7269638cf0a1ae7bd6465ea64e64bb34bf609d9a63fecba2b8bab123fbd74d787;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e9f496351ab53856b960be659bf0d02ffef26218c850c37455846319f953905fa635416db56159f7fbce5e396161fd04ce74bb510e0e4f6a17e9a95026589902a0af0bf63e15956bcfff03944a7b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h184404d7ca6fee7303c996910b1559bdcac7bcfe18cbfc038051ab746324a90e26c0ccd2a55f1260ad736a71eac1a1b2e500c87ae45030e9aa42f0c03cd0996ee7c082626a2374cc8210d4061f41a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb7d3c1baf53988306e13d277dbb8418cfa3c6f4115e0a84a8b1a6f85dded03f26640ed472abc3e13dfc7d47ded7ce52874389da8c2cbe9679b7d0ff37a36e642e47caff548f3194620e492157b85;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h148f2370c4cbae294d15b5f29c0fe8bf31bb64dc312ae24368b27a6d16c1f8407b3705c404b84feecc6cdf0f07901ba0c3edb2a9c30794f0ebde295bb8437728d685055639d960536bbec24683012;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h129f6040c8639409978bc92ac93705010700560c56ec78e001f0a7355fc51dbca47cc84b1717d869fc7d201897fe6bcf2ecf0e455529edda864969cae1c20c2c6decc2816020870138021e24addbb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ae6dd2108aa0f317d164814af0e99be93319512ff09b511b60d6d0b0923bd88be73e5834a763dc7809acbb9d4ff387abeedf9192e380ed0cd3842ed4d51cbb5926849e35271ff284a16de9e21e91;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h176d59d40adb8df6972ed65fd51c69a539ce5fec25788d5c91dcbce225aecb342da8aee1e635bbcf94ee035f3d798743874c74758a67524d77a2b5a304e32aeb896b50ab57d2260a6da5cd27e73d4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h70d425f49818a103b47ab5b782d15cb00bc5302834bf20fbe0ea20041dbb9e6f4bfa785211dd30fc1b0a5dc9322c6e71605d739554a23a1b75fa0a638e72366065d80eb5eebee1dd9a919c74a940;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15d55b89b5b23a2b3c203e247166425984a891149da44cc4159a9b44cc5d07094237b1c5bdc4c54a88f0b52ff4d40ad33f4c9c76d65e8bc580c71fe2d9ce463a7551beffd8766cb9e05cf13fae38;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcb32d15527b7be55e446c0e0ccf13bd1a06fca600ab183b284db0c5b9676ac815b05ccff565eb377632c167655af96b8b56376526461a64f472b4b422d2ec501699239f4dae280c184a37f8c468f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13c45f2549125127df4fc8fc3bf20bec6be412c99db6b8a6c5bca9a803a61c7e1933944549648f87ce2c8a55bd7e2678316e91f468868016815cb54aede8ca44e6ab944a73bb4ba35c38e3907f888;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1873da087732afd70ed8bffb49b8bace76bf0bca9eeeea5a740680e6b6ee2d5d0a2d8c39ea45469bfe31efb76ceda7313d742f295b47f46485473c5cad95e9e9b1c45c78828f9d3d94b7e008faa69;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h20173176296aa29529a33cffb1ded9b6dae60e12fd7881afb7bc971cd6faccd41f0e87378da4e0ed4b5a37192d2b6004aad605097b17dff550501ad492595479dd732154e9d9b7af6881d321b237;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fb099aaf5b8ea1387deb510e6efb2d67a57c977937fa2d8174097e0e5c4af1c991da3103d37111ce9806edd9823387825f5b3c379e8e368b99311ec156c03df9d4f422358420cd6375e8483dac8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a20257353f2c21a585d58eacf774e25921c5baf3e18650718372d836ee607b2cd517b704b98ba86812a651c9941bc03fc0df72df8b73c21a6978319d3693604f28104a8ebb044f7f81fbea17b1b2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bf0ddd91165d8f76fc7cee7235b27f9d35fccdc84bd4a422487213cd2cce09ad5cc16d1b8803f26e6d02b88098a4d2fce4e45da13d540804be638895d818d6931c2c17164deb0859721f4f76241c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bdae5aa3f2900872c504af2ca6fa518f0ed936af54525c6e95183b9b3803521f1cf66b3011b94736191eb62a144ec8ef14d639b3ff64a062dd49907290555995802696af42fec7e68643a4f08a6c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e6092218b017ca4e3c56e006196e18274243d0bd0e5667dd83ad4fab0cdf2f2cc821c637757058170c050d10a0f7928c58423ee6861b14dc9ffe222c493b9def7544953b4fdb2154c38d1827a29e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h121bdddae2d5b9148ea92e5ae1d5d10dbabde21b924e8a7a941f00ae5a63272daabef0b2a2deb72210c385fa2b04ded183124e92bcd28b8a5c99658d3fb690346f54ddccb573907be806833ed51a9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13105d82f48f4ee04db1d85e7852bf45281dc4f50180e765b968df8619e6a48994cef90d5a5a1001a6023a3e363c3d57dbf12d545f877eb850bfdb8cd2793848f68bdc07a465dd0aa4ab1043d1b62;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he0aed4ae6cf9ba97aec12ed8112e603a0d08c9044f94d1da1f7d55d14f86ec4634a6e6e99ae80fc984670213c0670d0e5396a8621d5c75cc4612e7fc8ba503620b7a25d413535e91d7833c5b08b5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1afa2d8cde5cbcffa1ae19fdb3e6943ad6acb0d01dd8c1c5e4611b96de66084fab492311e99e46524c14568eab94d12943398323909cedd2cd560762c796982c99201825d3a419374df20c9ac38c8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hff1730cbed4c9e1c8150ba6da0231572745ccd58c066129a762a92cffbb1c41c80c700e2c65b681611ec010ecb239053238c8fc953aea0a40aa6b7fbd35e2e16818097c5af055e0a948da82682e5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fd2c1fdbf0e4b3c5642341b897cfe1ed50a18fe34b7026f9b6f232b5edcf139942450ab4b7567f1e7ece3d535f4da83477c050af15cd816e93809e0fd39b73cee30c05852a0920659bf0ed2273d4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b04d8e3aa1623ecf3473f44b954f7212c690b2a59a90d7e22a32417d5444818292d446ea7fc21b3a4ea4c8a87dbe2fa07e4b2ba62329059bb3fa91f4045a5eb8aabf0bb3a91e7b1ecb2fad8371cb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1349277d0b18fe367d9f5f4db24888f2f22bf4ca5ac68284bd32262b2823dad511038a22d6f82b057be5931c5e389b9285a9ffba4e196d9102b573304e44505cfd9b554f8113b55e8e8d01571e87a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h795457b4ae9c3b8e6db5ec56efba2e0d3783f394e8859ebd4cbd7ec61fd5260e9ba3ca3d29ae08e962bff40468713c6cc9b10f76d7abdf2a57fcc7cc2060d9d1ab9f7ecc9df324ee653172321ddf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10feb6b83e37bdda984780b64d4874ddde644eb67210b70ce99eb3649f14fd1b705e1f15da9429b219f9677e888f1627ceec0ac86a2ceb47c2d5c0a3646d46762089be4bc8467ccd755b6c60ca461;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12741e1a429d3cd3f9a51ad701ea327436b4cf6b8510681641114dd4843785ebc9749617514e5c364d7de0f594b655c91bf851781c811100d3b646704ba646f7045b7ed19312878258978229c355e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h284e1529e9ee0235caceecbd35c5742bf65e69f777535f580eacb406de58761ba0d82965bac1ec81e7db037db171c48d600a8bf49718140acf6737cbf4842b15be32f7ac0faa5db6d9f11551265;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f18997fb531597995bd738138d4302b7bb47d8c5d5c655c5d263dd50c8d966e63c24e29c47dbd6b9085ebcc75d0a24b6188be1a52395204122fa08c4f1ffe6f46324f94879fde5ce49be7ced051e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd952c1013f44d5bde07fc799b92271c5261b4e39b52197a5aa2a36c4c22edc35a121edc6cc2e3d2d733d5aca4eeca0b94c8d7fb99cd176baa73634ac84ce1fd977c7ac163b5653e8bcfeba27632b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc4374e7721de4c35bec96bec24514913b82d19d062e93c277dc6041b662819c8b8cede9b9ab46a2fe9fd7f41d5856a39bee609c85de3d636a9554c9a64919cba26fba19bf5cc9eff376a09f502c9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc7db3ab8e8025ecadc2685aa796efc750a9766d2bb3cef68394ca2568a8d1f5eccd454ee472ee8c0f7efe4f181a8ef990a36a9521745efe48a640f3942c8201d8a4ae5fc8f79822dc162eae81dd5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc9495501f4288931ee866bd566fe0792f132d291ca5a40b00ca294fbd889262cb08ec7e8b24d691f725291dcde81610458d6c444db1c840ecb1881ccdf0d9fac1fa469ac6f9183cb82bce97e91f2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he96541ab2faa55a74169bc15cb366751e52804c95cbf8edac1fd943b8ae26ede6d84ac610862847016da2fe4daa6669507cc2709e7e281a78d427c1f956763c644697945a247f651a7175ccc188d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14686e11e92342100d3e2744479d36e4ff7e08c6d85c3d097e4ddc3407e44f68a90b3c92bb9d574e2e6116a6eeebcceb7a9f84bd56cae223513c4ed3465c2f23867111eb7fdba5874ad83c3272ee9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4dc9c3bb5da3c8b41533d9538e590f3786aefa83c41b60ab9b38fd58011c5f8831f5b9c19a592eb610c9a6983aca4cd1f7f4c51544ceca571710d40c8b54805ef47fdf068937dfaba02e19d04005;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e58eaabdcf32654f5665f89355842ab187637306b23154b1244a22a363dc387b80774ad80436a7436923197c7db16515100c12bbf9ac984fb7e111e6fae5f4b6aaae6a4eb29e95a0814360ece91e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c94e0977741df91f4e479754422640032e590b5a92150cb915034434496c4a4a115e1fbdf7b3849df3c165ead194794300ec356fff873e7094a665a5731043405ea652acf681465e1f4a053c3620;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdd75507b17996aed9e81c9a2b7f0d0b7e12e12b041a6d005de685c7155e8ee4a2708ac6cf9aed175a301c58feacfcbec9f1cbbb77bcd68f546e80f76e285c2cb584aef16332f637bfcd7fdb7182e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d25c3191af85a6ad117872176e1ebe2370aaf2f15aae04a5c9eb7d59558837ff231f2168789067c456c7365269d7e78231cacb68173774850a56ac0353f3266feab367ad11dc1d0616a455f55a84;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1968d8545a914b606717030e65dd1d377141131a7c6fe1f6aaa104a8e44b775fe8394082943fa4c08eaa8933aa3a259e73fcb454106ecf0eeacea708cf76f306bb777a2e079025574f13570a25395;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ccfa58ec6d14b4453fa23a4c5893cd077b35df8720334d0d5c0128fd2b7c7c239981a5e40741365c071a12cc08f5139f5b1f19172c23d8fcec388454b1cdf16e83e8f8a9078acc7d66d46fb8109;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf742119d7a40116c22cffb8f82b1b08cc9415c2aaf44117044fa2924b7856384e3f3c907a654c035d5cf93546eb8c8bf2d108ef91862fe0607eb4c058c8678eb5965ba5fb4a330e1df8dd6b88318;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8782f7282c6d89586246c51605a536f0889652e353fa06bd23bcb66a7df5091434df0095d9f74fa512c5d7f86c313c10dd842df557976a2851a269ea0387582ea82b09ae22d546a3782959c4e238;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb9433da883f285fefb3a856f49331f7fe232303f1f2a14270f1c4ef95a9de6e011547f1d63bdf53bd496e57ccb6909bb0058d41ff7d65778cb09ca8874ad1cd77117439b57fdd6e3b494fa1361d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h50ff162dc19b4787180fb5cf56b2a95dd97b22dc5394379797d64261edb51eac13bd86209c42d4a18908281f836b6aba6cbc0402b5e5920cc2d21eb3e5d19b76001728970f5376a27b04e71ef1b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h137abb74e9a295d0b233152546fef0fbf35631a436a0a7ca4cab3e06401accb1ac437475a888cd9bfd6f606b6ed357b96b30a6e1f1b4377efc8a35348364ed7a3b860421d6dbdd3e79776b72b9bd8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b364db8dc227fa7f44bbcaad7036d704ab1742b4fb899794fa3627e93ee4a3b589ceb4a3c00500c18d40f0d4d61ef02cb861262157f2edccaf5aa2eb8f8ee0fffd2cf3a64a0c9238dbf3fd75b883;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5427c471744591c2512f922a3af9c489483af17be00b0e7a510c5cf4c1d99853f4fabb8deebad6bf1f4bbc52f414bc5583131b7a59853426992580bca249bb54d7e83b5f39eba416f17336675ce8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a810ffaa021de3e7d3c065b05b3ff5c6a9083e3513f9218704333747f24bde5adaad36b80b6938711fc86420407947e174870fe92b3e17aaf0c8f9c2d0050a5f0ac304051c6e7c92499d492cda1f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h112b8baf9b35cf003762f6481e4a21447c6425e0ff346d4aa042912e794ee0c092bdc954c11267c037b1f34300003687db696387855889229e66efca1519b34b5d5480b3ef416bedad09a04fcd2f0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f9e8e7cb0db900dbd7ddd30e36ea548b20fe94eeedf0e320af461a2cf3bd74a411405362a3f9ee7da98710484f3d569a8c038d2dca3883070c9aae5804291594eb3c5f2b034b9ab7a1f6005de0b6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h129b974de694e1958ff531582e854bfe1bb3a28eca4fef31d2b8942838f868a4b057ee2593fe1263e9c69a9499fe49a1bd6145ee97b53e48aef0c9a56b59be7e7b7c9eaaff710c319bdc308d7e058;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15c1ebf3da976415276da0dd3abc51e27bf8cb30740826741e91b1a3db17c75b85bfdc56b28f2aa4baa09eeda253faf1183a057688b053a3767ef573c175e6a826e43cb5d208620f1d15318ab4418;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b27dfc08ad07218829ce0adb056167f3a6543cb1abbb179cc3585285532323dcf69ac2a594adc69c22b544375af63252c2b69709ffd0e0d66885acacf7d062b2fe60df7bad0cb2f7d2d34a11d683;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11ad3723905e780fd1dbdc05570ebec5c51431257e22f455cd763789c1a2d1b068813b21b492fa8679ec05f20fe832e346e61aaeebf5c299235df421ae48ef507d72d454400af67d7522f5bfa4648;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10ae18e06fce2fb0b5ac57669d8af7c7c03c8223b17c84e3533acc01faf3e2223e41c81cbf1fa3a0f8d139712504f2644b435626500d723db19d88fd272d82cb6ac5a9cb9ce78c06066565b471773;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bc02143be21a1c95645c216746c5fbcf4185016e5ded9dd691447778b76fdd4a045bd2c10eefc6d3cb4e7622b89044a24ad84c64586d4ff3998b2386d0d66432480d7565511554fd80fb5a20473a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h86c9d171828fdc0e62e5ba810c2b76f3d81080c320eed26034e3a56989ec8a1e84f5c3b104b052fac6e52c7b6970e49ebe6d3e189d68c12658da4ac064dbaf1b45690aa9ffbfd62550f456547e0b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5ccd8aeaf6e612cc385958450cd063be7cf20171223e88a0c239df13305c109a11e2a7322d5f44afb65e32a1233ae4cfa67e1f8315148b191cf79851d8ef7277ff0b6fc4d8288761416fd8779161;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17d68d7393186b44c2ada7c4478f21723a25c76e439017b9ed23da3acb47073401d83ad3f5160239747175d01a6316a2c3059def40765f0598006a77f56423a16b82a659c84d0a8f6ab93d4bbe155;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hedffa85ab806d85e6d07c6783fd020a3a43275e216d6a6aef951a2b88870a619151f741fe2a24250fda2721c6eab8ef464c6b14a1a1eb8384af117e26b34dd04865ed76d0c55192b5951a70b315e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h59a7d07fc79c53bf60260ac48f4b3c95af702a180dab9d7ee50d1f0024a82d2bf952bd85e9464754284bc9c38c297a126926ee0f2533bef3a90e37dd13b4185991802edf0fed03c9f667080ae4e5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8d1f4e3a0c295334435f748969aa74f3e2b031c2c459e626c7921440b68784c7797dec9c626715c9febbfce875433351ca77544ad24e5a661a802b66d6b6bcfd39252137b3df33a1ab792e760440;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14dce55c103a629dd4b8f58545f9519da12f94122971f83e74ad0dd4c8e6580461b34ec0c5ce75459faab02d6dfc9ec34e149196ff0f243398058126be744b30d3b71ac95360a0c8c292ec51c091c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha77d67b9d835bd5656115c3fc7d50a4ef786345c6de5cfd23425524e61a8a42548c13738a4aa72967f848c7d457c59b90bfaeaeb235d2983b340f2c87b45a2cde2c9cda7e17b4c0f31c764861d70;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb72f99f79c0aa253e7c6049e8db6485a0177a46c967cd3e28e02955e3dfabfd3e517310a4ba0ef1af8ee773897ede9527452a4ef93cf1466d70b69ba6cdab6ab5e6e1766bb01ff0312ef55278316;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7a5d7115a9fbd1fe65da24c773243b354c36b31e8c4788db1032621c11b7e94c5210a71fe752514dcb92d7adbef945eb07084e32e21250006226122ed5b68fe545a5b78a559ac3624e7b26ffef11;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5ce6db24cb625c1628ae33d6d010348bcfcc5546eff5eae76ca120d985fc499f9db3e9618028a771222cb53db4284912899788dc77f16aa2bd469a34fe4c3bac62d4c17586b3c60a819288cc44e2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h163fa9b40f037f7cd735a0e618b2d0dceea3488320e351d5c00dc34c0124334d9a24cb980f6aec5a6bc4a5210f7a8acf47345d42081032cf4cc62986fc008906c329ce47688455d5ccc47b1588573;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a3b41f3ef818897de4e9a6c220ef8bdcce7cc3adf2cf70715f7e868009cfd2378e2959cf92c0c1ce51d4d1b0aeb6817a639e12f59daef62fd43e1245f8408f5d23208abde4fa7c218dd99cf88a6f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9238f2fd644c10a1c3cd5a63c906b44292fe19337e80a858bf069f0a7e882c04264b0955c07210eef2d69d5fb3e3426c899505e617cb4227c5fee81ce5d341eb644d6081391e8b001a0146624a14;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h986ab7fed6c30b7e696effec4e8f37e483f21e913359e2303e025b60991120de157804c9a438ce92a13a20e3bce13437e425bc0a590c90799b78f2dd674f422c2d2399b246c1d1218c6909ca3bb8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb9743d812336bc37507b08ef6dfd09f49a412c92ded609809d05111798b71b73e9d3c5b94cd611f872f876b26e41603cc99a221ee3898ce182ec05b3abc4f41132e0c89aba392ca00064f75e8425;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h805ea5a44d0369347ddc312025f247719a1d075de38cbf4d297be21c6bac7c99d149d9eb9fe6620df88bf577970e6400303e009b228cb4853f114200bff32d404cd2278d110bd7b2f5b9a67e10ba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f29ae7d1f4008894491a5d8b61bd1ee4584e5c33744bb289bc0e853763ec4d7ef587c0eb03c42323ea205fe686d88b6b555ee52cf0ab91af8e94aab63f694bfe4c2abe7a80f32b7cddaa15174763;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hef34e7e61af4ba56e787a886f9b70db3134f730a558b69f734e5b58553b6d9865eb570457dca3a2e92204e6a458fb70e7fb25263156fff0e533825ddda5a2e2fe5d042fb0d5e4ca83fe7ea889227;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bbaad4727ee99218dacd732cfe58fc64dcda1116fc35f4f9d7410f3352387055cd137c488d41cabfbfb87db011e45af3ca09acd42167e4f19f618a32564c70e4115060532163f5c0628bb7be2bf6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb4273335fbb367ba417e986eac3a66411957260f13ca737749bc1e596997b6ccc29f62e12adb8b50810def54f1c44e1adfd8f9007088a1de3d2edc782ba8716eadcb9eeab1d1d8ce0c2caafc4095;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9bced77488f656b15cfc4769c5e9ce810b8ac7bd388e91c2fae6039b59e7727e6faade62e0b57cec51de3ebca3ca153c1e6f6a9e684e627e75ee46060fea7659469c7ed87d5368583d885372b5f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he2d26426b73b3467c35ad739e09385182efae3b612cc73ce8fbd44fc87003ab975f0b12ee134d537358ca3da7ab5d68bce537050c3352a787764cb92a544095d383edbe53a7b0074da736e4dd86a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcaf03b254d338ddfc14ae1b70e8d34e9440292eec1dce8754553b2be366b06b3e1bfe5abed8db022c03ce6e8e0defd15b8b729c15aca6bdb9718823cd6824e8e6f362bb78608cf602833dcef9445;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h21fa3af75bfb0a54a748cfe581c6834fc23cd662bb0c648d6ce0a4af6606f283d17155d9a43bd41670a60b2104c4716a430c24ddb8e3629c4914d48aa99261c5cb78ac5a4c163eb4264669082b79;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1706b2ae9ad390ca779686240b9ff3ca32c57ef73133b3d681ed843701adbbeb422808ef17f3563c05c879ad7159dea8ad6938d917e42c50a116c984a3228ed5b1f6164342df3593e893cc0f16b37;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1aab628c6df1372bc43ae07248c13d0ef1ea62ef3ae27614572bbe53608afcba7ee2a4eb0c570f50bcf455b74d4a24495b9bcee57b266307aa2d3495ec7abaf7b1f1294b2d8a5f2b2b239e6295766;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15e88056da52dc028ea3a93964cc44af75f5368f48bb258ee932dda75fdad11d97fe5f0d33097c9baa28b0e3991780c58690edcf8475f0cb9d32f74db4e438cca4fb9d00196b3c208fa4050bec65f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8f64c6ffe66ef1e74db72bd16b29c184ba33dc90e28d279e3b41ac866e6297a967976f4ccfcdedca596bcddd65e7defb3caa2698ee35234e9ff755c52f628db14f1da52c465205e4cd565eb8bfff;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9e79340e958e493b8b2a3856e136a7068ef5c8a500ef776c247a6e34cba7ce98133ccd839b01071659a744780b75c087405323467b30b04b7fbb0286291eb03c7da4148740bb994f902509a5ff19;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2745691cddcf97125be2573c0615ada5e71ca80a39a88ea5a3bb330128ae42e7e9ccdadc60e6b9c1ca604e9d6a23973877b3f3d14b2595114d1e5a87c2ca3def7865cac8505b6f22e1917ce0a1f9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d805561478afc2a7c436c4fa67e3773bce97ca6e55799cca86794c76342f7d9a1895c78d3b5366e1136771fa582575163b80bb4db0ec2a847547f10c9f2ea2b4a612306146450ee4956eb8a6ef3b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha221a55bb89dcbb2b3c97816f035cb90538be033059b3389504ade3a88fe05997d1365edf8c949f1d0fc3d0e543240fb187bf6206f2875fbc3311b3f92b979556b4e8fc6ce6521265902043f2535;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10dc772dfaaf28ff5d1df2abb62d1d0974cad742fbb7f8d9bbaac03488e88a2095ff3d99e2f54d4eae4e9331040b54ae9da507844d412a536abf9ad51eeec4d0149cd421043d052a09ee75e36cdb4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4818c8910ea4e945de2b9785dab4a374609e4c0491dc64c892d0aea0595a51c00967bf392255991b085f774c0cc643317a03d1baff19f8da6c9da61f94cc2ef7542e31b32c4c0bfafd51847e9bb4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h74bd765c8e3ce59d5266c65018ea3c9e107c02a46fb254a17986662ae1f043aadd60c9ab3185ad5d9b27b0e7415457265d916542d5582284aaf196dd92a10e031c582b0c339350d3a2293d67eae1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h123fa785b884af9516cb62be4f90ab2e503d7cca3610ae9694a0fce9dd27bed63099bc3bcf357ea8460bf478d7ca08fada3b164f3898c773ae4839dcb0796a365cce4d5363c9b638a303f349fa47c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hadec9c06b2a2019ccfe38fb6dc72433ef829a45c0b6256a15370c1a018fc7f9d7e0b41badb2623f6c43c5e747374a14101cad49121bcc97692e8b2e8545b0f0b2914faf0056764e8ce5c718904cc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf731a8ca1743914988d4677437918f124a0d07c6382f1cd30c6571da293c76bad846e3632b2cf2fb99bf47b3fcb14360a8beb0151e3e82f7ef8cf9cf2bcd61645f6b573b0cdeee53b6398a9db67;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f2074696b673e1ebda2198ac23dd07326222e20e1bf08f31f214d0ff56ade9373b63c3ac69920d2d17c040f7aa382c87710d884116e55b20f04af029b98808e7174796a20e1aaae949acca0abac;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc5afa7a5ee5da50ff6e28a5040a639ebca8f64b4a87c1ec145295cd0e45673038a6440313ed8437829fefc3094186b8f2ba14a91064cb8d5cf2c4303a15b226e82f62c38f6bdc30045452d94cf47;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he4f9fdfb2b88db59b1b70839baf5133a2f5aae174b2c5d6af1136299c3ad194197aff76d7452df092094b0f1669deac0d48a8ef9c70fd9ccf6141e9bf6392c3a42181429be6fade05e91db1cee38;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8a5d3723f6937d4c2142edc4508fde9eef0d0e58c21bb4221c433d58ab1d138722c96104f594997e3c025527ae8abcb4d5a4fc926a8fa3dfc482f5d00a0bf747efc2f81bebadef1b300c7981db09;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h8bb01ffe4a7fc2a93e11ef99b17583c9ba94d94a11d7576797bd705448f7f0a6ae1fd5c173207f49a2d40abeedf2279f9cc9731241a67202fb0550bc8b063ff30058d4c4e728dca954ce64dcb749;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h89c9d06eab73655064dfa0ec35fa9ac6d6a6bf8b2cf3bae6169e79f12755e067558368808a408a2126d208e7c9ec879cbedfe5bbb5a7d94321e490af65ff51d2f022d3d601fd74e9f7e57d28b324;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19dda3d66a6487df30edb97c3bd8c70242fd05875e47161963959cbdf124e9b9603a8d1a5b2eb8c3394e15e6cb83e79aa8bf47542af7a5cc1246a4ebe2a68b62dcddd01fa929702313c36e43ec7c8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14234f9584d5199233acb657c5f5f5bba398b5208156b20f061359402f2e6b0c3f49652b566fef99092e029cc3effa91810e70c70fa2a6be1158211ac62f7bde15093f79e1986b860c463e8fe85e0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ba5991f6328a5694d688aa12b109d5934b45048b985ff8876adf605e1ed291c07f1b9f4026e3a5cd7a7fe28f975437b4eac17395d9c567752a8e5008b76c4bd2fb7f1ffbc2c9a2730a77425e4c9a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5ef7ad375a5572b1e43ec306138856084e0de433e93b40b27766b9c349b37ba878475fdd365d9d1c854d903d92285a13d6849ee21a7dc228efa9a7253959acae7038af29c226ed504c584533d5c1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h46928d89ae1b24463c407dac7b2fbc00f8c38bbe80b0863fbb143cf4caf912ee63662fdf751a9cbd4f7417148e3f908845e4155e033e66983f8e16ad97e447ed5dc5d32bdbed88ec207b7f15a64;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16f5dd906a2855765fdb2fc54b3cc73ebf52756b8cf0e9aac9e8eb38f0a8527b7b1aceba6bfa893b9d4be27913f6e9205c253e446af217f297c5aa384fa73be0a9e06bd417228674d48cf6873a055;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16491069fbc2b378f26d6ec7c700e7bf7cc7224080449280172969a248f5587c4a757b758a122bde618479376154deb56ee4cd630dbe9ecf41d138b5c2aca38edcd2e52854a2d8b874f7bb091f163;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13971513627e76758515fbca5c98d9b7ca52e0fe38965c113ac35b0c42f0c96dfa3986bc2adc6bd1560cf8078eab1429f759cf55ba2d76ed53ba228ba8663cc35a90e89ab7e2b90a8f3712feab349;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10365c1fce6c091eb1e9fe6c3bac7f09dbb566a2f32afac87d53b5e6434de37e0c6f2fc07a8dd27c2531eeda49a291f199e6a90873658584c5f49805a450c6b57168d4b9a098770d69441e15604d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19224a77b2f7ca9cb5827fc4b00e3615c5a5cd5463d4bb803eb7ecb33171cde181f8a6dc3ec0a653a3746c06209530023e06dc6d98bfd0fe2cd64063d9646ec5de4d90d1bd8957b2a12b09ee11d9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11bb639053de98a267f6b57033885ff53b9e7897a1cc03b1cd89aeec58b63dad6806f2d366d3e27c4ac0bfe896a474ff9cb486be5a2a0a3f3348e06fb39499a20489b5d9410c975b4688a8eec4b65;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e99a4d6f9eedc48266b2effae5c102561847228cc5c50a45fc8646bb0bfff8532b119a3922b29b1760bea4be8c6a47bba8e7c9dc68a9953417177c46ba3e1bfabee41d13e8bfedda46ea84b40431;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h720f2966a20e4473e393f1582692b0442e991e263bd943c3762f40faafdab1ade8ee365ccac630fbe714e57376f3cfdb33c19aff0fdcd46a4bccb882fad2a28ff3f4c25762c6c893e1a46a338cbd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h83ba61816434bcb9f08f40acc90e2cf99c171013c7a7bb0bfed8df96da1900fd0eaae4bd84375897313f28f0634af3da4237f26c467594e0e5e5ab42a6d269bbb8d9a74cda38b248e1027f0daa04;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h498b3638da86e8840bf038916e2f9d44e2e2e9367a7ad38c8803895a9f92f591ffe8e80d11ca543dad68d939e7724580f38853a45d00d2d601cdf61b0c550829b3619169cb5e5989d8dbcbfd97f6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b61c52c15a1c214f2fede560d9e80b5505935e0021df034705c266fcc9fd2f4218933a926f789e5a47dd323d123ad9ebc6ee82f755ba8e3fbe2c3c9d010a7350caa37a892cdb88dba14ec7099718;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2e5416caf9fa30a1cb7400cc16bea8bdb8520310f5a27bb415e3aa97a69a193f4f5dc3281154490945f76f8800ec3be330acc25d388676ceb9d6c98a71289131b7efdf547c514dd60aca196aac61;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e3fbe3b3c106ba3ef2c516fb2ced05be78356e27ed581e227f637888415405379d0482754f4b68e42f9d56b616cc826d9a042bb83d88e2f33bdc0d8c49c597d56891425c3b4277d4ddd0bd9980f4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12c0ce5182975241997a68a55eb58f3f95a201c9a922d2072e4c07a7b4f5ea915ea15f3f959990f526c4a8d313b90137ff006e9a8e80c66b2cc73a7c6f0cf4739db70e984c8e63fc51ad8cae3b601;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17c6287a3cfc9036de9ca0dfe94469fe791628919cd20c17ab2abb0f0662646d382b91bdeb021e61969044df5bb3c561a70e28077e23a121ef5255f9f6789a3a412caa8a8ce84ad166a118b91eb10;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haafb35a3b57bf9594ad8196f07de3fde8ad43c41a1d0509342e49e7c5536dffe09e630a1b13a7fcd2aa65b30681b44090e815fc0fe5366e606de678ea9e8c5c95f007c23225d07f5b96a4eba806c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dffd9849d6c5fb7e3fa3513339b18b9fbcfe2c1a45c88d269a164350e2839cc56762ee229228a424c9280392aba169f21137414ef8f30b8b48bb881cb8a5bb0e8d899a67f4d2fe6f42ad339dac39;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f32349220a4c591ebce04c251224c7725253bdf0d208878bd504f25bd2e2732fd4a356f47931085fe7810970102e24fc0c3b0234fda7c0c8afe25aafae73556bacd01e18c12a7a6555a3080573be;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h137e9096bcc9955163a172ca590599129b5323083dc669bcdacb8adfeab66cbcded8c58f7cf5bbd8a73d820ce0d05b7e7cbf0b611ecafdc5e1b3e236887422418b0b1fa31a7ac366e3c8c85e4e9a1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hcbd47ec07b44b34010dded80d8c3e1b36ef4833a2eaaeed796355d94e7dab1fcc92284889ee67dde5bf39a14fe814ebcea1ef135012d89f4b9ac63a9a8c1cd304ffdc142ae8ed3a63f298ed9584c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11345e8593d56bfa46fb2d4cfe8c423f6c6446ce9fdf9f5f3a2a480c2176e2932c28dd3094233c09966e8e42095ab06342bf10a2145d368fd200e6dd62227dd788c45c0d16c937bd9071bdfdd7fac;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdd44d4b85ba16bf54bb7ad72ccf1483f1ab833737279d7b4c4bcc05b98df1d9168c9bff9628c1ff5b701bd9ae71bafd357c493329cae2a5a337a4e59218f2a7dedbdc673104f4bc064890c870cf8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h154e575ba67fa918150b4b9e4449280aebdea43e2120ee43f67aa53afbc00375b30c7e5cd953d66b580b6b243f5a27b3a1918abf590e4b4355a74c5375cbbd533720fb4640dc929fcca8c897978e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3160c0df5120df28410b68af89ec7eeb4744763df5c63344f399fb04c98d085e76a20a360c1c195ded24b9228cdc9b87058f59ff673bd701d215fbd538ec3020ce0ddaf2cfd08d7316cb84480c5a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h179b842475c42948c9f6796c49a307309c5c996ca41f021a52485582c93be035b5bbe6b807f08da1e023aaaf2b55a0e8404856d81883524bf8eacfab4ecc86e2abb660475a613cd468f29afbdc31;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16570f8d66cead1820527a8168562f72897c5efeb76c50cc8f0288ab51795248e61832ef6142e778f4da05ed905c526ba03a886605b7bcb48fed0f3d15399c507d702b7234258ac253d903f235dac;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18b3572c05249fdec2643897f39284c5b495f555bf386735b0856cd7bcebca17a73c772fed351668542c3f523e446123248fd4fa0c47be8544b567a0b761446931178af209a37aae1e4adab3e70bf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfa2d3b6d40414e007dc1f9f31fcea92e09e9ed0d7233714404352ee3d4cee7499285620b758ac9dc66a5651e044c93925a18cefec35b3b69bec847cac2b4a3c687875595ed8eb9a8dd3a96ee1b4d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he74d504fbacbe0eee3a547af30c00a40f216cfcec883b476026e2c2fc62f592d7c91abed5b7a8640fe76e45d5cc54b64b61bfd09846a75286f05f6f64e97d92121440151855516f1833f9e45d2d8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf499968ec6f19664bec6933abc6bbb67ce21190f89387fc2eeed235e3d8490a2f24ce4294d3d95392dffb8eda06c327adbf78626f09993b1e95ad7be2cf3b1727bfc11c86289b96362cde113fbc2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1a6ed48a41970339acdb4f180690cab3af3d0eb5ea68d8b6de49d919a4f18550cd10ba75e98bccae2007b2658517e2eefd02be40c3f4aab8027e6f3d4b86358c3f1af97e0f17d7c1aa2358d046f70;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h14c8fad9cc2c33cd5a274cfd1f7516b583bf9047ac9a6dd35c143f0c98bd61a10a16c1d3857e05f1d374d7faa34e9cf5d72dc37fcc70ed4e9e40b251ec276865ed46586f2940344e2a9d541bf1f7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'had53dfd22711b5ff17a06d39c4f3674669919fdd29d188bf073fa808fa9c40796e902c60c49480dfe02bf3b46ff1750c4ded1a4410cb5ef24a582ba68d303f7fa462396959e449b975cf93a7eea2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c28800892d676d5d091791cccd8275987b0ab6ec25a65c9c15125116564c0c60c4c48280f4e7c31f4dabcb27d41122670d596d62204867682532dc6bebb350c6a70fe06ac169cb7b3770537230a7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1212b61305857faed4554aab8571340d341d4d6b4dfb8827decabcccc0e38a3b0df48d5723a06172f7439e4eb5b0684b27a0bc2fd960210ac0c04e5cc597f2a76f31871884aeac1a18574509d5be4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12df39d87bda8bba202dd0f0f1472cab1792fb6f096b26965cc224e91c11136b6f9793dfe89d43c6eb116efabb80b7f51999b92bab913e046f9178773237f4ced252cc0ea4f2deb961b1c2cec2fda;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h45b0d4e81eba93691b36a676dec4890557640c3f4a0be9c16125cb1ae08398fdca58b49466952d85e492ee03aefb841166bf258e979afab1743824b72bcf7be08738c114dd633cede6a94b8a0d17;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11635e36dd75d823425adcf2b0d3b6369a40f42b89ef9cee4c3b7d85c7ef196b2a06c6f02cfafcd448ed9c01bfc9083141173c67a2b66e094102937098c552ebc4f3128cb3591a77439e8a019b7b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h19dc931f6ec1ae9509c03e2c8a0178cf1b53f8477533d2ed573f26cf354b91a3b269fe89740a9a61f439e1f6c8c1c5ff484faebc7cf440fcfce31b4ff3c36eebdf6ab4f9453b3ed0d6e227a889cca;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b789ed16561233fdafe4a39c4a874d17b2625261f5d5a8b30ded4198eae81faae0365d7ca1b1994b026102eb85dd3fe0566499a29c3e37a8b3b2e16efa11f5a94404572ddf5ba4f4a75f16d28370;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11a86c00fab0dc28a52f7e3769c102d88299ef80b101d5dc8d65b2a87d337dc01b2d7ccb9320816866d2a867a948faf42b2e7e98d9fd9649818a3d31b0965ae4bf2ca99e8338002d10f5793687ca6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h353559ec5efa9a5620162b4ca6194b7b68c47d2f05dc5ef195d27332567bf559b550809c3ff9b3e331b52a919226b16d7abe78ff6b58df56347c50ba8bf7150b63befaf83fe0db1e0999a9d9cd62;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h27b78ccd87798abdae77d090719741e3d63b621236b3dbad632c8f3e4923d2426e3ceb77b9658298e2896b8fbb10ff60b1e6eb2c67facd32f4a1c4f1d99279c7d72ff9d2b908e7f9caedd030bfb8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hbee536da8a139f0de0ab9f4ef876e24120613665bb9d3595aa1772875c6dd0b7b0a1b9037b076b573896ef4f54cc2720cfb8510022eaf90823bade77f41e40d6dba583032f41537006181f8d6d08;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15940ba29b6d4d86fd7bd9979b4a13cdcdfedff459ef2e9522f7562d04c9ba4bae2c932cb96409a7c6a7fd2415a83d2a941f323888c7d9d7665444c8238cea3cd8f2d1349696470da113ae5d5d1e5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd58d023e9843862d31811603d1d350077d6c129b6dc4e7c60d5091d83e919efcf7304c3aadda2051091049bc3873b93b4a87a17502a389af99b7420dfb0c947475c8183dc868adc556a3133433dd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h4eefbc666b63a7e58d5a21a708ea88e2d4d361853cb6a8311df9787340e4ea2c82f0a3965dedc85f1fc13781b9e5df164c16e94bdcaadbb27f0af24054a4c7603a84bb975b947091937556f0b846;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h182e3cbbbe43df58e7960d65ed3f9c08046937ecb6b2d6127448fc192e0fc0098ca07b6a2f9f78832f5937dc609ad1d1642b4606e0cd67e9ae96c8dad17b1fdc099e248d3f88f07943e5b962b4ac2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c63733cef5f248c8630b786fd8fef6e745646fb8b19ded6e48dd0f253e0eec66476075d0f10f2953fc54a991d570be0427042a098b2bdbd5e850506e3030607df3e44ba9108619a8e419fc3af6bc;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h21ddfb6a90604df5b23d7893c574addb90641a15d61b70bea42f118b2b65c3f7e15bfc5d06674c3c4506d869d7e3272a85357f3e6bdaab27741c548bda14b108b3833be44dfd0ed65ae89555d110;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12c8525401e34b24ff808f1f18d442d59dbe0b51cde66de86149bbd5ec5be226a95dffc2576f2d9eb610064b91d7e24420cbe5551538ddb126801e4a7c9b74880765992d6d656ce450e00968847e2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9fcfe441d9d72d29a9999a87f0582ce9c53c1972f8b605ddb555b0b43cfe0d50716b36a5af9b9b703e6c02808938e8fa51f6cded05a910038e3b5cdf352fcf4a7d25c46847e78330cc86087be959;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1667dc80059d1364168a29a6220487932a133b27619d06128541d0585394ac718ab4ec6717a33fca3c70769d4cbba778e99bba4d4938db22180cc7053780bb566cc51a5a6231e3d456e5ef7883219;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d837c38cfc597cb9fbbaeb42e0ec7e7d8468af9c74ac1a0a5b973291841eebcf6d1d5abc5f20bd0d438d3de3b08ced1f28b73bce3db61c00a9203b42ef73835aa7a6268e24438abad39048ad4601;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10cdcde9ab37528011e6338595fed625b24f99c525878ca4bd69e64bae03f4e420900608cd1c498fa177f0053b92ae387ea7dd81342738ecbb9e6e59f61e2036d963328d5d30ee7816ed54c0ed74f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d4c191707e4c6e2e3e9c66dade137af776d7c40e2ddfd13933cde8fbdf90e4607a6a8b8d31723a39c8225a62aaa8391101ce9288eb24899dfcab09818209805118a839dc160ea16ea18b3fe166db;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h144f5090126882ec21f89536d4e5f2640f0128985e24c2e68372c06e775d362bd04f0b1902f664d6822ca39d9af3a3ecca316ab51c858a2292bfa208f1c296859c647fdab5d98339be36267c9145d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hf32b483e98ff5db3339dd3b8ecfa3bc7d8350f7a781c3b6a4b961e1259342a594965748f0900592e522fffeb1cc18d6fdddb6c0fc41ce2760ee98f7b908e696536fc6d10e5becbd8e5d7ecdacec4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h26c42356cdcc4125ebb784dd843710fb529a63646dfc8693403613fd856db53a3ac5570204647593cfaaa90ba9d6a9093ae6df693c88ee1f69ce9b82a221dae7e4681fe61a75850569e6024aafeb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5c691c9cb638d5a11d47fccf698b539376e95c823cb3fa0a07a50f3656a4f806ab3c38be95f5432728147e8d97e5ea8a95428fbff5bd751c7f0bb48905d301c4e31602ced5695dfc7c303801e16;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1661bf44cb7bb1e00c12c275cb7af0b2effdaa1d2cce7c4cc4b6eeab8011b45604edb0cc9eae263ba274967333c05ec728b18b7d09a5552f711d5c9d6393eca33b7b4a2f520ee48a769ca656ce15e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17cce7caf7089bee51720964126327126876980638776346c04a13cfa5f4f004a5082eecf862aa73b78cecb1da8036cbbc335e4f146eb9385fdd31843ca505153de554043c788872ff60f13107ec9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17c66e054f6c5e0fc810bb8b65fe215e498cf76f5692b32f73a5f7bfc91704e1c90a9fe6d8a4c77902fcf4ac5a6eaf7fd9885586d724b7949efd6052ae28e9a675934ba097341a073ac77e8f2a8f8;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13f09a54cf92e3721bd8c1b6c3915488ec0cdd58a5ca96ce271e933dfd09a2c20da4485a2b315c0284dc32c260faf336728fa4ed195944b834fcfa50a4a0c590ebb1aafedb851759de7948a1f3a34;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h17facd5872d1ff2193751b35992b3ba3128aee46060e9d492abe4f159c850afa8f11e46a1753bc1ac4646de49e354c0884525a651d912dbee0ccc5653b8bbc40d57f8735f902ae5a731cd96a3015f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h112ec73e921b4e120b963c73da7c9885b73879fa08e1f04f24fa944b221be7a21f09b575a146c6ef4da1358d5e2e23e322d6f95760b91406e7d20f4615d87d89327e065c6e1b9fd84933c7e82094c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha68f0fef2f937eabf0b0e0e6717e74651b2fe7882a550546ab265a29aeb32781c10e4927154a5857b09a5ebbd1bd8ee34b2e1500b171304277eb9a73a9e63f5a70b120306f7a5b55d7b52e33ef7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18548ec4b343cdd85cc032322d13cf3e8be2b741fae4a57319a0c5d1b5c04722e695c3b30b9869b7e36d77f37125bf9cf8085f028aa40dd0b0982e15b8e68d245e57bae039a3f94cf1ed33c8b545d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10e3e3a7ae28c621962774a92bdc69165663d5000cc8d2c6809e2d60b9210a0bb9ed0dc704a8cdc3a6c7550d1eae990e4bbb092b6c0b4c089875566628ac53a57bb13d6ba601b501647dc746b013d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c5a38301e059b2c4bc196288cccb4ece5e7fab795b3a0faed7682604e8853ea462a16c29351f32c871b2462953b6957eaffdae14a6b09cd3cbfbd38e3718418cf065d94825180bbd2369e8128359;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h13c2da1b980fa9b0916ad5816981f027f00092bf2d3ce41c8441618fc6cb92bc4be837d7cc9ba78b91d490a9276c7a2f48e51231f9d78c8b7d7006b532a969b1b08bee828c1aeb68eaea6f2bdb7d5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10f9a6754b16c3d6b75914aef1c9bccf4720c8d9690bf9cc421619b7c9464bd740fedbca2d8fa14b8cc65a5ddc791eeed065b548b86a3aad72df670e77999d9a36a691b123e182d4035a875e8208c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h108c98110d49fe3f89a84710a00cbaa395b8aebf8771c18837d4df4c7d3507650bfaf4a948f2aa8b9143fd4e8969a5924a089635732ba274fc7c983c3bb0b25ad9476eca9f0fd58be4b45b99fcaca;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h107c98a60433876c172b50b0464ebe6bee6c4f86b3e381061e84f89cbf70b6785134fd666eb6ba0e54b40f277aea4ba27d97e0b953d38ace791a65b861a9c8baa2c798685fc76152de08239533e4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fc246ca353a22ca3b04b208fba010ae4c3a13ea620141421f8920c20f0cfd3ce14ca4985a6de6923a90c2b7f32f59efb4da133d2f26a64e7f69d9641704407bac5061fa055c2b92ba67a6aaa2c64;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d51b337735df5e83cd55a402eb36f5b158d1b695da25da7c9b97b717adf5e8ff6dd9a2965f70feb413fa81d4624dfd42c9f3eac9e820634327ab6971de61889cbab7dad64e013d5b8c7d0be87e47;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h86d47fc987e864089f4ce70af9388d22becf783159e24d2e66814855cf0fe004c6d3e8233cfa42749f373bf4c8bd2a683ece05e83a5d4de8f88bf905541c1868aa1172012522f7883bfa03462729;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18503fabd048b383099269171ed911beb7ed6867c9d8da0895c4bb7fd4fea2d59a04e86e20c61f27bc641320be8d65e7af418667e5e94965caf53e299e6a4199b4acb57d7b8d692d9f7ded9714f96;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1b4b028f16f5f6041831c9c15697fae705bfdc1954a7c4120a94c28221e33060612dea73d5c3911897d9c51c9787b43f7ceac92c1926f18c99196904d735e839bcb251960b2da1a516779abd4ffba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haaf79c90387f3b8b990a9afbe2d9f8146b75ac12a8dc8286996d564b4751fbd5e7441f1668d8c9e6d073e111d9a08dec80fd19c37f8a038702d0cfc1f88283777c1ce57f4eec49b67c120755da12;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h105600db71a9eee0923af50cf3b0c6e43bbad2c3cbafac5ae2dab9add280fbfe4e49e156b58bddfe9c6a0122e71128b1f19291fcb7e68fbc98ff40cf62dedd6dd6877f8a0b8a2d61430d008b6d79a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11527dd50538f55a15dc36dbd633b4b99694319bf7ae9f6e64cf58354b2a6cf61671108b5303336a3be2edbe2e4c0d44474ecac40d0b4b1d2bbf1ef6e74b41c7c176cc2ca0785d28140a885e1004f;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18bf6307fd16ff54e80d37a1ef9a8c5b0d82325fdd6865e36110e309d642db621746a6ecd7476219b839ef2bc34dcfaf66262277cdf49fcdcb58b876073562d77ff29d81028b3c0c65a76f633edbf;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haca2b892a99b5debb2b9f0100f3f6943ef1ddc913092dbc995488fff869cb0cc19593d0e613a266d06913aaff89f4f6d1cbc11e65cde05ae375e558274bd7be76cacbbb3ce4162f5ac097bca2df5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18cd40fd2b1cc5d119436f21c1ec0a943ae0883fdfd72a6d91d5ebf7c09f06bb19d93e1d7a3951a9c26c0cae95c6fbb4f26a88a063cc730c81e027d7f7634088ff521e5fe456344669d2d928deb0;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h163cdd2b891a294de98fed0f51df63ba3f4f3a33f556e96cf0988a7ea36dde51be2bc21515da13d7bb7efa4e616aa72ece266ad29dfc84c0b858acd8483ff87e2d81c751b0c60c3f35e2f8f21ef15;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h109ce8d0be8f07c3e12af28ab3288765871d4dc63a04fb14e41e5fa387f38a0a30d0ac5c2016edac9701ac31992eca33f76f7b21004d6798e6b80a30a34f9ab29734de008acc0e1eeab5df2fd01ee;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1eb913669dfe92df7da155ee061d4217232fdb890a82869da939271ba39a09de7106fe1b0e795f0b185de000cf56c6b6c67642351e8b7f145e4fe381213b1079ece7b192f917842141cb451bef996;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hfdd9252beb7f386a954d31d25784ca897dd2a0c0615b942e1c9d0cb872f47e4938ff708cf04c26e2f25b16e3b21533df55c9d400058a602f7daabe689c923699712570b493ac09f6ab4716a1d22e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h198327ea99e264f75cba92c24467dfa59673f4393da55e703cdf3db3066667b927e0552d6c5d21ce2f62f09b02beff923083e89dd9a933a8ffefde732748405e6b2af6108c9ebb210672c85fcfc46;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'ha211fa50b547608f8e141f7ca3042086ea71d6a061cae25abaf28ec93316e07d6534266f8f02f3b6bf9938a2caff522091dc76f0c4f2494664ae3fc267c06194dfb8d73b44ec898a1dfa3c14607a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15d06627d76733c09007e40a8ffa6b615865c1866694848fea411e7e947ddc43c66bb161eec20a0ec7a587c59d0ee1580f375e9e54716ba2a82fdb6ee282ce1b08a61ff50b19600c6fad13e9e37b9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h135a6f0ad67325de6d2e1c497c63df3f08d3da946e01f7b4a5afc1f7512045489f3e01c0a96cef683994bc5796bcf61621683847312965058cbdb545094222f7e3973f4b25a066af526472bbf25c1;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he13a2386273ac10ac770d173e4399bb4b4bc114e20048f7cf1090b3f0f1e18d3f05a0c1fd9114689de714517eb8c8fe399b69dd87bc3828690b5030565c27f3f23c6566004b94eba95d6207315c2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h24b2bd577e806386142bd43ae30bdba1edadfc2bc6ace0045a4532b3cdc1967eca2cdf3e7b0f702486bcb336fde6dc3759b2e5e5d3fa83b5d0ce9ce3fcaf2719c389330dd77ef91cd3cce54f6d6d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h12cf7d9d4a7743607a538cde2733c14d540489502afeb396aff047895a4e1e4bd9e5d3dc98832aba66ca5fca74ad1584fb4959120f1151fc33b2e92f27ffce77b2f468ce938a8a6392022193b4ace;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ff6f1858cd09eac910e16b4a26a25315b0d522add020c4c99c54447a25dfb5982f6e5d80f0a713b95f76fa9a824f7776974afafb381b9a3c35007550f672d9e2d926bb681443e2e6f855964a3d7d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h18bf29f8eaf249fbdededfa58483e75022f0a8fb9f115108feac43a584af7955ea28dade3c16d2b8808f8a825889e3b97305bde4645c167bda1bd4a132b3cd1b2dfec1b599d30bb389a6e20189163;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h35abf0a7e7ec183ac21079972a69602b17f9e93d21a52af12eea090fc1d44bc5a2de37838890db2303d92be4f418d24a84fb03d008c3c1906076c0083b12bafa489d385b04f37f225a5dbc283661;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10fa0e055ed32e1f810756c139fde24dec4461ebb8841447e70a10ec058983400c581747156d6f24590fa1f785d1f9c4ad35bd230f5d9707b69c729296cf84dc9e85c85845c00a0d8e33bef2c9809;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'haaba484d80d9f08a94318c61c9b9d99e22de76362871ba17ba206cb3030786e3ce3e597b8ec1cc99603156c94485752112fefe573d2459dc30b0de1fc529df988bfc645de4625da6ae7a9bb5fc86;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1bd9865c02a54cdf7c5bc5ef53d515ff25bff5f0b46d365b82f54489652ef22c67f4f4ed9232be632883df29b9343191f5a80a07c739ff2ff0930c4da5b6f15d1bf7d7e7819c4017747b67cec0991;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1825167cc0d4f389005aeb8d55c44fdca9686c53b2aeb1f25ebe16665bdcce37aa8c2262e233236d2d8c42a8fd1fbc744dd00d4df0154074a8d7c1f77497eb88f45cfe718a93348d41df2d56ae6bb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h11d63595ef29da3a13b39df22850769cca7082fee28015a93f6c9dea6764ababd6b0a5288f982d37d2c0425c8271c7c259420ddb0483eaf97ae0d784782e41f67b0670ea383eae6588efbb354bb63;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h150df156f10332921352530ae5e9e867170b88ad1c0555f3b3a3498fa99521cabc8907396f4666c459f35f4efc8908bfe596fd064f4abb5268d99d4a98680bf141097c281ea53b3bf6c3aa06d03ba;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fd468094dd601d20e31e954bbfcdb147b91b6e5bdaafc9151665ad1af10a29fca3de9774b05ce89944f00d263d0b3acd9158b1e597a97f75aa2a0d0974752a4aa06ed1f1b9d851e3525b58097170;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h16aa9635b62a973551692495c312679e1063439e320fbef98c8429e7cd64a37f7385863dd34f0b578b2e779713525de79adf83e6259cb5c4334652c06b2ea4669c1490619fcaca6a49bf07a12044d;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1f1cb77c5e91eeeea8046e9921b41f1b8f4f7fc5dd7ef2f68c29df9c3f12df14c3b50f0ad7a5f8d37135e7ec41d2b6bf539ec63417f29ca4bd58fddc17c2fc484a9561d5ee71250c3f23178cd8b80;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1dff1349fb875a91ddcdccc7ce14c6326d16e9d4faa18a9636f76ffde5afbe77560bdda905c4d5a7251b5f825ad934d067b11d7f0576b793f93cc28d93dd5b51d5a9258b5a815bade3d90df638d2c;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h688b08475e957cfad1a57394334eab25a3b2d4b4bc76e3bb0bb9439a8db6f8565948d4b1c574dd91a21dfd6c85671ae3734aae9a7d34b05621a5d76267247d1378829d5f43e5dae105dda73fc8b2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1504b9ddc5b8f4a21493cb24fcf81a66f77493f31f81904a30bb1f0dc3274e28a3df5e4e388eaec822f9b0b8a8dda5b48478017bfea93ef02582db0e5d4c6632559a3cbd9f52ce1425a5b7c000232;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h283de753ff647c4f60c95c75095e11c077c541664e365914240576ca38dd131942d709627d5a969941afae8a01376d5bdaef27b27d0f027e5c263bb245026888752999c121151ae2956e6c2b5678;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1c670dd6bb47b74a0319f6a681137106c4132edfa871026a6e636b463bf1d6badce1fc6b3b7cb7aa33e6b213ac7efae04b7ad2a8d49566363c2cd06ff0f050ad1e37e5010322db0a3d1f394b0ced5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1266696ed3c82e35ae31848c007c6320ce20a9c1c2bce76b8462eab4c67b4a1b3c2b5eb274b6e6c7d7d27aac77c4cbc481e1e3c3241c39c9536d5f4216724da7f9f8a5dabab202b34f60f03b48e6e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15abb655b054e62cbc1bfb4b879271bda0f4417a2b50c1186d2e249efed7c198a7247cca30a6ccec8afdeafdaff518eafe7a9381b113358fce6bada0ca1bef96b70fb6e4fa23e5c2348ef1d27c5a4;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he231639d79da4e112cbe5e2bf60a0a1bfb667bff8688a8712302efa8a718559b64f52bf2679a379180785797de5ef38c08eb30d66f6cfb159905460899079601be33d393d4a2b12569395933dba2;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h119685da34bf9b8ce8fd5e8191613ff7d80e1b2a36474d0bfca666fc06cf715b6895fc256754339b04b68124345fefa7cd4bcba57fbc3413bae528ef556754a49d2553959ab458c8137f3ae07cc86;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fb0a505088911c8f5c3da0fc0b39f3ba7cdd5b488cc83c75a130dda48e011a16083ba2ec741ab30011649a1a999a711fb967683ee7f18e015f6328a6a293a185ac6fbbd8b29cfd689e48c3aca833;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he7709c866ab366d58e7657a79c794471ab6a43c21f33d50215a69481dfe8ab2a547d7547bd7c5bff1ba8b629f7a07e3967df4870c08bf6eaeba178a964be44d2fe6065a6aeaebc5499266157266a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'he1398cad3e28c046fd75ab8b2ef788fbc75757b815edd363f47c89d312817a6eeb3ebe2b223965bff09f6a2de9070c87ffb231be8119afadf24450901ea90d7b4d2f2fdc85b7c785b8f2d8647c15;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1de51e985f8993285666e770899ddaed64c68e0c5a61f8dce9345324b47ef5f71cc849e6bd32dc505e4754d38c67fef072d1733c865996ee2d701e2d6c34e4e4f61c16cfadaad8475a081c30285c9;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h15d3f4f2d40abdf5c5a38524b40787f6496f26954fda0f93b8554d8aacab500a72e926863d103a47ae03fc97b1188b8269e57d0b11d9a2e9b2bf96ed8f7cc399ebcb74be9b9e47402d0c1371f6573;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h968bb60ef212bdefa72aa728adecf42bd739ccbc947d4d48b6671ccb4bcfee889d8f73f1bd706c5cc98f333dc21cdbcb08dd30d07d2b6d94776ee7c8435a5f73a5e1422c68e633fc42417e45c530;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd7b2c28a7d7abb0f131d4828c2d81ed13bd992219ef50ed262ee94ce9f29f3096651b2eea4b340ea44fa418726e32c70556e1d231f74cdc5e03a7bb469dc0c02d227cee5a450eb22ea7ac5ca71e6;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h3f65a4b43e9556c706a39435035a9063ab9012f270d46c1b560a3e34c5acc0cc614ba3aa6590715543a7c4fd88066e1c110a446e019c69fadf9bfdabb087d49814077d56c4b47ba744e1fdc89c5b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1d34cf0c6111593d5b507c34af51e3f3993b8d8780c6a56c42eeaf32a4173f51608dbe8ee95cab1d809be4daa656b12b1b840ce073a80d14d86b1bd0692e4ef06b488b9422376f351c450a4d73121;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h567295e8f7ebc6893ad3abad3b1c1bf1bee8e0319e0225d8c7b49acfa9cd9945173fc973a70a4dab49574dd778a4da172de62ea726419359a9536c5c2ceef5ab6879dfcafb006a6fc421eec7122;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hdccd5ab0c48bfdaa981f29ee78bc3599f20cd8b9a8e10c97eed2676922cf884630e2c00534d75712c9030df16c955ebeb82ee36f43c256aaa8d75d4c05d8829a88b98a0fc842ce791b334e6db6a5;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h2a9532f47e4ec0b4822feabc0ac74ed86bd6e7e7833c02db9ddadf259f581fc504ba025bf81f715b1040f24e34fd0fe034994abdb26866a6ddd4ae37ed3d482704e7562ac53b94c0d5fd59b8475e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h9bf6cc3325931df1b57d6cabea6746833ae87e590665d904122e7ea86a3870f540a2938174f499dee99c36f412c6dac90a5821581ffe292c83d75bf6f77baea5651786e3de378c3fc4a4f56db7d7;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h389ffea082e7ae37dc9b4d4c3421c368285447302a28d17bd26db33f9f3eb810273d740d2a415c5f0001e5e2ebdc73e467124ecfb65ad11863c9cea341187f0e333782cf9ee3e2e35b3b135e487a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h133a4c067cc12ee5c17d9eb40cca2023ce0837d6f7fd41da3b04d7e691ec1300c0dcf68af3cfb5fd38808a31688404c248d9a508d565215a5a28268329668ca113f16b5a600f5d2a8f4b50d1bf50e;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1cb265dc0dc133bcf43a8ec8cccfbbc969131064284cea42b7403f619f729c071ed50d3b506621bdfef49369c56f2c3e8ed19c6fe640f4f6bca07c3cbf9177530a52148cb0eb9f50fec5d088db82a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hd38b3e10863b15400851ce6bf6de4a954ab8b7d1fc4e1cd9b8a1f2f7703809b78952bc2516271a8d18601ad286271f4487ae0a40139877edb090c54683bb165f41a418b1030af463f1ae9e608aaa;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1fed44521019ac9d1423c01d967bd0c99f35e7ca987032b618d221837a7a57530eeaeb94d98448a8e1e70153a48ab5e921e49a7ad2d5fee18c9331fd31430514e50134b5f682a102f002bdf9c5055;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h10eda82c741eeba8a1512d85e6648350873dbfffef5b5e7bf22a8961edf17ddc9ec7d5fc732cac4ef94f404060a9201941b25669b3969240093cd603b9dc7bd4124c43d401cd637c0cfaa9e50ddfb;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7c88e47d3b4cb2dfe7a34bb567cfdff431d90ce110c6287e94c9810a812ceeba56123f069a717e842f1ceec209e66443f81fcc6efc41b60e1fa016118bfc1788cdc31f46bf094c7088dc531afcd;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1788c53b01c8b4d0471fe5a1cca2a95bcef7511ed4c71246d86b2bab5cc4ac358a7603ec2c4d2ad2ba89bc15bd8b330bb8bc6523c760867e8d908ba66c51b42e0f2f941e20925ebaf7dc7d784e327;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h88c32c53f214b702f49080af8f8c8f53faca1b21fa77449d442b4b30a5c704e2dd5a8b395544ae307afdb8e17beb6221372b17635d2712da93d6b00df24d31d8223b35e4b0baa9076c2a2a8a052b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1e82f966db02e385beaea4dd264d1828a2174d82d46367ee48917506580c91f12d00c362a7836d1dd18b983531cf88e02a7c029c2e8728a669e84eeea7bb539e86edea119930a8dd3e7efd075226a;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h5920794cda0f4da7517664b49e052bd5a857fd2060a9ff23588d57399f82f22e33007ae645735ecdb32b93bba529f5475a49dbb5afd35affaf7fd32803e2a30ba982cdcb375da8016ad444e27a21;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h1ce1655dae65d0551e73a57b1d2494924e35e49056da78ce4052e9fbfd34bba82857a2564450b105aab4d81abde26970e0d47cffb0c8d008cf4b2d674572e7f47dbd84530b8242cf45a48cdb9fb74;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hc47d19cfad38e80c151709db24e4679a5b4eeb3ad067a5ccfa7feaedfb6156f429718de8b0bdec535b3eb95f889742227a3acba78467527445f46fa69ce5bb0c2ac63d8df2085cb6a5d0381ada67;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h7f339bbe1c24e79e491ac66b8543d40b9447a004f6cdcef9e789f54bd7672b2065c830063a22321cdca462c95aa47a9242639b23b7e029bbec03afde28e9aa2458e514a98526cab741434f0bd05b;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'h189a59494a55d53498fcd8a1e2245c45e6063b6645beb6464a15f40146479b9130bdbedd05520be4b7d1fef002fb94d759b48afe9068cfe7e8392cc7bae885b8ad25c72ab918487b0dd8518622177;
        #1
        {src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 625'hb41bcdf4d39d0b88d07ea2c87604b673cf03fd0ad55791066b1e7a5a455190dadac1da0bfd513c2cf7dea3da57aa1446406c737c72a2db2941caa4f0117060585cbfdf457eb02883e2ecd41d2d08;
        #1
        $finish();
    end
endmodule
