module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69);
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    reg [53:0] src12;
    reg [53:0] src13;
    reg [53:0] src14;
    reg [53:0] src15;
    reg [53:0] src16;
    reg [53:0] src17;
    reg [53:0] src18;
    reg [53:0] src19;
    reg [53:0] src20;
    reg [53:0] src21;
    reg [53:0] src22;
    reg [53:0] src23;
    reg [53:0] src24;
    reg [53:0] src25;
    reg [53:0] src26;
    reg [53:0] src27;
    reg [53:0] src28;
    reg [53:0] src29;
    reg [53:0] src30;
    reg [53:0] src31;
    reg [53:0] src32;
    reg [53:0] src33;
    reg [53:0] src34;
    reg [53:0] src35;
    reg [53:0] src36;
    reg [53:0] src37;
    reg [53:0] src38;
    reg [53:0] src39;
    reg [53:0] src40;
    reg [53:0] src41;
    reg [53:0] src42;
    reg [53:0] src43;
    reg [53:0] src44;
    reg [53:0] src45;
    reg [53:0] src46;
    reg [53:0] src47;
    reg [53:0] src48;
    reg [53:0] src49;
    reg [53:0] src50;
    reg [53:0] src51;
    reg [53:0] src52;
    reg [53:0] src53;
    reg [53:0] src54;
    reg [53:0] src55;
    reg [53:0] src56;
    reg [53:0] src57;
    reg [53:0] src58;
    reg [53:0] src59;
    reg [53:0] src60;
    reg [53:0] src61;
    reg [53:0] src62;
    reg [53:0] src63;
    compressor_CLA54_64 compressor_CLA54_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69));
    initial begin
        src0 <= 54'h0;
        src1 <= 54'h0;
        src2 <= 54'h0;
        src3 <= 54'h0;
        src4 <= 54'h0;
        src5 <= 54'h0;
        src6 <= 54'h0;
        src7 <= 54'h0;
        src8 <= 54'h0;
        src9 <= 54'h0;
        src10 <= 54'h0;
        src11 <= 54'h0;
        src12 <= 54'h0;
        src13 <= 54'h0;
        src14 <= 54'h0;
        src15 <= 54'h0;
        src16 <= 54'h0;
        src17 <= 54'h0;
        src18 <= 54'h0;
        src19 <= 54'h0;
        src20 <= 54'h0;
        src21 <= 54'h0;
        src22 <= 54'h0;
        src23 <= 54'h0;
        src24 <= 54'h0;
        src25 <= 54'h0;
        src26 <= 54'h0;
        src27 <= 54'h0;
        src28 <= 54'h0;
        src29 <= 54'h0;
        src30 <= 54'h0;
        src31 <= 54'h0;
        src32 <= 54'h0;
        src33 <= 54'h0;
        src34 <= 54'h0;
        src35 <= 54'h0;
        src36 <= 54'h0;
        src37 <= 54'h0;
        src38 <= 54'h0;
        src39 <= 54'h0;
        src40 <= 54'h0;
        src41 <= 54'h0;
        src42 <= 54'h0;
        src43 <= 54'h0;
        src44 <= 54'h0;
        src45 <= 54'h0;
        src46 <= 54'h0;
        src47 <= 54'h0;
        src48 <= 54'h0;
        src49 <= 54'h0;
        src50 <= 54'h0;
        src51 <= 54'h0;
        src52 <= 54'h0;
        src53 <= 54'h0;
        src54 <= 54'h0;
        src55 <= 54'h0;
        src56 <= 54'h0;
        src57 <= 54'h0;
        src58 <= 54'h0;
        src59 <= 54'h0;
        src60 <= 54'h0;
        src61 <= 54'h0;
        src62 <= 54'h0;
        src63 <= 54'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor_CLA54_64(
    input [53:0]src0,
    input [53:0]src1,
    input [53:0]src2,
    input [53:0]src3,
    input [53:0]src4,
    input [53:0]src5,
    input [53:0]src6,
    input [53:0]src7,
    input [53:0]src8,
    input [53:0]src9,
    input [53:0]src10,
    input [53:0]src11,
    input [53:0]src12,
    input [53:0]src13,
    input [53:0]src14,
    input [53:0]src15,
    input [53:0]src16,
    input [53:0]src17,
    input [53:0]src18,
    input [53:0]src19,
    input [53:0]src20,
    input [53:0]src21,
    input [53:0]src22,
    input [53:0]src23,
    input [53:0]src24,
    input [53:0]src25,
    input [53:0]src26,
    input [53:0]src27,
    input [53:0]src28,
    input [53:0]src29,
    input [53:0]src30,
    input [53:0]src31,
    input [53:0]src32,
    input [53:0]src33,
    input [53:0]src34,
    input [53:0]src35,
    input [53:0]src36,
    input [53:0]src37,
    input [53:0]src38,
    input [53:0]src39,
    input [53:0]src40,
    input [53:0]src41,
    input [53:0]src42,
    input [53:0]src43,
    input [53:0]src44,
    input [53:0]src45,
    input [53:0]src46,
    input [53:0]src47,
    input [53:0]src48,
    input [53:0]src49,
    input [53:0]src50,
    input [53:0]src51,
    input [53:0]src52,
    input [53:0]src53,
    input [53:0]src54,
    input [53:0]src55,
    input [53:0]src56,
    input [53:0]src57,
    input [53:0]src58,
    input [53:0]src59,
    input [53:0]src60,
    input [53:0]src61,
    input [53:0]src62,
    input [53:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [0:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [0:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [1:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [1:0] comp_out67;
    wire [0:0] comp_out68;
    wire [0:0] comp_out69;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69)
    );
    LookAheadCarryUnit256 LCU256(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out67[1], comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], comp_out62[1], comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], 1'h0, comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], 1'h0, comp_out3[1], 1'h0, comp_out1[1], comp_out0[1]}),
        .dst({dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [53:0] src0,
      input wire [53:0] src1,
      input wire [53:0] src2,
      input wire [53:0] src3,
      input wire [53:0] src4,
      input wire [53:0] src5,
      input wire [53:0] src6,
      input wire [53:0] src7,
      input wire [53:0] src8,
      input wire [53:0] src9,
      input wire [53:0] src10,
      input wire [53:0] src11,
      input wire [53:0] src12,
      input wire [53:0] src13,
      input wire [53:0] src14,
      input wire [53:0] src15,
      input wire [53:0] src16,
      input wire [53:0] src17,
      input wire [53:0] src18,
      input wire [53:0] src19,
      input wire [53:0] src20,
      input wire [53:0] src21,
      input wire [53:0] src22,
      input wire [53:0] src23,
      input wire [53:0] src24,
      input wire [53:0] src25,
      input wire [53:0] src26,
      input wire [53:0] src27,
      input wire [53:0] src28,
      input wire [53:0] src29,
      input wire [53:0] src30,
      input wire [53:0] src31,
      input wire [53:0] src32,
      input wire [53:0] src33,
      input wire [53:0] src34,
      input wire [53:0] src35,
      input wire [53:0] src36,
      input wire [53:0] src37,
      input wire [53:0] src38,
      input wire [53:0] src39,
      input wire [53:0] src40,
      input wire [53:0] src41,
      input wire [53:0] src42,
      input wire [53:0] src43,
      input wire [53:0] src44,
      input wire [53:0] src45,
      input wire [53:0] src46,
      input wire [53:0] src47,
      input wire [53:0] src48,
      input wire [53:0] src49,
      input wire [53:0] src50,
      input wire [53:0] src51,
      input wire [53:0] src52,
      input wire [53:0] src53,
      input wire [53:0] src54,
      input wire [53:0] src55,
      input wire [53:0] src56,
      input wire [53:0] src57,
      input wire [53:0] src58,
      input wire [53:0] src59,
      input wire [53:0] src60,
      input wire [53:0] src61,
      input wire [53:0] src62,
      input wire [53:0] src63,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [0:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [0:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [0:0] dst68,
      output wire [0:0] dst69);

   wire [53:0] stage0_0;
   wire [53:0] stage0_1;
   wire [53:0] stage0_2;
   wire [53:0] stage0_3;
   wire [53:0] stage0_4;
   wire [53:0] stage0_5;
   wire [53:0] stage0_6;
   wire [53:0] stage0_7;
   wire [53:0] stage0_8;
   wire [53:0] stage0_9;
   wire [53:0] stage0_10;
   wire [53:0] stage0_11;
   wire [53:0] stage0_12;
   wire [53:0] stage0_13;
   wire [53:0] stage0_14;
   wire [53:0] stage0_15;
   wire [53:0] stage0_16;
   wire [53:0] stage0_17;
   wire [53:0] stage0_18;
   wire [53:0] stage0_19;
   wire [53:0] stage0_20;
   wire [53:0] stage0_21;
   wire [53:0] stage0_22;
   wire [53:0] stage0_23;
   wire [53:0] stage0_24;
   wire [53:0] stage0_25;
   wire [53:0] stage0_26;
   wire [53:0] stage0_27;
   wire [53:0] stage0_28;
   wire [53:0] stage0_29;
   wire [53:0] stage0_30;
   wire [53:0] stage0_31;
   wire [53:0] stage0_32;
   wire [53:0] stage0_33;
   wire [53:0] stage0_34;
   wire [53:0] stage0_35;
   wire [53:0] stage0_36;
   wire [53:0] stage0_37;
   wire [53:0] stage0_38;
   wire [53:0] stage0_39;
   wire [53:0] stage0_40;
   wire [53:0] stage0_41;
   wire [53:0] stage0_42;
   wire [53:0] stage0_43;
   wire [53:0] stage0_44;
   wire [53:0] stage0_45;
   wire [53:0] stage0_46;
   wire [53:0] stage0_47;
   wire [53:0] stage0_48;
   wire [53:0] stage0_49;
   wire [53:0] stage0_50;
   wire [53:0] stage0_51;
   wire [53:0] stage0_52;
   wire [53:0] stage0_53;
   wire [53:0] stage0_54;
   wire [53:0] stage0_55;
   wire [53:0] stage0_56;
   wire [53:0] stage0_57;
   wire [53:0] stage0_58;
   wire [53:0] stage0_59;
   wire [53:0] stage0_60;
   wire [53:0] stage0_61;
   wire [53:0] stage0_62;
   wire [53:0] stage0_63;
   wire [16:0] stage1_0;
   wire [19:0] stage1_1;
   wire [24:0] stage1_2;
   wire [23:0] stage1_3;
   wire [32:0] stage1_4;
   wire [35:0] stage1_5;
   wire [18:0] stage1_6;
   wire [24:0] stage1_7;
   wire [30:0] stage1_8;
   wire [17:0] stage1_9;
   wire [25:0] stage1_10;
   wire [28:0] stage1_11;
   wire [20:0] stage1_12;
   wire [29:0] stage1_13;
   wire [23:0] stage1_14;
   wire [42:0] stage1_15;
   wire [23:0] stage1_16;
   wire [17:0] stage1_17;
   wire [33:0] stage1_18;
   wire [20:0] stage1_19;
   wire [19:0] stage1_20;
   wire [25:0] stage1_21;
   wire [22:0] stage1_22;
   wire [21:0] stage1_23;
   wire [31:0] stage1_24;
   wire [24:0] stage1_25;
   wire [31:0] stage1_26;
   wire [23:0] stage1_27;
   wire [17:0] stage1_28;
   wire [25:0] stage1_29;
   wire [34:0] stage1_30;
   wire [33:0] stage1_31;
   wire [18:0] stage1_32;
   wire [45:0] stage1_33;
   wire [18:0] stage1_34;
   wire [27:0] stage1_35;
   wire [33:0] stage1_36;
   wire [24:0] stage1_37;
   wire [23:0] stage1_38;
   wire [30:0] stage1_39;
   wire [38:0] stage1_40;
   wire [19:0] stage1_41;
   wire [20:0] stage1_42;
   wire [22:0] stage1_43;
   wire [21:0] stage1_44;
   wire [31:0] stage1_45;
   wire [29:0] stage1_46;
   wire [33:0] stage1_47;
   wire [17:0] stage1_48;
   wire [23:0] stage1_49;
   wire [42:0] stage1_50;
   wire [47:0] stage1_51;
   wire [21:0] stage1_52;
   wire [40:0] stage1_53;
   wire [16:0] stage1_54;
   wire [37:0] stage1_55;
   wire [20:0] stage1_56;
   wire [40:0] stage1_57;
   wire [14:0] stage1_58;
   wire [34:0] stage1_59;
   wire [22:0] stage1_60;
   wire [20:0] stage1_61;
   wire [23:0] stage1_62;
   wire [34:0] stage1_63;
   wire [13:0] stage1_64;
   wire [5:0] stage1_65;
   wire [5:0] stage2_0;
   wire [6:0] stage2_1;
   wire [13:0] stage2_2;
   wire [8:0] stage2_3;
   wire [22:0] stage2_4;
   wire [9:0] stage2_5;
   wire [10:0] stage2_6;
   wire [12:0] stage2_7;
   wire [10:0] stage2_8;
   wire [19:0] stage2_9;
   wire [9:0] stage2_10;
   wire [12:0] stage2_11;
   wire [9:0] stage2_12;
   wire [9:0] stage2_13;
   wire [14:0] stage2_14;
   wire [13:0] stage2_15;
   wire [10:0] stage2_16;
   wire [11:0] stage2_17;
   wire [19:0] stage2_18;
   wire [8:0] stage2_19;
   wire [8:0] stage2_20;
   wire [21:0] stage2_21;
   wire [10:0] stage2_22;
   wire [20:0] stage2_23;
   wire [9:0] stage2_24;
   wire [12:0] stage2_25;
   wire [18:0] stage2_26;
   wire [6:0] stage2_27;
   wire [13:0] stage2_28;
   wire [17:0] stage2_29;
   wire [9:0] stage2_30;
   wire [16:0] stage2_31;
   wire [11:0] stage2_32;
   wire [15:0] stage2_33;
   wire [15:0] stage2_34;
   wire [10:0] stage2_35;
   wire [18:0] stage2_36;
   wire [16:0] stage2_37;
   wire [12:0] stage2_38;
   wire [16:0] stage2_39;
   wire [11:0] stage2_40;
   wire [12:0] stage2_41;
   wire [13:0] stage2_42;
   wire [9:0] stage2_43;
   wire [14:0] stage2_44;
   wire [11:0] stage2_45;
   wire [17:0] stage2_46;
   wire [21:0] stage2_47;
   wire [12:0] stage2_48;
   wire [17:0] stage2_49;
   wire [10:0] stage2_50;
   wire [16:0] stage2_51;
   wire [18:0] stage2_52;
   wire [12:0] stage2_53;
   wire [14:0] stage2_54;
   wire [18:0] stage2_55;
   wire [12:0] stage2_56;
   wire [12:0] stage2_57;
   wire [17:0] stage2_58;
   wire [12:0] stage2_59;
   wire [12:0] stage2_60;
   wire [11:0] stage2_61;
   wire [17:0] stage2_62;
   wire [16:0] stage2_63;
   wire [5:0] stage2_64;
   wire [9:0] stage2_65;
   wire [3:0] stage2_66;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [4:0] stage3_2;
   wire [5:0] stage3_3;
   wire [14:0] stage3_4;
   wire [8:0] stage3_5;
   wire [4:0] stage3_6;
   wire [13:0] stage3_7;
   wire [6:0] stage3_8;
   wire [10:0] stage3_9;
   wire [6:0] stage3_10;
   wire [3:0] stage3_11;
   wire [4:0] stage3_12;
   wire [7:0] stage3_13;
   wire [3:0] stage3_14;
   wire [5:0] stage3_15;
   wire [5:0] stage3_16;
   wire [7:0] stage3_17;
   wire [5:0] stage3_18;
   wire [7:0] stage3_19;
   wire [4:0] stage3_20;
   wire [6:0] stage3_21;
   wire [6:0] stage3_22;
   wire [4:0] stage3_23;
   wire [5:0] stage3_24;
   wire [7:0] stage3_25;
   wire [5:0] stage3_26;
   wire [4:0] stage3_27;
   wire [4:0] stage3_28;
   wire [11:0] stage3_29;
   wire [5:0] stage3_30;
   wire [6:0] stage3_31;
   wire [3:0] stage3_32;
   wire [14:0] stage3_33;
   wire [8:0] stage3_34;
   wire [3:0] stage3_35;
   wire [5:0] stage3_36;
   wire [6:0] stage3_37;
   wire [6:0] stage3_38;
   wire [5:0] stage3_39;
   wire [6:0] stage3_40;
   wire [6:0] stage3_41;
   wire [5:0] stage3_42;
   wire [7:0] stage3_43;
   wire [7:0] stage3_44;
   wire [4:0] stage3_45;
   wire [5:0] stage3_46;
   wire [8:0] stage3_47;
   wire [12:0] stage3_48;
   wire [5:0] stage3_49;
   wire [10:0] stage3_50;
   wire [7:0] stage3_51;
   wire [10:0] stage3_52;
   wire [6:0] stage3_53;
   wire [5:0] stage3_54;
   wire [5:0] stage3_55;
   wire [10:0] stage3_56;
   wire [7:0] stage3_57;
   wire [3:0] stage3_58;
   wire [13:0] stage3_59;
   wire [5:0] stage3_60;
   wire [9:0] stage3_61;
   wire [3:0] stage3_62;
   wire [9:0] stage3_63;
   wire [4:0] stage3_64;
   wire [6:0] stage3_65;
   wire [5:0] stage3_66;
   wire [0:0] stage3_67;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [0:0] stage4_2;
   wire [1:0] stage4_3;
   wire [5:0] stage4_4;
   wire [2:0] stage4_5;
   wire [3:0] stage4_6;
   wire [5:0] stage4_7;
   wire [3:0] stage4_8;
   wire [2:0] stage4_9;
   wire [3:0] stage4_10;
   wire [3:0] stage4_11;
   wire [3:0] stage4_12;
   wire [1:0] stage4_13;
   wire [2:0] stage4_14;
   wire [4:0] stage4_15;
   wire [3:0] stage4_16;
   wire [1:0] stage4_17;
   wire [6:0] stage4_18;
   wire [2:0] stage4_19;
   wire [2:0] stage4_20;
   wire [3:0] stage4_21;
   wire [1:0] stage4_22;
   wire [2:0] stage4_23;
   wire [2:0] stage4_24;
   wire [2:0] stage4_25;
   wire [3:0] stage4_26;
   wire [5:0] stage4_27;
   wire [0:0] stage4_28;
   wire [5:0] stage4_29;
   wire [2:0] stage4_30;
   wire [1:0] stage4_31;
   wire [2:0] stage4_32;
   wire [5:0] stage4_33;
   wire [2:0] stage4_34;
   wire [3:0] stage4_35;
   wire [2:0] stage4_36;
   wire [5:0] stage4_37;
   wire [6:0] stage4_38;
   wire [0:0] stage4_39;
   wire [2:0] stage4_40;
   wire [2:0] stage4_41;
   wire [2:0] stage4_42;
   wire [3:0] stage4_43;
   wire [5:0] stage4_44;
   wire [1:0] stage4_45;
   wire [2:0] stage4_46;
   wire [3:0] stage4_47;
   wire [3:0] stage4_48;
   wire [2:0] stage4_49;
   wire [3:0] stage4_50;
   wire [4:0] stage4_51;
   wire [3:0] stage4_52;
   wire [2:0] stage4_53;
   wire [2:0] stage4_54;
   wire [3:0] stage4_55;
   wire [5:0] stage4_56;
   wire [2:0] stage4_57;
   wire [2:0] stage4_58;
   wire [5:0] stage4_59;
   wire [2:0] stage4_60;
   wire [5:0] stage4_61;
   wire [2:0] stage4_62;
   wire [5:0] stage4_63;
   wire [2:0] stage4_64;
   wire [2:0] stage4_65;
   wire [2:0] stage4_66;
   wire [2:0] stage4_67;
   wire [0:0] stage4_68;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [0:0] stage5_2;
   wire [1:0] stage5_3;
   wire [0:0] stage5_4;
   wire [1:0] stage5_5;
   wire [1:0] stage5_6;
   wire [1:0] stage5_7;
   wire [1:0] stage5_8;
   wire [1:0] stage5_9;
   wire [1:0] stage5_10;
   wire [1:0] stage5_11;
   wire [1:0] stage5_12;
   wire [1:0] stage5_13;
   wire [1:0] stage5_14;
   wire [1:0] stage5_15;
   wire [1:0] stage5_16;
   wire [1:0] stage5_17;
   wire [1:0] stage5_18;
   wire [1:0] stage5_19;
   wire [1:0] stage5_20;
   wire [1:0] stage5_21;
   wire [1:0] stage5_22;
   wire [1:0] stage5_23;
   wire [1:0] stage5_24;
   wire [1:0] stage5_25;
   wire [1:0] stage5_26;
   wire [1:0] stage5_27;
   wire [1:0] stage5_28;
   wire [0:0] stage5_29;
   wire [1:0] stage5_30;
   wire [1:0] stage5_31;
   wire [1:0] stage5_32;
   wire [1:0] stage5_33;
   wire [1:0] stage5_34;
   wire [1:0] stage5_35;
   wire [1:0] stage5_36;
   wire [1:0] stage5_37;
   wire [1:0] stage5_38;
   wire [1:0] stage5_39;
   wire [1:0] stage5_40;
   wire [1:0] stage5_41;
   wire [1:0] stage5_42;
   wire [1:0] stage5_43;
   wire [1:0] stage5_44;
   wire [1:0] stage5_45;
   wire [1:0] stage5_46;
   wire [1:0] stage5_47;
   wire [1:0] stage5_48;
   wire [1:0] stage5_49;
   wire [1:0] stage5_50;
   wire [1:0] stage5_51;
   wire [1:0] stage5_52;
   wire [1:0] stage5_53;
   wire [1:0] stage5_54;
   wire [1:0] stage5_55;
   wire [1:0] stage5_56;
   wire [1:0] stage5_57;
   wire [1:0] stage5_58;
   wire [1:0] stage5_59;
   wire [1:0] stage5_60;
   wire [1:0] stage5_61;
   wire [1:0] stage5_62;
   wire [1:0] stage5_63;
   wire [1:0] stage5_64;
   wire [1:0] stage5_65;
   wire [1:0] stage5_66;
   wire [1:0] stage5_67;
   wire [0:0] stage5_68;
   wire [0:0] stage5_69;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage5_0;
   assign dst1 = stage5_1;
   assign dst2 = stage5_2;
   assign dst3 = stage5_3;
   assign dst4 = stage5_4;
   assign dst5 = stage5_5;
   assign dst6 = stage5_6;
   assign dst7 = stage5_7;
   assign dst8 = stage5_8;
   assign dst9 = stage5_9;
   assign dst10 = stage5_10;
   assign dst11 = stage5_11;
   assign dst12 = stage5_12;
   assign dst13 = stage5_13;
   assign dst14 = stage5_14;
   assign dst15 = stage5_15;
   assign dst16 = stage5_16;
   assign dst17 = stage5_17;
   assign dst18 = stage5_18;
   assign dst19 = stage5_19;
   assign dst20 = stage5_20;
   assign dst21 = stage5_21;
   assign dst22 = stage5_22;
   assign dst23 = stage5_23;
   assign dst24 = stage5_24;
   assign dst25 = stage5_25;
   assign dst26 = stage5_26;
   assign dst27 = stage5_27;
   assign dst28 = stage5_28;
   assign dst29 = stage5_29;
   assign dst30 = stage5_30;
   assign dst31 = stage5_31;
   assign dst32 = stage5_32;
   assign dst33 = stage5_33;
   assign dst34 = stage5_34;
   assign dst35 = stage5_35;
   assign dst36 = stage5_36;
   assign dst37 = stage5_37;
   assign dst38 = stage5_38;
   assign dst39 = stage5_39;
   assign dst40 = stage5_40;
   assign dst41 = stage5_41;
   assign dst42 = stage5_42;
   assign dst43 = stage5_43;
   assign dst44 = stage5_44;
   assign dst45 = stage5_45;
   assign dst46 = stage5_46;
   assign dst47 = stage5_47;
   assign dst48 = stage5_48;
   assign dst49 = stage5_49;
   assign dst50 = stage5_50;
   assign dst51 = stage5_51;
   assign dst52 = stage5_52;
   assign dst53 = stage5_53;
   assign dst54 = stage5_54;
   assign dst55 = stage5_55;
   assign dst56 = stage5_56;
   assign dst57 = stage5_57;
   assign dst58 = stage5_58;
   assign dst59 = stage5_59;
   assign dst60 = stage5_60;
   assign dst61 = stage5_61;
   assign dst62 = stage5_62;
   assign dst63 = stage5_63;
   assign dst64 = stage5_64;
   assign dst65 = stage5_65;
   assign dst66 = stage5_66;
   assign dst67 = stage5_67;
   assign dst68 = stage5_68;
   assign dst69 = stage5_69;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1163_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[1]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[2]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc7_3 gpc3 (
      {stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14], stage0_0[15]},
      {stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc606_5 gpc4 (
      {stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20], stage0_0[21]},
      {stage0_2[3], stage0_2[4], stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8]},
      {stage1_4[3],stage1_3[3],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27]},
      {stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14]},
      {stage1_4[4],stage1_3[4],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33]},
      {stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19], stage0_2[20]},
      {stage1_4[5],stage1_3[5],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc606_5 gpc7 (
      {stage0_0[34], stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25], stage0_2[26]},
      {stage1_4[6],stage1_3[6],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45]},
      {stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31], stage0_2[32]},
      {stage1_4[7],stage1_3[7],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_3[3], stage0_3[4], stage0_3[5], stage0_3[6], stage0_3[7], stage0_3[8]},
      {stage1_5[0],stage1_4[8],stage1_3[8],stage1_2[9],stage1_1[9]}
   );
   gpc606_5 gpc10 (
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13], stage0_3[14]},
      {stage1_5[1],stage1_4[9],stage1_3[9],stage1_2[10],stage1_1[10]}
   );
   gpc606_5 gpc11 (
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19], stage0_3[20]},
      {stage1_5[2],stage1_4[10],stage1_3[10],stage1_2[11],stage1_1[11]}
   );
   gpc606_5 gpc12 (
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26]},
      {stage1_5[3],stage1_4[11],stage1_3[11],stage1_2[12],stage1_1[12]}
   );
   gpc606_5 gpc13 (
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32]},
      {stage1_5[4],stage1_4[12],stage1_3[12],stage1_2[13],stage1_1[13]}
   );
   gpc606_5 gpc14 (
      {stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37], stage0_2[38]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[5],stage1_4[13],stage1_3[13],stage1_2[14]}
   );
   gpc606_5 gpc15 (
      {stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43], stage0_2[44]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[6],stage1_4[14],stage1_3[14],stage1_2[15]}
   );
   gpc615_5 gpc16 (
      {stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37]},
      {stage0_4[12]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[2],stage1_5[7],stage1_4[15],stage1_3[15]}
   );
   gpc615_5 gpc17 (
      {stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42]},
      {stage0_4[13]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[3],stage1_5[8],stage1_4[16],stage1_3[16]}
   );
   gpc615_5 gpc18 (
      {stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47]},
      {stage0_4[14]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[4],stage1_5[9],stage1_4[17],stage1_3[17]}
   );
   gpc615_5 gpc19 (
      {stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18], stage0_4[19]},
      {stage0_5[18]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[3],stage1_6[5],stage1_5[10],stage1_4[18]}
   );
   gpc615_5 gpc20 (
      {stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24]},
      {stage0_5[19]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[4],stage1_6[6],stage1_5[11],stage1_4[19]}
   );
   gpc615_5 gpc21 (
      {stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage0_5[20]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[5],stage1_6[7],stage1_5[12],stage1_4[20]}
   );
   gpc615_5 gpc22 (
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34]},
      {stage0_5[21]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[6],stage1_6[8],stage1_5[13],stage1_4[21]}
   );
   gpc615_5 gpc23 (
      {stage0_4[35], stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39]},
      {stage0_5[22]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[7],stage1_6[9],stage1_5[14],stage1_4[22]}
   );
   gpc615_5 gpc24 (
      {stage0_4[40], stage0_4[41], stage0_4[42], stage0_4[43], stage0_4[44]},
      {stage0_5[23]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[8],stage1_6[10],stage1_5[15],stage1_4[23]}
   );
   gpc606_5 gpc25 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[6],stage1_7[9],stage1_6[11],stage1_5[16]}
   );
   gpc606_5 gpc26 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[7],stage1_7[10],stage1_6[12],stage1_5[17]}
   );
   gpc615_5 gpc27 (
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40]},
      {stage0_7[12]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[2],stage1_8[8],stage1_7[11],stage1_6[13]}
   );
   gpc615_5 gpc28 (
      {stage0_6[41], stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45]},
      {stage0_7[13]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[3],stage1_8[9],stage1_7[12],stage1_6[14]}
   );
   gpc615_5 gpc29 (
      {stage0_6[46], stage0_6[47], stage0_6[48], stage0_6[49], stage0_6[50]},
      {stage0_7[14]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[4],stage1_8[10],stage1_7[13],stage1_6[15]}
   );
   gpc606_5 gpc30 (
      {stage0_7[15], stage0_7[16], stage0_7[17], stage0_7[18], stage0_7[19], stage0_7[20]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[3],stage1_9[5],stage1_8[11],stage1_7[14]}
   );
   gpc606_5 gpc31 (
      {stage0_7[21], stage0_7[22], stage0_7[23], stage0_7[24], stage0_7[25], stage0_7[26]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[4],stage1_9[6],stage1_8[12],stage1_7[15]}
   );
   gpc606_5 gpc32 (
      {stage0_7[27], stage0_7[28], stage0_7[29], stage0_7[30], stage0_7[31], stage0_7[32]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[5],stage1_9[7],stage1_8[13],stage1_7[16]}
   );
   gpc606_5 gpc33 (
      {stage0_7[33], stage0_7[34], stage0_7[35], stage0_7[36], stage0_7[37], stage0_7[38]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[6],stage1_9[8],stage1_8[14],stage1_7[17]}
   );
   gpc615_5 gpc34 (
      {stage0_7[39], stage0_7[40], stage0_7[41], stage0_7[42], stage0_7[43]},
      {stage0_8[18]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[7],stage1_9[9],stage1_8[15],stage1_7[18]}
   );
   gpc615_5 gpc35 (
      {stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47], stage0_7[48]},
      {stage0_8[19]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[8],stage1_9[10],stage1_8[16],stage1_7[19]}
   );
   gpc606_5 gpc36 (
      {stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[6],stage1_10[9],stage1_9[11],stage1_8[17]}
   );
   gpc606_5 gpc37 (
      {stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[7],stage1_10[10],stage1_9[12],stage1_8[18]}
   );
   gpc606_5 gpc38 (
      {stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[8],stage1_10[11],stage1_9[13],stage1_8[19]}
   );
   gpc606_5 gpc39 (
      {stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[9],stage1_10[12],stage1_9[14],stage1_8[20]}
   );
   gpc606_5 gpc40 (
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[4],stage1_11[10],stage1_10[13],stage1_9[15]}
   );
   gpc606_5 gpc41 (
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[5],stage1_11[11],stage1_10[14],stage1_9[16]}
   );
   gpc606_5 gpc42 (
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[6],stage1_11[12],stage1_10[15],stage1_9[17]}
   );
   gpc615_5 gpc43 (
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28]},
      {stage0_11[18]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[3],stage1_12[7],stage1_11[13],stage1_10[16]}
   );
   gpc615_5 gpc44 (
      {stage0_10[29], stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33]},
      {stage0_11[19]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[4],stage1_12[8],stage1_11[14],stage1_10[17]}
   );
   gpc615_5 gpc45 (
      {stage0_10[34], stage0_10[35], stage0_10[36], stage0_10[37], stage0_10[38]},
      {stage0_11[20]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[5],stage1_12[9],stage1_11[15],stage1_10[18]}
   );
   gpc615_5 gpc46 (
      {stage0_10[39], stage0_10[40], stage0_10[41], stage0_10[42], stage0_10[43]},
      {stage0_11[21]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[6],stage1_12[10],stage1_11[16],stage1_10[19]}
   );
   gpc615_5 gpc47 (
      {stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47], stage0_10[48]},
      {stage0_11[22]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[7],stage1_12[11],stage1_11[17],stage1_10[20]}
   );
   gpc615_5 gpc48 (
      {stage0_11[23], stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27]},
      {stage0_12[30]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[5],stage1_13[8],stage1_12[12],stage1_11[18]}
   );
   gpc615_5 gpc49 (
      {stage0_11[28], stage0_11[29], stage0_11[30], stage0_11[31], stage0_11[32]},
      {stage0_12[31]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[6],stage1_13[9],stage1_12[13],stage1_11[19]}
   );
   gpc615_5 gpc50 (
      {stage0_11[33], stage0_11[34], stage0_11[35], stage0_11[36], stage0_11[37]},
      {stage0_12[32]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[7],stage1_13[10],stage1_12[14],stage1_11[20]}
   );
   gpc615_5 gpc51 (
      {stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41], stage0_11[42]},
      {stage0_12[33]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[8],stage1_13[11],stage1_12[15],stage1_11[21]}
   );
   gpc615_5 gpc52 (
      {stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage0_12[34]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[9],stage1_13[12],stage1_12[16],stage1_11[22]}
   );
   gpc606_5 gpc53 (
      {stage0_12[35], stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[5],stage1_14[10],stage1_13[13],stage1_12[17]}
   );
   gpc606_5 gpc54 (
      {stage0_12[41], stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[6],stage1_14[11],stage1_13[14],stage1_12[18]}
   );
   gpc606_5 gpc55 (
      {stage0_12[47], stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[7],stage1_14[12],stage1_13[15],stage1_12[19]}
   );
   gpc606_5 gpc56 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[3],stage1_15[8],stage1_14[13],stage1_13[16]}
   );
   gpc606_5 gpc57 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[4],stage1_15[9],stage1_14[14],stage1_13[17]}
   );
   gpc606_5 gpc58 (
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[2],stage1_16[5],stage1_15[10],stage1_14[15]}
   );
   gpc606_5 gpc59 (
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[3],stage1_16[6],stage1_15[11],stage1_14[16]}
   );
   gpc606_5 gpc60 (
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[4],stage1_16[7],stage1_15[12],stage1_14[17]}
   );
   gpc615_5 gpc61 (
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40]},
      {stage0_15[12]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23]},
      {stage1_18[3],stage1_17[5],stage1_16[8],stage1_15[13],stage1_14[18]}
   );
   gpc615_5 gpc62 (
      {stage0_14[41], stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45]},
      {stage0_15[13]},
      {stage0_16[24], stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29]},
      {stage1_18[4],stage1_17[6],stage1_16[9],stage1_15[14],stage1_14[19]}
   );
   gpc615_5 gpc63 (
      {stage0_14[46], stage0_14[47], stage0_14[48], stage0_14[49], stage0_14[50]},
      {stage0_15[14]},
      {stage0_16[30], stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35]},
      {stage1_18[5],stage1_17[7],stage1_16[10],stage1_15[15],stage1_14[20]}
   );
   gpc615_5 gpc64 (
      {stage0_15[15], stage0_15[16], stage0_15[17], stage0_15[18], stage0_15[19]},
      {stage0_16[36]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[6],stage1_17[8],stage1_16[11],stage1_15[16]}
   );
   gpc615_5 gpc65 (
      {stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23], stage0_15[24]},
      {stage0_16[37]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[7],stage1_17[9],stage1_16[12],stage1_15[17]}
   );
   gpc615_5 gpc66 (
      {stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage0_16[38]},
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage1_19[2],stage1_18[8],stage1_17[10],stage1_16[13],stage1_15[18]}
   );
   gpc606_5 gpc67 (
      {stage0_16[39], stage0_16[40], stage0_16[41], stage0_16[42], stage0_16[43], stage0_16[44]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[3],stage1_18[9],stage1_17[11],stage1_16[14]}
   );
   gpc606_5 gpc68 (
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[1],stage1_19[4],stage1_18[10],stage1_17[12]}
   );
   gpc606_5 gpc69 (
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[2],stage1_19[5],stage1_18[11],stage1_17[13]}
   );
   gpc606_5 gpc70 (
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[3],stage1_19[6],stage1_18[12],stage1_17[14]}
   );
   gpc606_5 gpc71 (
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[4],stage1_19[7],stage1_18[13],stage1_17[15]}
   );
   gpc606_5 gpc72 (
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[5],stage1_19[8],stage1_18[14],stage1_17[16]}
   );
   gpc606_5 gpc73 (
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[6],stage1_19[9],stage1_18[15],stage1_17[17]}
   );
   gpc606_5 gpc74 (
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[6],stage1_20[7],stage1_19[10],stage1_18[16]}
   );
   gpc606_5 gpc75 (
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[7],stage1_20[8],stage1_19[11],stage1_18[17]}
   );
   gpc606_5 gpc76 (
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[8],stage1_20[9],stage1_19[12],stage1_18[18]}
   );
   gpc606_5 gpc77 (
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[9],stage1_20[10],stage1_19[13],stage1_18[19]}
   );
   gpc606_5 gpc78 (
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29]},
      {stage1_22[4],stage1_21[10],stage1_20[11],stage1_19[14],stage1_18[20]}
   );
   gpc606_5 gpc79 (
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35]},
      {stage1_22[5],stage1_21[11],stage1_20[12],stage1_19[15],stage1_18[21]}
   );
   gpc606_5 gpc80 (
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[6],stage1_21[12],stage1_20[13],stage1_19[16]}
   );
   gpc615_5 gpc81 (
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46]},
      {stage0_20[36]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[7],stage1_21[13],stage1_20[14],stage1_19[17]}
   );
   gpc615_5 gpc82 (
      {stage0_19[47], stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51]},
      {stage0_20[37]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[8],stage1_21[14],stage1_20[15],stage1_19[18]}
   );
   gpc615_5 gpc83 (
      {stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41], stage0_20[42]},
      {stage0_21[18]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[3],stage1_22[9],stage1_21[15],stage1_20[16]}
   );
   gpc615_5 gpc84 (
      {stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage0_21[19]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[4],stage1_22[10],stage1_21[16],stage1_20[17]}
   );
   gpc615_5 gpc85 (
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52]},
      {stage0_21[20]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[5],stage1_22[11],stage1_21[17],stage1_20[18]}
   );
   gpc606_5 gpc86 (
      {stage0_21[21], stage0_21[22], stage0_21[23], stage0_21[24], stage0_21[25], stage0_21[26]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[3],stage1_23[6],stage1_22[12],stage1_21[18]}
   );
   gpc606_5 gpc87 (
      {stage0_21[27], stage0_21[28], stage0_21[29], stage0_21[30], stage0_21[31], stage0_21[32]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[4],stage1_23[7],stage1_22[13],stage1_21[19]}
   );
   gpc606_5 gpc88 (
      {stage0_21[33], stage0_21[34], stage0_21[35], stage0_21[36], stage0_21[37], stage0_21[38]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[5],stage1_23[8],stage1_22[14],stage1_21[20]}
   );
   gpc606_5 gpc89 (
      {stage0_21[39], stage0_21[40], stage0_21[41], stage0_21[42], stage0_21[43], stage0_21[44]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[6],stage1_23[9],stage1_22[15],stage1_21[21]}
   );
   gpc606_5 gpc90 (
      {stage0_21[45], stage0_21[46], stage0_21[47], stage0_21[48], stage0_21[49], stage0_21[50]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[7],stage1_23[10],stage1_22[16],stage1_21[22]}
   );
   gpc606_5 gpc91 (
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[5],stage1_24[8],stage1_23[11],stage1_22[17]}
   );
   gpc606_5 gpc92 (
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[6],stage1_24[9],stage1_23[12],stage1_22[18]}
   );
   gpc606_5 gpc93 (
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[7],stage1_24[10],stage1_23[13],stage1_22[19]}
   );
   gpc606_5 gpc94 (
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[8],stage1_24[11],stage1_23[14],stage1_22[20]}
   );
   gpc606_5 gpc95 (
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[9],stage1_24[12],stage1_23[15],stage1_22[21]}
   );
   gpc606_5 gpc96 (
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[10],stage1_24[13],stage1_23[16],stage1_22[22]}
   );
   gpc615_5 gpc97 (
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34]},
      {stage0_24[36]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[6],stage1_25[11],stage1_24[14],stage1_23[17]}
   );
   gpc615_5 gpc98 (
      {stage0_23[35], stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39]},
      {stage0_24[37]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[7],stage1_25[12],stage1_24[15],stage1_23[18]}
   );
   gpc615_5 gpc99 (
      {stage0_23[40], stage0_23[41], stage0_23[42], stage0_23[43], stage0_23[44]},
      {stage0_24[38]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[8],stage1_25[13],stage1_24[16],stage1_23[19]}
   );
   gpc615_5 gpc100 (
      {stage0_23[45], stage0_23[46], stage0_23[47], stage0_23[48], stage0_23[49]},
      {stage0_24[39]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[9],stage1_25[14],stage1_24[17],stage1_23[20]}
   );
   gpc615_5 gpc101 (
      {stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53], 1'b0},
      {stage0_24[40]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[10],stage1_25[15],stage1_24[18],stage1_23[21]}
   );
   gpc606_5 gpc102 (
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[0],stage1_27[5],stage1_26[11],stage1_25[16]}
   );
   gpc606_5 gpc103 (
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[1],stage1_27[6],stage1_26[12],stage1_25[17]}
   );
   gpc606_5 gpc104 (
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[2],stage1_27[7],stage1_26[13],stage1_25[18]}
   );
   gpc2135_5 gpc105 (
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4]},
      {stage0_27[18], stage0_27[19], stage0_27[20]},
      {stage0_28[0]},
      {stage0_29[0], stage0_29[1]},
      {stage1_30[0],stage1_29[3],stage1_28[3],stage1_27[8],stage1_26[14]}
   );
   gpc2135_5 gpc106 (
      {stage0_26[5], stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9]},
      {stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage0_28[1]},
      {stage0_29[2], stage0_29[3]},
      {stage1_30[1],stage1_29[4],stage1_28[4],stage1_27[9],stage1_26[15]}
   );
   gpc2135_5 gpc107 (
      {stage0_26[10], stage0_26[11], stage0_26[12], stage0_26[13], stage0_26[14]},
      {stage0_27[24], stage0_27[25], stage0_27[26]},
      {stage0_28[2]},
      {stage0_29[4], stage0_29[5]},
      {stage1_30[2],stage1_29[5],stage1_28[5],stage1_27[10],stage1_26[16]}
   );
   gpc2135_5 gpc108 (
      {stage0_26[15], stage0_26[16], stage0_26[17], stage0_26[18], stage0_26[19]},
      {stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage0_28[3]},
      {stage0_29[6], stage0_29[7]},
      {stage1_30[3],stage1_29[6],stage1_28[6],stage1_27[11],stage1_26[17]}
   );
   gpc615_5 gpc109 (
      {stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23], stage0_26[24]},
      {stage0_27[30]},
      {stage0_28[4], stage0_28[5], stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9]},
      {stage1_30[4],stage1_29[7],stage1_28[7],stage1_27[12],stage1_26[18]}
   );
   gpc615_5 gpc110 (
      {stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage0_27[31]},
      {stage0_28[10], stage0_28[11], stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15]},
      {stage1_30[5],stage1_29[8],stage1_28[8],stage1_27[13],stage1_26[19]}
   );
   gpc615_5 gpc111 (
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34]},
      {stage0_27[32]},
      {stage0_28[16], stage0_28[17], stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21]},
      {stage1_30[6],stage1_29[9],stage1_28[9],stage1_27[14],stage1_26[20]}
   );
   gpc615_5 gpc112 (
      {stage0_26[35], stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39]},
      {stage0_27[33]},
      {stage0_28[22], stage0_28[23], stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27]},
      {stage1_30[7],stage1_29[10],stage1_28[10],stage1_27[15],stage1_26[21]}
   );
   gpc615_5 gpc113 (
      {stage0_26[40], stage0_26[41], stage0_26[42], stage0_26[43], stage0_26[44]},
      {stage0_27[34]},
      {stage0_28[28], stage0_28[29], stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33]},
      {stage1_30[8],stage1_29[11],stage1_28[11],stage1_27[16],stage1_26[22]}
   );
   gpc615_5 gpc114 (
      {stage0_27[35], stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39]},
      {stage0_28[34]},
      {stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11], stage0_29[12], stage0_29[13]},
      {stage1_31[0],stage1_30[9],stage1_29[12],stage1_28[12],stage1_27[17]}
   );
   gpc615_5 gpc115 (
      {stage0_27[40], stage0_27[41], stage0_27[42], stage0_27[43], stage0_27[44]},
      {stage0_28[35]},
      {stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17], stage0_29[18], stage0_29[19]},
      {stage1_31[1],stage1_30[10],stage1_29[13],stage1_28[13],stage1_27[18]}
   );
   gpc615_5 gpc116 (
      {stage0_27[45], stage0_27[46], stage0_27[47], stage0_27[48], stage0_27[49]},
      {stage0_28[36]},
      {stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23], stage0_29[24], stage0_29[25]},
      {stage1_31[2],stage1_30[11],stage1_29[14],stage1_28[14],stage1_27[19]}
   );
   gpc606_5 gpc117 (
      {stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41], stage0_28[42]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[3],stage1_30[12],stage1_29[15],stage1_28[15]}
   );
   gpc606_5 gpc118 (
      {stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46], stage0_28[47], stage0_28[48]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[4],stage1_30[13],stage1_29[16],stage1_28[16]}
   );
   gpc606_5 gpc119 (
      {stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52], stage0_28[53], 1'b0},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[5],stage1_30[14],stage1_29[17],stage1_28[17]}
   );
   gpc606_5 gpc120 (
      {stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29], stage0_29[30], stage0_29[31]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[3],stage1_31[6],stage1_30[15],stage1_29[18]}
   );
   gpc606_5 gpc121 (
      {stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35], stage0_29[36], stage0_29[37]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[4],stage1_31[7],stage1_30[16],stage1_29[19]}
   );
   gpc606_5 gpc122 (
      {stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41], stage0_29[42], stage0_29[43]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[5],stage1_31[8],stage1_30[17],stage1_29[20]}
   );
   gpc606_5 gpc123 (
      {stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47], stage0_29[48], stage0_29[49]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[6],stage1_31[9],stage1_30[18],stage1_29[21]}
   );
   gpc606_5 gpc124 (
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3], stage0_32[4], stage0_32[5]},
      {stage1_34[0],stage1_33[4],stage1_32[7],stage1_31[10],stage1_30[19]}
   );
   gpc606_5 gpc125 (
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage0_32[6], stage0_32[7], stage0_32[8], stage0_32[9], stage0_32[10], stage0_32[11]},
      {stage1_34[1],stage1_33[5],stage1_32[8],stage1_31[11],stage1_30[20]}
   );
   gpc606_5 gpc126 (
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage0_32[12], stage0_32[13], stage0_32[14], stage0_32[15], stage0_32[16], stage0_32[17]},
      {stage1_34[2],stage1_33[6],stage1_32[9],stage1_31[12],stage1_30[21]}
   );
   gpc606_5 gpc127 (
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage0_32[18], stage0_32[19], stage0_32[20], stage0_32[21], stage0_32[22], stage0_32[23]},
      {stage1_34[3],stage1_33[7],stage1_32[10],stage1_31[13],stage1_30[22]}
   );
   gpc606_5 gpc128 (
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage0_33[0], stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5]},
      {stage1_35[0],stage1_34[4],stage1_33[8],stage1_32[11],stage1_31[14]}
   );
   gpc606_5 gpc129 (
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage0_33[6], stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11]},
      {stage1_35[1],stage1_34[5],stage1_33[9],stage1_32[12],stage1_31[15]}
   );
   gpc606_5 gpc130 (
      {stage0_32[24], stage0_32[25], stage0_32[26], stage0_32[27], stage0_32[28], stage0_32[29]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[2],stage1_34[6],stage1_33[10],stage1_32[13]}
   );
   gpc606_5 gpc131 (
      {stage0_32[30], stage0_32[31], stage0_32[32], stage0_32[33], stage0_32[34], stage0_32[35]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[3],stage1_34[7],stage1_33[11],stage1_32[14]}
   );
   gpc606_5 gpc132 (
      {stage0_32[36], stage0_32[37], stage0_32[38], stage0_32[39], stage0_32[40], stage0_32[41]},
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17]},
      {stage1_36[2],stage1_35[4],stage1_34[8],stage1_33[12],stage1_32[15]}
   );
   gpc606_5 gpc133 (
      {stage0_32[42], stage0_32[43], stage0_32[44], stage0_32[45], stage0_32[46], stage0_32[47]},
      {stage0_34[18], stage0_34[19], stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23]},
      {stage1_36[3],stage1_35[5],stage1_34[9],stage1_33[13],stage1_32[16]}
   );
   gpc615_5 gpc134 (
      {stage0_32[48], stage0_32[49], stage0_32[50], stage0_32[51], stage0_32[52]},
      {stage0_33[12]},
      {stage0_34[24], stage0_34[25], stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29]},
      {stage1_36[4],stage1_35[6],stage1_34[10],stage1_33[14],stage1_32[17]}
   );
   gpc606_5 gpc135 (
      {stage0_33[13], stage0_33[14], stage0_33[15], stage0_33[16], stage0_33[17], stage0_33[18]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[5],stage1_35[7],stage1_34[11],stage1_33[15]}
   );
   gpc606_5 gpc136 (
      {stage0_33[19], stage0_33[20], stage0_33[21], stage0_33[22], stage0_33[23], stage0_33[24]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[6],stage1_35[8],stage1_34[12],stage1_33[16]}
   );
   gpc117_4 gpc137 (
      {stage0_34[30], stage0_34[31], stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35], stage0_34[36]},
      {stage0_35[12]},
      {stage0_36[0]},
      {stage1_37[2],stage1_36[7],stage1_35[9],stage1_34[13]}
   );
   gpc117_4 gpc138 (
      {stage0_34[37], stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41], stage0_34[42], stage0_34[43]},
      {stage0_35[13]},
      {stage0_36[1]},
      {stage1_37[3],stage1_36[8],stage1_35[10],stage1_34[14]}
   );
   gpc117_4 gpc139 (
      {stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47], stage0_34[48], stage0_34[49], stage0_34[50]},
      {stage0_35[14]},
      {stage0_36[2]},
      {stage1_37[4],stage1_36[9],stage1_35[11],stage1_34[15]}
   );
   gpc606_5 gpc140 (
      {stage0_35[15], stage0_35[16], stage0_35[17], stage0_35[18], stage0_35[19], stage0_35[20]},
      {stage0_37[0], stage0_37[1], stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5]},
      {stage1_39[0],stage1_38[0],stage1_37[5],stage1_36[10],stage1_35[12]}
   );
   gpc606_5 gpc141 (
      {stage0_35[21], stage0_35[22], stage0_35[23], stage0_35[24], stage0_35[25], stage0_35[26]},
      {stage0_37[6], stage0_37[7], stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11]},
      {stage1_39[1],stage1_38[1],stage1_37[6],stage1_36[11],stage1_35[13]}
   );
   gpc606_5 gpc142 (
      {stage0_35[27], stage0_35[28], stage0_35[29], stage0_35[30], stage0_35[31], stage0_35[32]},
      {stage0_37[12], stage0_37[13], stage0_37[14], stage0_37[15], stage0_37[16], stage0_37[17]},
      {stage1_39[2],stage1_38[2],stage1_37[7],stage1_36[12],stage1_35[14]}
   );
   gpc615_5 gpc143 (
      {stage0_35[33], stage0_35[34], stage0_35[35], stage0_35[36], stage0_35[37]},
      {stage0_36[3]},
      {stage0_37[18], stage0_37[19], stage0_37[20], stage0_37[21], stage0_37[22], stage0_37[23]},
      {stage1_39[3],stage1_38[3],stage1_37[8],stage1_36[13],stage1_35[15]}
   );
   gpc615_5 gpc144 (
      {stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41], stage0_35[42]},
      {stage0_36[4]},
      {stage0_37[24], stage0_37[25], stage0_37[26], stage0_37[27], stage0_37[28], stage0_37[29]},
      {stage1_39[4],stage1_38[4],stage1_37[9],stage1_36[14],stage1_35[16]}
   );
   gpc606_5 gpc145 (
      {stage0_36[5], stage0_36[6], stage0_36[7], stage0_36[8], stage0_36[9], stage0_36[10]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[5],stage1_38[5],stage1_37[10],stage1_36[15]}
   );
   gpc606_5 gpc146 (
      {stage0_36[11], stage0_36[12], stage0_36[13], stage0_36[14], stage0_36[15], stage0_36[16]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[6],stage1_38[6],stage1_37[11],stage1_36[16]}
   );
   gpc606_5 gpc147 (
      {stage0_36[17], stage0_36[18], stage0_36[19], stage0_36[20], stage0_36[21], stage0_36[22]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[7],stage1_38[7],stage1_37[12],stage1_36[17]}
   );
   gpc606_5 gpc148 (
      {stage0_36[23], stage0_36[24], stage0_36[25], stage0_36[26], stage0_36[27], stage0_36[28]},
      {stage0_38[18], stage0_38[19], stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23]},
      {stage1_40[3],stage1_39[8],stage1_38[8],stage1_37[13],stage1_36[18]}
   );
   gpc606_5 gpc149 (
      {stage0_36[29], stage0_36[30], stage0_36[31], stage0_36[32], stage0_36[33], stage0_36[34]},
      {stage0_38[24], stage0_38[25], stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29]},
      {stage1_40[4],stage1_39[9],stage1_38[9],stage1_37[14],stage1_36[19]}
   );
   gpc606_5 gpc150 (
      {stage0_36[35], stage0_36[36], stage0_36[37], stage0_36[38], stage0_36[39], stage0_36[40]},
      {stage0_38[30], stage0_38[31], stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35]},
      {stage1_40[5],stage1_39[10],stage1_38[10],stage1_37[15],stage1_36[20]}
   );
   gpc606_5 gpc151 (
      {stage0_37[30], stage0_37[31], stage0_37[32], stage0_37[33], stage0_37[34], stage0_37[35]},
      {stage0_39[0], stage0_39[1], stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5]},
      {stage1_41[0],stage1_40[6],stage1_39[11],stage1_38[11],stage1_37[16]}
   );
   gpc606_5 gpc152 (
      {stage0_37[36], stage0_37[37], stage0_37[38], stage0_37[39], stage0_37[40], stage0_37[41]},
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage1_41[1],stage1_40[7],stage1_39[12],stage1_38[12],stage1_37[17]}
   );
   gpc606_5 gpc153 (
      {stage0_37[42], stage0_37[43], stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47]},
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage1_41[2],stage1_40[8],stage1_39[13],stage1_38[13],stage1_37[18]}
   );
   gpc615_5 gpc154 (
      {stage0_38[36], stage0_38[37], stage0_38[38], stage0_38[39], stage0_38[40]},
      {stage0_39[18]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[3],stage1_40[9],stage1_39[14],stage1_38[14]}
   );
   gpc615_5 gpc155 (
      {stage0_38[41], stage0_38[42], stage0_38[43], stage0_38[44], stage0_38[45]},
      {stage0_39[19]},
      {stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11]},
      {stage1_42[1],stage1_41[4],stage1_40[10],stage1_39[15],stage1_38[15]}
   );
   gpc606_5 gpc156 (
      {stage0_39[20], stage0_39[21], stage0_39[22], stage0_39[23], stage0_39[24], stage0_39[25]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[2],stage1_41[5],stage1_40[11],stage1_39[16]}
   );
   gpc606_5 gpc157 (
      {stage0_39[26], stage0_39[27], stage0_39[28], stage0_39[29], stage0_39[30], stage0_39[31]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[3],stage1_41[6],stage1_40[12],stage1_39[17]}
   );
   gpc606_5 gpc158 (
      {stage0_39[32], stage0_39[33], stage0_39[34], stage0_39[35], stage0_39[36], stage0_39[37]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[4],stage1_41[7],stage1_40[13],stage1_39[18]}
   );
   gpc615_5 gpc159 (
      {stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41], stage0_39[42]},
      {stage0_40[12]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[5],stage1_41[8],stage1_40[14],stage1_39[19]}
   );
   gpc1406_5 gpc160 (
      {stage0_40[13], stage0_40[14], stage0_40[15], stage0_40[16], stage0_40[17], stage0_40[18]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3]},
      {stage0_43[0]},
      {stage1_44[0],stage1_43[4],stage1_42[6],stage1_41[9],stage1_40[15]}
   );
   gpc615_5 gpc161 (
      {stage0_40[19], stage0_40[20], stage0_40[21], stage0_40[22], stage0_40[23]},
      {stage0_41[24]},
      {stage0_42[4], stage0_42[5], stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9]},
      {stage1_44[1],stage1_43[5],stage1_42[7],stage1_41[10],stage1_40[16]}
   );
   gpc615_5 gpc162 (
      {stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27], stage0_40[28]},
      {stage0_41[25]},
      {stage0_42[10], stage0_42[11], stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15]},
      {stage1_44[2],stage1_43[6],stage1_42[8],stage1_41[11],stage1_40[17]}
   );
   gpc615_5 gpc163 (
      {stage0_40[29], stage0_40[30], stage0_40[31], stage0_40[32], stage0_40[33]},
      {stage0_41[26]},
      {stage0_42[16], stage0_42[17], stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21]},
      {stage1_44[3],stage1_43[7],stage1_42[9],stage1_41[12],stage1_40[18]}
   );
   gpc606_5 gpc164 (
      {stage0_41[27], stage0_41[28], stage0_41[29], stage0_41[30], stage0_41[31], stage0_41[32]},
      {stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5], stage0_43[6]},
      {stage1_45[0],stage1_44[4],stage1_43[8],stage1_42[10],stage1_41[13]}
   );
   gpc606_5 gpc165 (
      {stage0_41[33], stage0_41[34], stage0_41[35], stage0_41[36], stage0_41[37], stage0_41[38]},
      {stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11], stage0_43[12]},
      {stage1_45[1],stage1_44[5],stage1_43[9],stage1_42[11],stage1_41[14]}
   );
   gpc606_5 gpc166 (
      {stage0_41[39], stage0_41[40], stage0_41[41], stage0_41[42], stage0_41[43], stage0_41[44]},
      {stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17], stage0_43[18]},
      {stage1_45[2],stage1_44[6],stage1_43[10],stage1_42[12],stage1_41[15]}
   );
   gpc606_5 gpc167 (
      {stage0_41[45], stage0_41[46], stage0_41[47], stage0_41[48], stage0_41[49], stage0_41[50]},
      {stage0_43[19], stage0_43[20], stage0_43[21], stage0_43[22], stage0_43[23], stage0_43[24]},
      {stage1_45[3],stage1_44[7],stage1_43[11],stage1_42[13],stage1_41[16]}
   );
   gpc606_5 gpc168 (
      {stage0_42[22], stage0_42[23], stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[4],stage1_44[8],stage1_43[12],stage1_42[14]}
   );
   gpc606_5 gpc169 (
      {stage0_42[28], stage0_42[29], stage0_42[30], stage0_42[31], stage0_42[32], stage0_42[33]},
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11]},
      {stage1_46[1],stage1_45[5],stage1_44[9],stage1_43[13],stage1_42[15]}
   );
   gpc606_5 gpc170 (
      {stage0_42[34], stage0_42[35], stage0_42[36], stage0_42[37], stage0_42[38], stage0_42[39]},
      {stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15], stage0_44[16], stage0_44[17]},
      {stage1_46[2],stage1_45[6],stage1_44[10],stage1_43[14],stage1_42[16]}
   );
   gpc606_5 gpc171 (
      {stage0_42[40], stage0_42[41], stage0_42[42], stage0_42[43], stage0_42[44], stage0_42[45]},
      {stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21], stage0_44[22], stage0_44[23]},
      {stage1_46[3],stage1_45[7],stage1_44[11],stage1_43[15],stage1_42[17]}
   );
   gpc606_5 gpc172 (
      {stage0_42[46], stage0_42[47], stage0_42[48], stage0_42[49], stage0_42[50], stage0_42[51]},
      {stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27], stage0_44[28], stage0_44[29]},
      {stage1_46[4],stage1_45[8],stage1_44[12],stage1_43[16],stage1_42[18]}
   );
   gpc615_5 gpc173 (
      {stage0_43[25], stage0_43[26], stage0_43[27], stage0_43[28], stage0_43[29]},
      {stage0_44[30]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[5],stage1_45[9],stage1_44[13],stage1_43[17]}
   );
   gpc615_5 gpc174 (
      {stage0_43[30], stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34]},
      {stage0_44[31]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[6],stage1_45[10],stage1_44[14],stage1_43[18]}
   );
   gpc615_5 gpc175 (
      {stage0_43[35], stage0_43[36], stage0_43[37], stage0_43[38], stage0_43[39]},
      {stage0_44[32]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[7],stage1_45[11],stage1_44[15],stage1_43[19]}
   );
   gpc615_5 gpc176 (
      {stage0_43[40], stage0_43[41], stage0_43[42], stage0_43[43], stage0_43[44]},
      {stage0_44[33]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[8],stage1_45[12],stage1_44[16],stage1_43[20]}
   );
   gpc615_5 gpc177 (
      {stage0_43[45], stage0_43[46], stage0_43[47], stage0_43[48], stage0_43[49]},
      {stage0_44[34]},
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage1_47[4],stage1_46[9],stage1_45[13],stage1_44[17],stage1_43[21]}
   );
   gpc615_5 gpc178 (
      {stage0_43[50], stage0_43[51], stage0_43[52], stage0_43[53], 1'b0},
      {stage0_44[35]},
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage1_47[5],stage1_46[10],stage1_45[14],stage1_44[18],stage1_43[22]}
   );
   gpc606_5 gpc179 (
      {stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39], stage0_44[40], stage0_44[41]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[6],stage1_46[11],stage1_45[15],stage1_44[19]}
   );
   gpc606_5 gpc180 (
      {stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45], stage0_44[46], stage0_44[47]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[7],stage1_46[12],stage1_45[16],stage1_44[20]}
   );
   gpc606_5 gpc181 (
      {stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51], stage0_44[52], stage0_44[53]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[8],stage1_46[13],stage1_45[17],stage1_44[21]}
   );
   gpc615_5 gpc182 (
      {stage0_45[36], stage0_45[37], stage0_45[38], stage0_45[39], stage0_45[40]},
      {stage0_46[18]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[3],stage1_47[9],stage1_46[14],stage1_45[18]}
   );
   gpc615_5 gpc183 (
      {stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage0_47[6]},
      {stage0_48[0], stage0_48[1], stage0_48[2], stage0_48[3], stage0_48[4], stage0_48[5]},
      {stage1_50[0],stage1_49[1],stage1_48[4],stage1_47[10],stage1_46[15]}
   );
   gpc615_5 gpc184 (
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28]},
      {stage0_47[7]},
      {stage0_48[6], stage0_48[7], stage0_48[8], stage0_48[9], stage0_48[10], stage0_48[11]},
      {stage1_50[1],stage1_49[2],stage1_48[5],stage1_47[11],stage1_46[16]}
   );
   gpc615_5 gpc185 (
      {stage0_46[29], stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33]},
      {stage0_47[8]},
      {stage0_48[12], stage0_48[13], stage0_48[14], stage0_48[15], stage0_48[16], stage0_48[17]},
      {stage1_50[2],stage1_49[3],stage1_48[6],stage1_47[12],stage1_46[17]}
   );
   gpc615_5 gpc186 (
      {stage0_46[34], stage0_46[35], stage0_46[36], stage0_46[37], stage0_46[38]},
      {stage0_47[9]},
      {stage0_48[18], stage0_48[19], stage0_48[20], stage0_48[21], stage0_48[22], stage0_48[23]},
      {stage1_50[3],stage1_49[4],stage1_48[7],stage1_47[13],stage1_46[18]}
   );
   gpc615_5 gpc187 (
      {stage0_46[39], stage0_46[40], stage0_46[41], stage0_46[42], stage0_46[43]},
      {stage0_47[10]},
      {stage0_48[24], stage0_48[25], stage0_48[26], stage0_48[27], stage0_48[28], stage0_48[29]},
      {stage1_50[4],stage1_49[5],stage1_48[8],stage1_47[14],stage1_46[19]}
   );
   gpc615_5 gpc188 (
      {stage0_47[11], stage0_47[12], stage0_47[13], stage0_47[14], stage0_47[15]},
      {stage0_48[30]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[5],stage1_49[6],stage1_48[9],stage1_47[15]}
   );
   gpc615_5 gpc189 (
      {stage0_47[16], stage0_47[17], stage0_47[18], stage0_47[19], stage0_47[20]},
      {stage0_48[31]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[6],stage1_49[7],stage1_48[10],stage1_47[16]}
   );
   gpc615_5 gpc190 (
      {stage0_47[21], stage0_47[22], stage0_47[23], stage0_47[24], stage0_47[25]},
      {stage0_48[32]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[7],stage1_49[8],stage1_48[11],stage1_47[17]}
   );
   gpc615_5 gpc191 (
      {stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29], stage0_47[30]},
      {stage0_48[33]},
      {stage0_49[18], stage0_49[19], stage0_49[20], stage0_49[21], stage0_49[22], stage0_49[23]},
      {stage1_51[3],stage1_50[8],stage1_49[9],stage1_48[12],stage1_47[18]}
   );
   gpc615_5 gpc192 (
      {stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage0_48[34]},
      {stage0_49[24], stage0_49[25], stage0_49[26], stage0_49[27], stage0_49[28], stage0_49[29]},
      {stage1_51[4],stage1_50[9],stage1_49[10],stage1_48[13],stage1_47[19]}
   );
   gpc615_5 gpc193 (
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40]},
      {stage0_48[35]},
      {stage0_49[30], stage0_49[31], stage0_49[32], stage0_49[33], stage0_49[34], stage0_49[35]},
      {stage1_51[5],stage1_50[10],stage1_49[11],stage1_48[14],stage1_47[20]}
   );
   gpc606_5 gpc194 (
      {stage0_48[36], stage0_48[37], stage0_48[38], stage0_48[39], stage0_48[40], stage0_48[41]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[6],stage1_50[11],stage1_49[12],stage1_48[15]}
   );
   gpc606_5 gpc195 (
      {stage0_48[42], stage0_48[43], stage0_48[44], stage0_48[45], stage0_48[46], stage0_48[47]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[7],stage1_50[12],stage1_49[13],stage1_48[16]}
   );
   gpc606_5 gpc196 (
      {stage0_48[48], stage0_48[49], stage0_48[50], stage0_48[51], stage0_48[52], stage0_48[53]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[8],stage1_50[13],stage1_49[14],stage1_48[17]}
   );
   gpc606_5 gpc197 (
      {stage0_49[36], stage0_49[37], stage0_49[38], stage0_49[39], stage0_49[40], stage0_49[41]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[3],stage1_51[9],stage1_50[14],stage1_49[15]}
   );
   gpc615_5 gpc198 (
      {stage0_49[42], stage0_49[43], stage0_49[44], stage0_49[45], stage0_49[46]},
      {stage0_50[18]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[4],stage1_51[10],stage1_50[15],stage1_49[16]}
   );
   gpc615_5 gpc199 (
      {stage0_50[19], stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23]},
      {stage0_51[12]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[2],stage1_52[5],stage1_51[11],stage1_50[16]}
   );
   gpc615_5 gpc200 (
      {stage0_50[24], stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28]},
      {stage0_51[13]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[3],stage1_52[6],stage1_51[12],stage1_50[17]}
   );
   gpc606_5 gpc201 (
      {stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17], stage0_51[18], stage0_51[19]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[2],stage1_53[4],stage1_52[7],stage1_51[13]}
   );
   gpc615_5 gpc202 (
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16]},
      {stage0_53[6]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[1],stage1_54[3],stage1_53[5],stage1_52[8]}
   );
   gpc615_5 gpc203 (
      {stage0_52[17], stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21]},
      {stage0_53[7]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[2],stage1_54[4],stage1_53[6],stage1_52[9]}
   );
   gpc615_5 gpc204 (
      {stage0_52[22], stage0_52[23], stage0_52[24], stage0_52[25], stage0_52[26]},
      {stage0_53[8]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[3],stage1_54[5],stage1_53[7],stage1_52[10]}
   );
   gpc615_5 gpc205 (
      {stage0_52[27], stage0_52[28], stage0_52[29], stage0_52[30], stage0_52[31]},
      {stage0_53[9]},
      {stage0_54[18], stage0_54[19], stage0_54[20], stage0_54[21], stage0_54[22], stage0_54[23]},
      {stage1_56[3],stage1_55[4],stage1_54[6],stage1_53[8],stage1_52[11]}
   );
   gpc615_5 gpc206 (
      {stage0_52[32], stage0_52[33], stage0_52[34], stage0_52[35], stage0_52[36]},
      {stage0_53[10]},
      {stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27], stage0_54[28], stage0_54[29]},
      {stage1_56[4],stage1_55[5],stage1_54[7],stage1_53[9],stage1_52[12]}
   );
   gpc615_5 gpc207 (
      {stage0_52[37], stage0_52[38], stage0_52[39], stage0_52[40], stage0_52[41]},
      {stage0_53[11]},
      {stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33], stage0_54[34], stage0_54[35]},
      {stage1_56[5],stage1_55[6],stage1_54[8],stage1_53[10],stage1_52[13]}
   );
   gpc615_5 gpc208 (
      {stage0_52[42], stage0_52[43], stage0_52[44], stage0_52[45], stage0_52[46]},
      {stage0_53[12]},
      {stage0_54[36], stage0_54[37], stage0_54[38], stage0_54[39], stage0_54[40], stage0_54[41]},
      {stage1_56[6],stage1_55[7],stage1_54[9],stage1_53[11],stage1_52[14]}
   );
   gpc615_5 gpc209 (
      {stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage0_54[42]},
      {stage0_55[0], stage0_55[1], stage0_55[2], stage0_55[3], stage0_55[4], stage0_55[5]},
      {stage1_57[0],stage1_56[7],stage1_55[8],stage1_54[10],stage1_53[12]}
   );
   gpc615_5 gpc210 (
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22]},
      {stage0_54[43]},
      {stage0_55[6], stage0_55[7], stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11]},
      {stage1_57[1],stage1_56[8],stage1_55[9],stage1_54[11],stage1_53[13]}
   );
   gpc615_5 gpc211 (
      {stage0_53[23], stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27]},
      {stage0_54[44]},
      {stage0_55[12], stage0_55[13], stage0_55[14], stage0_55[15], stage0_55[16], stage0_55[17]},
      {stage1_57[2],stage1_56[9],stage1_55[10],stage1_54[12],stage1_53[14]}
   );
   gpc606_5 gpc212 (
      {stage0_54[45], stage0_54[46], stage0_54[47], stage0_54[48], stage0_54[49], stage0_54[50]},
      {stage0_56[0], stage0_56[1], stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5]},
      {stage1_58[0],stage1_57[3],stage1_56[10],stage1_55[11],stage1_54[13]}
   );
   gpc606_5 gpc213 (
      {stage0_55[18], stage0_55[19], stage0_55[20], stage0_55[21], stage0_55[22], stage0_55[23]},
      {stage0_57[0], stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5]},
      {stage1_59[0],stage1_58[1],stage1_57[4],stage1_56[11],stage1_55[12]}
   );
   gpc606_5 gpc214 (
      {stage0_55[24], stage0_55[25], stage0_55[26], stage0_55[27], stage0_55[28], stage0_55[29]},
      {stage0_57[6], stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11]},
      {stage1_59[1],stage1_58[2],stage1_57[5],stage1_56[12],stage1_55[13]}
   );
   gpc606_5 gpc215 (
      {stage0_56[6], stage0_56[7], stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11]},
      {stage0_58[0], stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5]},
      {stage1_60[0],stage1_59[2],stage1_58[3],stage1_57[6],stage1_56[13]}
   );
   gpc606_5 gpc216 (
      {stage0_56[12], stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17]},
      {stage0_58[6], stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11]},
      {stage1_60[1],stage1_59[3],stage1_58[4],stage1_57[7],stage1_56[14]}
   );
   gpc606_5 gpc217 (
      {stage0_56[18], stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23]},
      {stage0_58[12], stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17]},
      {stage1_60[2],stage1_59[4],stage1_58[5],stage1_57[8],stage1_56[15]}
   );
   gpc606_5 gpc218 (
      {stage0_56[24], stage0_56[25], stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29]},
      {stage0_58[18], stage0_58[19], stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23]},
      {stage1_60[3],stage1_59[5],stage1_58[6],stage1_57[9],stage1_56[16]}
   );
   gpc606_5 gpc219 (
      {stage0_56[30], stage0_56[31], stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35]},
      {stage0_58[24], stage0_58[25], stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29]},
      {stage1_60[4],stage1_59[6],stage1_58[7],stage1_57[10],stage1_56[17]}
   );
   gpc606_5 gpc220 (
      {stage0_56[36], stage0_56[37], stage0_56[38], stage0_56[39], stage0_56[40], stage0_56[41]},
      {stage0_58[30], stage0_58[31], stage0_58[32], stage0_58[33], stage0_58[34], stage0_58[35]},
      {stage1_60[5],stage1_59[7],stage1_58[8],stage1_57[11],stage1_56[18]}
   );
   gpc606_5 gpc221 (
      {stage0_56[42], stage0_56[43], stage0_56[44], stage0_56[45], stage0_56[46], stage0_56[47]},
      {stage0_58[36], stage0_58[37], stage0_58[38], stage0_58[39], stage0_58[40], stage0_58[41]},
      {stage1_60[6],stage1_59[8],stage1_58[9],stage1_57[12],stage1_56[19]}
   );
   gpc606_5 gpc222 (
      {stage0_56[48], stage0_56[49], stage0_56[50], stage0_56[51], stage0_56[52], stage0_56[53]},
      {stage0_58[42], stage0_58[43], stage0_58[44], stage0_58[45], stage0_58[46], stage0_58[47]},
      {stage1_60[7],stage1_59[9],stage1_58[10],stage1_57[13],stage1_56[20]}
   );
   gpc606_5 gpc223 (
      {stage0_57[12], stage0_57[13], stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[8],stage1_59[10],stage1_58[11],stage1_57[14]}
   );
   gpc606_5 gpc224 (
      {stage0_57[18], stage0_57[19], stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[9],stage1_59[11],stage1_58[12],stage1_57[15]}
   );
   gpc606_5 gpc225 (
      {stage0_57[24], stage0_57[25], stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[10],stage1_59[12],stage1_58[13],stage1_57[16]}
   );
   gpc606_5 gpc226 (
      {stage0_58[48], stage0_58[49], stage0_58[50], stage0_58[51], stage0_58[52], stage0_58[53]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3], stage0_60[4], stage0_60[5]},
      {stage1_62[0],stage1_61[3],stage1_60[11],stage1_59[13],stage1_58[14]}
   );
   gpc606_5 gpc227 (
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage0_61[0], stage0_61[1], stage0_61[2], stage0_61[3], stage0_61[4], stage0_61[5]},
      {stage1_63[0],stage1_62[1],stage1_61[4],stage1_60[12],stage1_59[14]}
   );
   gpc606_5 gpc228 (
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage0_61[6], stage0_61[7], stage0_61[8], stage0_61[9], stage0_61[10], stage0_61[11]},
      {stage1_63[1],stage1_62[2],stage1_61[5],stage1_60[13],stage1_59[15]}
   );
   gpc606_5 gpc229 (
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage0_61[12], stage0_61[13], stage0_61[14], stage0_61[15], stage0_61[16], stage0_61[17]},
      {stage1_63[2],stage1_62[3],stage1_61[6],stage1_60[14],stage1_59[16]}
   );
   gpc606_5 gpc230 (
      {stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9], stage0_60[10], stage0_60[11]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5]},
      {stage1_64[0],stage1_63[3],stage1_62[4],stage1_61[7],stage1_60[15]}
   );
   gpc606_5 gpc231 (
      {stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15], stage0_60[16], stage0_60[17]},
      {stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11]},
      {stage1_64[1],stage1_63[4],stage1_62[5],stage1_61[8],stage1_60[16]}
   );
   gpc606_5 gpc232 (
      {stage0_60[18], stage0_60[19], stage0_60[20], stage0_60[21], stage0_60[22], stage0_60[23]},
      {stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17]},
      {stage1_64[2],stage1_63[5],stage1_62[6],stage1_61[9],stage1_60[17]}
   );
   gpc606_5 gpc233 (
      {stage0_60[24], stage0_60[25], stage0_60[26], stage0_60[27], stage0_60[28], stage0_60[29]},
      {stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23]},
      {stage1_64[3],stage1_63[6],stage1_62[7],stage1_61[10],stage1_60[18]}
   );
   gpc606_5 gpc234 (
      {stage0_60[30], stage0_60[31], stage0_60[32], stage0_60[33], stage0_60[34], stage0_60[35]},
      {stage0_62[24], stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29]},
      {stage1_64[4],stage1_63[7],stage1_62[8],stage1_61[11],stage1_60[19]}
   );
   gpc606_5 gpc235 (
      {stage0_60[36], stage0_60[37], stage0_60[38], stage0_60[39], stage0_60[40], stage0_60[41]},
      {stage0_62[30], stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35]},
      {stage1_64[5],stage1_63[8],stage1_62[9],stage1_61[12],stage1_60[20]}
   );
   gpc606_5 gpc236 (
      {stage0_60[42], stage0_60[43], stage0_60[44], stage0_60[45], stage0_60[46], stage0_60[47]},
      {stage0_62[36], stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41]},
      {stage1_64[6],stage1_63[9],stage1_62[10],stage1_61[13],stage1_60[21]}
   );
   gpc606_5 gpc237 (
      {stage0_60[48], stage0_60[49], stage0_60[50], stage0_60[51], stage0_60[52], stage0_60[53]},
      {stage0_62[42], stage0_62[43], stage0_62[44], stage0_62[45], stage0_62[46], stage0_62[47]},
      {stage1_64[7],stage1_63[10],stage1_62[11],stage1_61[14],stage1_60[22]}
   );
   gpc606_5 gpc238 (
      {stage0_61[18], stage0_61[19], stage0_61[20], stage0_61[21], stage0_61[22], stage0_61[23]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[8],stage1_63[11],stage1_62[12],stage1_61[15]}
   );
   gpc606_5 gpc239 (
      {stage0_61[24], stage0_61[25], stage0_61[26], stage0_61[27], stage0_61[28], stage0_61[29]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[9],stage1_63[12],stage1_62[13],stage1_61[16]}
   );
   gpc606_5 gpc240 (
      {stage0_61[30], stage0_61[31], stage0_61[32], stage0_61[33], stage0_61[34], stage0_61[35]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[10],stage1_63[13],stage1_62[14],stage1_61[17]}
   );
   gpc606_5 gpc241 (
      {stage0_61[36], stage0_61[37], stage0_61[38], stage0_61[39], stage0_61[40], stage0_61[41]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[11],stage1_63[14],stage1_62[15],stage1_61[18]}
   );
   gpc606_5 gpc242 (
      {stage0_61[42], stage0_61[43], stage0_61[44], stage0_61[45], stage0_61[46], stage0_61[47]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[12],stage1_63[15],stage1_62[16],stage1_61[19]}
   );
   gpc606_5 gpc243 (
      {stage0_61[48], stage0_61[49], stage0_61[50], stage0_61[51], stage0_61[52], stage0_61[53]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[13],stage1_63[16],stage1_62[17],stage1_61[20]}
   );
   gpc1_1 gpc244 (
      {stage0_0[46]},
      {stage1_0[9]}
   );
   gpc1_1 gpc245 (
      {stage0_0[47]},
      {stage1_0[10]}
   );
   gpc1_1 gpc246 (
      {stage0_0[48]},
      {stage1_0[11]}
   );
   gpc1_1 gpc247 (
      {stage0_0[49]},
      {stage1_0[12]}
   );
   gpc1_1 gpc248 (
      {stage0_0[50]},
      {stage1_0[13]}
   );
   gpc1_1 gpc249 (
      {stage0_0[51]},
      {stage1_0[14]}
   );
   gpc1_1 gpc250 (
      {stage0_0[52]},
      {stage1_0[15]}
   );
   gpc1_1 gpc251 (
      {stage0_0[53]},
      {stage1_0[16]}
   );
   gpc1_1 gpc252 (
      {stage0_1[48]},
      {stage1_1[14]}
   );
   gpc1_1 gpc253 (
      {stage0_1[49]},
      {stage1_1[15]}
   );
   gpc1_1 gpc254 (
      {stage0_1[50]},
      {stage1_1[16]}
   );
   gpc1_1 gpc255 (
      {stage0_1[51]},
      {stage1_1[17]}
   );
   gpc1_1 gpc256 (
      {stage0_1[52]},
      {stage1_1[18]}
   );
   gpc1_1 gpc257 (
      {stage0_1[53]},
      {stage1_1[19]}
   );
   gpc1_1 gpc258 (
      {stage0_2[45]},
      {stage1_2[16]}
   );
   gpc1_1 gpc259 (
      {stage0_2[46]},
      {stage1_2[17]}
   );
   gpc1_1 gpc260 (
      {stage0_2[47]},
      {stage1_2[18]}
   );
   gpc1_1 gpc261 (
      {stage0_2[48]},
      {stage1_2[19]}
   );
   gpc1_1 gpc262 (
      {stage0_2[49]},
      {stage1_2[20]}
   );
   gpc1_1 gpc263 (
      {stage0_2[50]},
      {stage1_2[21]}
   );
   gpc1_1 gpc264 (
      {stage0_2[51]},
      {stage1_2[22]}
   );
   gpc1_1 gpc265 (
      {stage0_2[52]},
      {stage1_2[23]}
   );
   gpc1_1 gpc266 (
      {stage0_2[53]},
      {stage1_2[24]}
   );
   gpc1_1 gpc267 (
      {stage0_3[48]},
      {stage1_3[18]}
   );
   gpc1_1 gpc268 (
      {stage0_3[49]},
      {stage1_3[19]}
   );
   gpc1_1 gpc269 (
      {stage0_3[50]},
      {stage1_3[20]}
   );
   gpc1_1 gpc270 (
      {stage0_3[51]},
      {stage1_3[21]}
   );
   gpc1_1 gpc271 (
      {stage0_3[52]},
      {stage1_3[22]}
   );
   gpc1_1 gpc272 (
      {stage0_3[53]},
      {stage1_3[23]}
   );
   gpc1_1 gpc273 (
      {stage0_4[45]},
      {stage1_4[24]}
   );
   gpc1_1 gpc274 (
      {stage0_4[46]},
      {stage1_4[25]}
   );
   gpc1_1 gpc275 (
      {stage0_4[47]},
      {stage1_4[26]}
   );
   gpc1_1 gpc276 (
      {stage0_4[48]},
      {stage1_4[27]}
   );
   gpc1_1 gpc277 (
      {stage0_4[49]},
      {stage1_4[28]}
   );
   gpc1_1 gpc278 (
      {stage0_4[50]},
      {stage1_4[29]}
   );
   gpc1_1 gpc279 (
      {stage0_4[51]},
      {stage1_4[30]}
   );
   gpc1_1 gpc280 (
      {stage0_4[52]},
      {stage1_4[31]}
   );
   gpc1_1 gpc281 (
      {stage0_4[53]},
      {stage1_4[32]}
   );
   gpc1_1 gpc282 (
      {stage0_5[36]},
      {stage1_5[18]}
   );
   gpc1_1 gpc283 (
      {stage0_5[37]},
      {stage1_5[19]}
   );
   gpc1_1 gpc284 (
      {stage0_5[38]},
      {stage1_5[20]}
   );
   gpc1_1 gpc285 (
      {stage0_5[39]},
      {stage1_5[21]}
   );
   gpc1_1 gpc286 (
      {stage0_5[40]},
      {stage1_5[22]}
   );
   gpc1_1 gpc287 (
      {stage0_5[41]},
      {stage1_5[23]}
   );
   gpc1_1 gpc288 (
      {stage0_5[42]},
      {stage1_5[24]}
   );
   gpc1_1 gpc289 (
      {stage0_5[43]},
      {stage1_5[25]}
   );
   gpc1_1 gpc290 (
      {stage0_5[44]},
      {stage1_5[26]}
   );
   gpc1_1 gpc291 (
      {stage0_5[45]},
      {stage1_5[27]}
   );
   gpc1_1 gpc292 (
      {stage0_5[46]},
      {stage1_5[28]}
   );
   gpc1_1 gpc293 (
      {stage0_5[47]},
      {stage1_5[29]}
   );
   gpc1_1 gpc294 (
      {stage0_5[48]},
      {stage1_5[30]}
   );
   gpc1_1 gpc295 (
      {stage0_5[49]},
      {stage1_5[31]}
   );
   gpc1_1 gpc296 (
      {stage0_5[50]},
      {stage1_5[32]}
   );
   gpc1_1 gpc297 (
      {stage0_5[51]},
      {stage1_5[33]}
   );
   gpc1_1 gpc298 (
      {stage0_5[52]},
      {stage1_5[34]}
   );
   gpc1_1 gpc299 (
      {stage0_5[53]},
      {stage1_5[35]}
   );
   gpc1_1 gpc300 (
      {stage0_6[51]},
      {stage1_6[16]}
   );
   gpc1_1 gpc301 (
      {stage0_6[52]},
      {stage1_6[17]}
   );
   gpc1_1 gpc302 (
      {stage0_6[53]},
      {stage1_6[18]}
   );
   gpc1_1 gpc303 (
      {stage0_7[49]},
      {stage1_7[20]}
   );
   gpc1_1 gpc304 (
      {stage0_7[50]},
      {stage1_7[21]}
   );
   gpc1_1 gpc305 (
      {stage0_7[51]},
      {stage1_7[22]}
   );
   gpc1_1 gpc306 (
      {stage0_7[52]},
      {stage1_7[23]}
   );
   gpc1_1 gpc307 (
      {stage0_7[53]},
      {stage1_7[24]}
   );
   gpc1_1 gpc308 (
      {stage0_8[44]},
      {stage1_8[21]}
   );
   gpc1_1 gpc309 (
      {stage0_8[45]},
      {stage1_8[22]}
   );
   gpc1_1 gpc310 (
      {stage0_8[46]},
      {stage1_8[23]}
   );
   gpc1_1 gpc311 (
      {stage0_8[47]},
      {stage1_8[24]}
   );
   gpc1_1 gpc312 (
      {stage0_8[48]},
      {stage1_8[25]}
   );
   gpc1_1 gpc313 (
      {stage0_8[49]},
      {stage1_8[26]}
   );
   gpc1_1 gpc314 (
      {stage0_8[50]},
      {stage1_8[27]}
   );
   gpc1_1 gpc315 (
      {stage0_8[51]},
      {stage1_8[28]}
   );
   gpc1_1 gpc316 (
      {stage0_8[52]},
      {stage1_8[29]}
   );
   gpc1_1 gpc317 (
      {stage0_8[53]},
      {stage1_8[30]}
   );
   gpc1_1 gpc318 (
      {stage0_10[49]},
      {stage1_10[21]}
   );
   gpc1_1 gpc319 (
      {stage0_10[50]},
      {stage1_10[22]}
   );
   gpc1_1 gpc320 (
      {stage0_10[51]},
      {stage1_10[23]}
   );
   gpc1_1 gpc321 (
      {stage0_10[52]},
      {stage1_10[24]}
   );
   gpc1_1 gpc322 (
      {stage0_10[53]},
      {stage1_10[25]}
   );
   gpc1_1 gpc323 (
      {stage0_11[48]},
      {stage1_11[23]}
   );
   gpc1_1 gpc324 (
      {stage0_11[49]},
      {stage1_11[24]}
   );
   gpc1_1 gpc325 (
      {stage0_11[50]},
      {stage1_11[25]}
   );
   gpc1_1 gpc326 (
      {stage0_11[51]},
      {stage1_11[26]}
   );
   gpc1_1 gpc327 (
      {stage0_11[52]},
      {stage1_11[27]}
   );
   gpc1_1 gpc328 (
      {stage0_11[53]},
      {stage1_11[28]}
   );
   gpc1_1 gpc329 (
      {stage0_12[53]},
      {stage1_12[20]}
   );
   gpc1_1 gpc330 (
      {stage0_13[42]},
      {stage1_13[18]}
   );
   gpc1_1 gpc331 (
      {stage0_13[43]},
      {stage1_13[19]}
   );
   gpc1_1 gpc332 (
      {stage0_13[44]},
      {stage1_13[20]}
   );
   gpc1_1 gpc333 (
      {stage0_13[45]},
      {stage1_13[21]}
   );
   gpc1_1 gpc334 (
      {stage0_13[46]},
      {stage1_13[22]}
   );
   gpc1_1 gpc335 (
      {stage0_13[47]},
      {stage1_13[23]}
   );
   gpc1_1 gpc336 (
      {stage0_13[48]},
      {stage1_13[24]}
   );
   gpc1_1 gpc337 (
      {stage0_13[49]},
      {stage1_13[25]}
   );
   gpc1_1 gpc338 (
      {stage0_13[50]},
      {stage1_13[26]}
   );
   gpc1_1 gpc339 (
      {stage0_13[51]},
      {stage1_13[27]}
   );
   gpc1_1 gpc340 (
      {stage0_13[52]},
      {stage1_13[28]}
   );
   gpc1_1 gpc341 (
      {stage0_13[53]},
      {stage1_13[29]}
   );
   gpc1_1 gpc342 (
      {stage0_14[51]},
      {stage1_14[21]}
   );
   gpc1_1 gpc343 (
      {stage0_14[52]},
      {stage1_14[22]}
   );
   gpc1_1 gpc344 (
      {stage0_14[53]},
      {stage1_14[23]}
   );
   gpc1_1 gpc345 (
      {stage0_15[30]},
      {stage1_15[19]}
   );
   gpc1_1 gpc346 (
      {stage0_15[31]},
      {stage1_15[20]}
   );
   gpc1_1 gpc347 (
      {stage0_15[32]},
      {stage1_15[21]}
   );
   gpc1_1 gpc348 (
      {stage0_15[33]},
      {stage1_15[22]}
   );
   gpc1_1 gpc349 (
      {stage0_15[34]},
      {stage1_15[23]}
   );
   gpc1_1 gpc350 (
      {stage0_15[35]},
      {stage1_15[24]}
   );
   gpc1_1 gpc351 (
      {stage0_15[36]},
      {stage1_15[25]}
   );
   gpc1_1 gpc352 (
      {stage0_15[37]},
      {stage1_15[26]}
   );
   gpc1_1 gpc353 (
      {stage0_15[38]},
      {stage1_15[27]}
   );
   gpc1_1 gpc354 (
      {stage0_15[39]},
      {stage1_15[28]}
   );
   gpc1_1 gpc355 (
      {stage0_15[40]},
      {stage1_15[29]}
   );
   gpc1_1 gpc356 (
      {stage0_15[41]},
      {stage1_15[30]}
   );
   gpc1_1 gpc357 (
      {stage0_15[42]},
      {stage1_15[31]}
   );
   gpc1_1 gpc358 (
      {stage0_15[43]},
      {stage1_15[32]}
   );
   gpc1_1 gpc359 (
      {stage0_15[44]},
      {stage1_15[33]}
   );
   gpc1_1 gpc360 (
      {stage0_15[45]},
      {stage1_15[34]}
   );
   gpc1_1 gpc361 (
      {stage0_15[46]},
      {stage1_15[35]}
   );
   gpc1_1 gpc362 (
      {stage0_15[47]},
      {stage1_15[36]}
   );
   gpc1_1 gpc363 (
      {stage0_15[48]},
      {stage1_15[37]}
   );
   gpc1_1 gpc364 (
      {stage0_15[49]},
      {stage1_15[38]}
   );
   gpc1_1 gpc365 (
      {stage0_15[50]},
      {stage1_15[39]}
   );
   gpc1_1 gpc366 (
      {stage0_15[51]},
      {stage1_15[40]}
   );
   gpc1_1 gpc367 (
      {stage0_15[52]},
      {stage1_15[41]}
   );
   gpc1_1 gpc368 (
      {stage0_15[53]},
      {stage1_15[42]}
   );
   gpc1_1 gpc369 (
      {stage0_16[45]},
      {stage1_16[15]}
   );
   gpc1_1 gpc370 (
      {stage0_16[46]},
      {stage1_16[16]}
   );
   gpc1_1 gpc371 (
      {stage0_16[47]},
      {stage1_16[17]}
   );
   gpc1_1 gpc372 (
      {stage0_16[48]},
      {stage1_16[18]}
   );
   gpc1_1 gpc373 (
      {stage0_16[49]},
      {stage1_16[19]}
   );
   gpc1_1 gpc374 (
      {stage0_16[50]},
      {stage1_16[20]}
   );
   gpc1_1 gpc375 (
      {stage0_16[51]},
      {stage1_16[21]}
   );
   gpc1_1 gpc376 (
      {stage0_16[52]},
      {stage1_16[22]}
   );
   gpc1_1 gpc377 (
      {stage0_16[53]},
      {stage1_16[23]}
   );
   gpc1_1 gpc378 (
      {stage0_18[42]},
      {stage1_18[22]}
   );
   gpc1_1 gpc379 (
      {stage0_18[43]},
      {stage1_18[23]}
   );
   gpc1_1 gpc380 (
      {stage0_18[44]},
      {stage1_18[24]}
   );
   gpc1_1 gpc381 (
      {stage0_18[45]},
      {stage1_18[25]}
   );
   gpc1_1 gpc382 (
      {stage0_18[46]},
      {stage1_18[26]}
   );
   gpc1_1 gpc383 (
      {stage0_18[47]},
      {stage1_18[27]}
   );
   gpc1_1 gpc384 (
      {stage0_18[48]},
      {stage1_18[28]}
   );
   gpc1_1 gpc385 (
      {stage0_18[49]},
      {stage1_18[29]}
   );
   gpc1_1 gpc386 (
      {stage0_18[50]},
      {stage1_18[30]}
   );
   gpc1_1 gpc387 (
      {stage0_18[51]},
      {stage1_18[31]}
   );
   gpc1_1 gpc388 (
      {stage0_18[52]},
      {stage1_18[32]}
   );
   gpc1_1 gpc389 (
      {stage0_18[53]},
      {stage1_18[33]}
   );
   gpc1_1 gpc390 (
      {stage0_19[52]},
      {stage1_19[19]}
   );
   gpc1_1 gpc391 (
      {stage0_19[53]},
      {stage1_19[20]}
   );
   gpc1_1 gpc392 (
      {stage0_20[53]},
      {stage1_20[19]}
   );
   gpc1_1 gpc393 (
      {stage0_21[51]},
      {stage1_21[23]}
   );
   gpc1_1 gpc394 (
      {stage0_21[52]},
      {stage1_21[24]}
   );
   gpc1_1 gpc395 (
      {stage0_21[53]},
      {stage1_21[25]}
   );
   gpc1_1 gpc396 (
      {stage0_24[41]},
      {stage1_24[19]}
   );
   gpc1_1 gpc397 (
      {stage0_24[42]},
      {stage1_24[20]}
   );
   gpc1_1 gpc398 (
      {stage0_24[43]},
      {stage1_24[21]}
   );
   gpc1_1 gpc399 (
      {stage0_24[44]},
      {stage1_24[22]}
   );
   gpc1_1 gpc400 (
      {stage0_24[45]},
      {stage1_24[23]}
   );
   gpc1_1 gpc401 (
      {stage0_24[46]},
      {stage1_24[24]}
   );
   gpc1_1 gpc402 (
      {stage0_24[47]},
      {stage1_24[25]}
   );
   gpc1_1 gpc403 (
      {stage0_24[48]},
      {stage1_24[26]}
   );
   gpc1_1 gpc404 (
      {stage0_24[49]},
      {stage1_24[27]}
   );
   gpc1_1 gpc405 (
      {stage0_24[50]},
      {stage1_24[28]}
   );
   gpc1_1 gpc406 (
      {stage0_24[51]},
      {stage1_24[29]}
   );
   gpc1_1 gpc407 (
      {stage0_24[52]},
      {stage1_24[30]}
   );
   gpc1_1 gpc408 (
      {stage0_24[53]},
      {stage1_24[31]}
   );
   gpc1_1 gpc409 (
      {stage0_25[48]},
      {stage1_25[19]}
   );
   gpc1_1 gpc410 (
      {stage0_25[49]},
      {stage1_25[20]}
   );
   gpc1_1 gpc411 (
      {stage0_25[50]},
      {stage1_25[21]}
   );
   gpc1_1 gpc412 (
      {stage0_25[51]},
      {stage1_25[22]}
   );
   gpc1_1 gpc413 (
      {stage0_25[52]},
      {stage1_25[23]}
   );
   gpc1_1 gpc414 (
      {stage0_25[53]},
      {stage1_25[24]}
   );
   gpc1_1 gpc415 (
      {stage0_26[45]},
      {stage1_26[23]}
   );
   gpc1_1 gpc416 (
      {stage0_26[46]},
      {stage1_26[24]}
   );
   gpc1_1 gpc417 (
      {stage0_26[47]},
      {stage1_26[25]}
   );
   gpc1_1 gpc418 (
      {stage0_26[48]},
      {stage1_26[26]}
   );
   gpc1_1 gpc419 (
      {stage0_26[49]},
      {stage1_26[27]}
   );
   gpc1_1 gpc420 (
      {stage0_26[50]},
      {stage1_26[28]}
   );
   gpc1_1 gpc421 (
      {stage0_26[51]},
      {stage1_26[29]}
   );
   gpc1_1 gpc422 (
      {stage0_26[52]},
      {stage1_26[30]}
   );
   gpc1_1 gpc423 (
      {stage0_26[53]},
      {stage1_26[31]}
   );
   gpc1_1 gpc424 (
      {stage0_27[50]},
      {stage1_27[20]}
   );
   gpc1_1 gpc425 (
      {stage0_27[51]},
      {stage1_27[21]}
   );
   gpc1_1 gpc426 (
      {stage0_27[52]},
      {stage1_27[22]}
   );
   gpc1_1 gpc427 (
      {stage0_27[53]},
      {stage1_27[23]}
   );
   gpc1_1 gpc428 (
      {stage0_29[50]},
      {stage1_29[22]}
   );
   gpc1_1 gpc429 (
      {stage0_29[51]},
      {stage1_29[23]}
   );
   gpc1_1 gpc430 (
      {stage0_29[52]},
      {stage1_29[24]}
   );
   gpc1_1 gpc431 (
      {stage0_29[53]},
      {stage1_29[25]}
   );
   gpc1_1 gpc432 (
      {stage0_30[42]},
      {stage1_30[23]}
   );
   gpc1_1 gpc433 (
      {stage0_30[43]},
      {stage1_30[24]}
   );
   gpc1_1 gpc434 (
      {stage0_30[44]},
      {stage1_30[25]}
   );
   gpc1_1 gpc435 (
      {stage0_30[45]},
      {stage1_30[26]}
   );
   gpc1_1 gpc436 (
      {stage0_30[46]},
      {stage1_30[27]}
   );
   gpc1_1 gpc437 (
      {stage0_30[47]},
      {stage1_30[28]}
   );
   gpc1_1 gpc438 (
      {stage0_30[48]},
      {stage1_30[29]}
   );
   gpc1_1 gpc439 (
      {stage0_30[49]},
      {stage1_30[30]}
   );
   gpc1_1 gpc440 (
      {stage0_30[50]},
      {stage1_30[31]}
   );
   gpc1_1 gpc441 (
      {stage0_30[51]},
      {stage1_30[32]}
   );
   gpc1_1 gpc442 (
      {stage0_30[52]},
      {stage1_30[33]}
   );
   gpc1_1 gpc443 (
      {stage0_30[53]},
      {stage1_30[34]}
   );
   gpc1_1 gpc444 (
      {stage0_31[36]},
      {stage1_31[16]}
   );
   gpc1_1 gpc445 (
      {stage0_31[37]},
      {stage1_31[17]}
   );
   gpc1_1 gpc446 (
      {stage0_31[38]},
      {stage1_31[18]}
   );
   gpc1_1 gpc447 (
      {stage0_31[39]},
      {stage1_31[19]}
   );
   gpc1_1 gpc448 (
      {stage0_31[40]},
      {stage1_31[20]}
   );
   gpc1_1 gpc449 (
      {stage0_31[41]},
      {stage1_31[21]}
   );
   gpc1_1 gpc450 (
      {stage0_31[42]},
      {stage1_31[22]}
   );
   gpc1_1 gpc451 (
      {stage0_31[43]},
      {stage1_31[23]}
   );
   gpc1_1 gpc452 (
      {stage0_31[44]},
      {stage1_31[24]}
   );
   gpc1_1 gpc453 (
      {stage0_31[45]},
      {stage1_31[25]}
   );
   gpc1_1 gpc454 (
      {stage0_31[46]},
      {stage1_31[26]}
   );
   gpc1_1 gpc455 (
      {stage0_31[47]},
      {stage1_31[27]}
   );
   gpc1_1 gpc456 (
      {stage0_31[48]},
      {stage1_31[28]}
   );
   gpc1_1 gpc457 (
      {stage0_31[49]},
      {stage1_31[29]}
   );
   gpc1_1 gpc458 (
      {stage0_31[50]},
      {stage1_31[30]}
   );
   gpc1_1 gpc459 (
      {stage0_31[51]},
      {stage1_31[31]}
   );
   gpc1_1 gpc460 (
      {stage0_31[52]},
      {stage1_31[32]}
   );
   gpc1_1 gpc461 (
      {stage0_31[53]},
      {stage1_31[33]}
   );
   gpc1_1 gpc462 (
      {stage0_32[53]},
      {stage1_32[18]}
   );
   gpc1_1 gpc463 (
      {stage0_33[25]},
      {stage1_33[17]}
   );
   gpc1_1 gpc464 (
      {stage0_33[26]},
      {stage1_33[18]}
   );
   gpc1_1 gpc465 (
      {stage0_33[27]},
      {stage1_33[19]}
   );
   gpc1_1 gpc466 (
      {stage0_33[28]},
      {stage1_33[20]}
   );
   gpc1_1 gpc467 (
      {stage0_33[29]},
      {stage1_33[21]}
   );
   gpc1_1 gpc468 (
      {stage0_33[30]},
      {stage1_33[22]}
   );
   gpc1_1 gpc469 (
      {stage0_33[31]},
      {stage1_33[23]}
   );
   gpc1_1 gpc470 (
      {stage0_33[32]},
      {stage1_33[24]}
   );
   gpc1_1 gpc471 (
      {stage0_33[33]},
      {stage1_33[25]}
   );
   gpc1_1 gpc472 (
      {stage0_33[34]},
      {stage1_33[26]}
   );
   gpc1_1 gpc473 (
      {stage0_33[35]},
      {stage1_33[27]}
   );
   gpc1_1 gpc474 (
      {stage0_33[36]},
      {stage1_33[28]}
   );
   gpc1_1 gpc475 (
      {stage0_33[37]},
      {stage1_33[29]}
   );
   gpc1_1 gpc476 (
      {stage0_33[38]},
      {stage1_33[30]}
   );
   gpc1_1 gpc477 (
      {stage0_33[39]},
      {stage1_33[31]}
   );
   gpc1_1 gpc478 (
      {stage0_33[40]},
      {stage1_33[32]}
   );
   gpc1_1 gpc479 (
      {stage0_33[41]},
      {stage1_33[33]}
   );
   gpc1_1 gpc480 (
      {stage0_33[42]},
      {stage1_33[34]}
   );
   gpc1_1 gpc481 (
      {stage0_33[43]},
      {stage1_33[35]}
   );
   gpc1_1 gpc482 (
      {stage0_33[44]},
      {stage1_33[36]}
   );
   gpc1_1 gpc483 (
      {stage0_33[45]},
      {stage1_33[37]}
   );
   gpc1_1 gpc484 (
      {stage0_33[46]},
      {stage1_33[38]}
   );
   gpc1_1 gpc485 (
      {stage0_33[47]},
      {stage1_33[39]}
   );
   gpc1_1 gpc486 (
      {stage0_33[48]},
      {stage1_33[40]}
   );
   gpc1_1 gpc487 (
      {stage0_33[49]},
      {stage1_33[41]}
   );
   gpc1_1 gpc488 (
      {stage0_33[50]},
      {stage1_33[42]}
   );
   gpc1_1 gpc489 (
      {stage0_33[51]},
      {stage1_33[43]}
   );
   gpc1_1 gpc490 (
      {stage0_33[52]},
      {stage1_33[44]}
   );
   gpc1_1 gpc491 (
      {stage0_33[53]},
      {stage1_33[45]}
   );
   gpc1_1 gpc492 (
      {stage0_34[51]},
      {stage1_34[16]}
   );
   gpc1_1 gpc493 (
      {stage0_34[52]},
      {stage1_34[17]}
   );
   gpc1_1 gpc494 (
      {stage0_34[53]},
      {stage1_34[18]}
   );
   gpc1_1 gpc495 (
      {stage0_35[43]},
      {stage1_35[17]}
   );
   gpc1_1 gpc496 (
      {stage0_35[44]},
      {stage1_35[18]}
   );
   gpc1_1 gpc497 (
      {stage0_35[45]},
      {stage1_35[19]}
   );
   gpc1_1 gpc498 (
      {stage0_35[46]},
      {stage1_35[20]}
   );
   gpc1_1 gpc499 (
      {stage0_35[47]},
      {stage1_35[21]}
   );
   gpc1_1 gpc500 (
      {stage0_35[48]},
      {stage1_35[22]}
   );
   gpc1_1 gpc501 (
      {stage0_35[49]},
      {stage1_35[23]}
   );
   gpc1_1 gpc502 (
      {stage0_35[50]},
      {stage1_35[24]}
   );
   gpc1_1 gpc503 (
      {stage0_35[51]},
      {stage1_35[25]}
   );
   gpc1_1 gpc504 (
      {stage0_35[52]},
      {stage1_35[26]}
   );
   gpc1_1 gpc505 (
      {stage0_35[53]},
      {stage1_35[27]}
   );
   gpc1_1 gpc506 (
      {stage0_36[41]},
      {stage1_36[21]}
   );
   gpc1_1 gpc507 (
      {stage0_36[42]},
      {stage1_36[22]}
   );
   gpc1_1 gpc508 (
      {stage0_36[43]},
      {stage1_36[23]}
   );
   gpc1_1 gpc509 (
      {stage0_36[44]},
      {stage1_36[24]}
   );
   gpc1_1 gpc510 (
      {stage0_36[45]},
      {stage1_36[25]}
   );
   gpc1_1 gpc511 (
      {stage0_36[46]},
      {stage1_36[26]}
   );
   gpc1_1 gpc512 (
      {stage0_36[47]},
      {stage1_36[27]}
   );
   gpc1_1 gpc513 (
      {stage0_36[48]},
      {stage1_36[28]}
   );
   gpc1_1 gpc514 (
      {stage0_36[49]},
      {stage1_36[29]}
   );
   gpc1_1 gpc515 (
      {stage0_36[50]},
      {stage1_36[30]}
   );
   gpc1_1 gpc516 (
      {stage0_36[51]},
      {stage1_36[31]}
   );
   gpc1_1 gpc517 (
      {stage0_36[52]},
      {stage1_36[32]}
   );
   gpc1_1 gpc518 (
      {stage0_36[53]},
      {stage1_36[33]}
   );
   gpc1_1 gpc519 (
      {stage0_37[48]},
      {stage1_37[19]}
   );
   gpc1_1 gpc520 (
      {stage0_37[49]},
      {stage1_37[20]}
   );
   gpc1_1 gpc521 (
      {stage0_37[50]},
      {stage1_37[21]}
   );
   gpc1_1 gpc522 (
      {stage0_37[51]},
      {stage1_37[22]}
   );
   gpc1_1 gpc523 (
      {stage0_37[52]},
      {stage1_37[23]}
   );
   gpc1_1 gpc524 (
      {stage0_37[53]},
      {stage1_37[24]}
   );
   gpc1_1 gpc525 (
      {stage0_38[46]},
      {stage1_38[16]}
   );
   gpc1_1 gpc526 (
      {stage0_38[47]},
      {stage1_38[17]}
   );
   gpc1_1 gpc527 (
      {stage0_38[48]},
      {stage1_38[18]}
   );
   gpc1_1 gpc528 (
      {stage0_38[49]},
      {stage1_38[19]}
   );
   gpc1_1 gpc529 (
      {stage0_38[50]},
      {stage1_38[20]}
   );
   gpc1_1 gpc530 (
      {stage0_38[51]},
      {stage1_38[21]}
   );
   gpc1_1 gpc531 (
      {stage0_38[52]},
      {stage1_38[22]}
   );
   gpc1_1 gpc532 (
      {stage0_38[53]},
      {stage1_38[23]}
   );
   gpc1_1 gpc533 (
      {stage0_39[43]},
      {stage1_39[20]}
   );
   gpc1_1 gpc534 (
      {stage0_39[44]},
      {stage1_39[21]}
   );
   gpc1_1 gpc535 (
      {stage0_39[45]},
      {stage1_39[22]}
   );
   gpc1_1 gpc536 (
      {stage0_39[46]},
      {stage1_39[23]}
   );
   gpc1_1 gpc537 (
      {stage0_39[47]},
      {stage1_39[24]}
   );
   gpc1_1 gpc538 (
      {stage0_39[48]},
      {stage1_39[25]}
   );
   gpc1_1 gpc539 (
      {stage0_39[49]},
      {stage1_39[26]}
   );
   gpc1_1 gpc540 (
      {stage0_39[50]},
      {stage1_39[27]}
   );
   gpc1_1 gpc541 (
      {stage0_39[51]},
      {stage1_39[28]}
   );
   gpc1_1 gpc542 (
      {stage0_39[52]},
      {stage1_39[29]}
   );
   gpc1_1 gpc543 (
      {stage0_39[53]},
      {stage1_39[30]}
   );
   gpc1_1 gpc544 (
      {stage0_40[34]},
      {stage1_40[19]}
   );
   gpc1_1 gpc545 (
      {stage0_40[35]},
      {stage1_40[20]}
   );
   gpc1_1 gpc546 (
      {stage0_40[36]},
      {stage1_40[21]}
   );
   gpc1_1 gpc547 (
      {stage0_40[37]},
      {stage1_40[22]}
   );
   gpc1_1 gpc548 (
      {stage0_40[38]},
      {stage1_40[23]}
   );
   gpc1_1 gpc549 (
      {stage0_40[39]},
      {stage1_40[24]}
   );
   gpc1_1 gpc550 (
      {stage0_40[40]},
      {stage1_40[25]}
   );
   gpc1_1 gpc551 (
      {stage0_40[41]},
      {stage1_40[26]}
   );
   gpc1_1 gpc552 (
      {stage0_40[42]},
      {stage1_40[27]}
   );
   gpc1_1 gpc553 (
      {stage0_40[43]},
      {stage1_40[28]}
   );
   gpc1_1 gpc554 (
      {stage0_40[44]},
      {stage1_40[29]}
   );
   gpc1_1 gpc555 (
      {stage0_40[45]},
      {stage1_40[30]}
   );
   gpc1_1 gpc556 (
      {stage0_40[46]},
      {stage1_40[31]}
   );
   gpc1_1 gpc557 (
      {stage0_40[47]},
      {stage1_40[32]}
   );
   gpc1_1 gpc558 (
      {stage0_40[48]},
      {stage1_40[33]}
   );
   gpc1_1 gpc559 (
      {stage0_40[49]},
      {stage1_40[34]}
   );
   gpc1_1 gpc560 (
      {stage0_40[50]},
      {stage1_40[35]}
   );
   gpc1_1 gpc561 (
      {stage0_40[51]},
      {stage1_40[36]}
   );
   gpc1_1 gpc562 (
      {stage0_40[52]},
      {stage1_40[37]}
   );
   gpc1_1 gpc563 (
      {stage0_40[53]},
      {stage1_40[38]}
   );
   gpc1_1 gpc564 (
      {stage0_41[51]},
      {stage1_41[17]}
   );
   gpc1_1 gpc565 (
      {stage0_41[52]},
      {stage1_41[18]}
   );
   gpc1_1 gpc566 (
      {stage0_41[53]},
      {stage1_41[19]}
   );
   gpc1_1 gpc567 (
      {stage0_42[52]},
      {stage1_42[19]}
   );
   gpc1_1 gpc568 (
      {stage0_42[53]},
      {stage1_42[20]}
   );
   gpc1_1 gpc569 (
      {stage0_45[41]},
      {stage1_45[19]}
   );
   gpc1_1 gpc570 (
      {stage0_45[42]},
      {stage1_45[20]}
   );
   gpc1_1 gpc571 (
      {stage0_45[43]},
      {stage1_45[21]}
   );
   gpc1_1 gpc572 (
      {stage0_45[44]},
      {stage1_45[22]}
   );
   gpc1_1 gpc573 (
      {stage0_45[45]},
      {stage1_45[23]}
   );
   gpc1_1 gpc574 (
      {stage0_45[46]},
      {stage1_45[24]}
   );
   gpc1_1 gpc575 (
      {stage0_45[47]},
      {stage1_45[25]}
   );
   gpc1_1 gpc576 (
      {stage0_45[48]},
      {stage1_45[26]}
   );
   gpc1_1 gpc577 (
      {stage0_45[49]},
      {stage1_45[27]}
   );
   gpc1_1 gpc578 (
      {stage0_45[50]},
      {stage1_45[28]}
   );
   gpc1_1 gpc579 (
      {stage0_45[51]},
      {stage1_45[29]}
   );
   gpc1_1 gpc580 (
      {stage0_45[52]},
      {stage1_45[30]}
   );
   gpc1_1 gpc581 (
      {stage0_45[53]},
      {stage1_45[31]}
   );
   gpc1_1 gpc582 (
      {stage0_46[44]},
      {stage1_46[20]}
   );
   gpc1_1 gpc583 (
      {stage0_46[45]},
      {stage1_46[21]}
   );
   gpc1_1 gpc584 (
      {stage0_46[46]},
      {stage1_46[22]}
   );
   gpc1_1 gpc585 (
      {stage0_46[47]},
      {stage1_46[23]}
   );
   gpc1_1 gpc586 (
      {stage0_46[48]},
      {stage1_46[24]}
   );
   gpc1_1 gpc587 (
      {stage0_46[49]},
      {stage1_46[25]}
   );
   gpc1_1 gpc588 (
      {stage0_46[50]},
      {stage1_46[26]}
   );
   gpc1_1 gpc589 (
      {stage0_46[51]},
      {stage1_46[27]}
   );
   gpc1_1 gpc590 (
      {stage0_46[52]},
      {stage1_46[28]}
   );
   gpc1_1 gpc591 (
      {stage0_46[53]},
      {stage1_46[29]}
   );
   gpc1_1 gpc592 (
      {stage0_47[41]},
      {stage1_47[21]}
   );
   gpc1_1 gpc593 (
      {stage0_47[42]},
      {stage1_47[22]}
   );
   gpc1_1 gpc594 (
      {stage0_47[43]},
      {stage1_47[23]}
   );
   gpc1_1 gpc595 (
      {stage0_47[44]},
      {stage1_47[24]}
   );
   gpc1_1 gpc596 (
      {stage0_47[45]},
      {stage1_47[25]}
   );
   gpc1_1 gpc597 (
      {stage0_47[46]},
      {stage1_47[26]}
   );
   gpc1_1 gpc598 (
      {stage0_47[47]},
      {stage1_47[27]}
   );
   gpc1_1 gpc599 (
      {stage0_47[48]},
      {stage1_47[28]}
   );
   gpc1_1 gpc600 (
      {stage0_47[49]},
      {stage1_47[29]}
   );
   gpc1_1 gpc601 (
      {stage0_47[50]},
      {stage1_47[30]}
   );
   gpc1_1 gpc602 (
      {stage0_47[51]},
      {stage1_47[31]}
   );
   gpc1_1 gpc603 (
      {stage0_47[52]},
      {stage1_47[32]}
   );
   gpc1_1 gpc604 (
      {stage0_47[53]},
      {stage1_47[33]}
   );
   gpc1_1 gpc605 (
      {stage0_49[47]},
      {stage1_49[17]}
   );
   gpc1_1 gpc606 (
      {stage0_49[48]},
      {stage1_49[18]}
   );
   gpc1_1 gpc607 (
      {stage0_49[49]},
      {stage1_49[19]}
   );
   gpc1_1 gpc608 (
      {stage0_49[50]},
      {stage1_49[20]}
   );
   gpc1_1 gpc609 (
      {stage0_49[51]},
      {stage1_49[21]}
   );
   gpc1_1 gpc610 (
      {stage0_49[52]},
      {stage1_49[22]}
   );
   gpc1_1 gpc611 (
      {stage0_49[53]},
      {stage1_49[23]}
   );
   gpc1_1 gpc612 (
      {stage0_50[29]},
      {stage1_50[18]}
   );
   gpc1_1 gpc613 (
      {stage0_50[30]},
      {stage1_50[19]}
   );
   gpc1_1 gpc614 (
      {stage0_50[31]},
      {stage1_50[20]}
   );
   gpc1_1 gpc615 (
      {stage0_50[32]},
      {stage1_50[21]}
   );
   gpc1_1 gpc616 (
      {stage0_50[33]},
      {stage1_50[22]}
   );
   gpc1_1 gpc617 (
      {stage0_50[34]},
      {stage1_50[23]}
   );
   gpc1_1 gpc618 (
      {stage0_50[35]},
      {stage1_50[24]}
   );
   gpc1_1 gpc619 (
      {stage0_50[36]},
      {stage1_50[25]}
   );
   gpc1_1 gpc620 (
      {stage0_50[37]},
      {stage1_50[26]}
   );
   gpc1_1 gpc621 (
      {stage0_50[38]},
      {stage1_50[27]}
   );
   gpc1_1 gpc622 (
      {stage0_50[39]},
      {stage1_50[28]}
   );
   gpc1_1 gpc623 (
      {stage0_50[40]},
      {stage1_50[29]}
   );
   gpc1_1 gpc624 (
      {stage0_50[41]},
      {stage1_50[30]}
   );
   gpc1_1 gpc625 (
      {stage0_50[42]},
      {stage1_50[31]}
   );
   gpc1_1 gpc626 (
      {stage0_50[43]},
      {stage1_50[32]}
   );
   gpc1_1 gpc627 (
      {stage0_50[44]},
      {stage1_50[33]}
   );
   gpc1_1 gpc628 (
      {stage0_50[45]},
      {stage1_50[34]}
   );
   gpc1_1 gpc629 (
      {stage0_50[46]},
      {stage1_50[35]}
   );
   gpc1_1 gpc630 (
      {stage0_50[47]},
      {stage1_50[36]}
   );
   gpc1_1 gpc631 (
      {stage0_50[48]},
      {stage1_50[37]}
   );
   gpc1_1 gpc632 (
      {stage0_50[49]},
      {stage1_50[38]}
   );
   gpc1_1 gpc633 (
      {stage0_50[50]},
      {stage1_50[39]}
   );
   gpc1_1 gpc634 (
      {stage0_50[51]},
      {stage1_50[40]}
   );
   gpc1_1 gpc635 (
      {stage0_50[52]},
      {stage1_50[41]}
   );
   gpc1_1 gpc636 (
      {stage0_50[53]},
      {stage1_50[42]}
   );
   gpc1_1 gpc637 (
      {stage0_51[20]},
      {stage1_51[14]}
   );
   gpc1_1 gpc638 (
      {stage0_51[21]},
      {stage1_51[15]}
   );
   gpc1_1 gpc639 (
      {stage0_51[22]},
      {stage1_51[16]}
   );
   gpc1_1 gpc640 (
      {stage0_51[23]},
      {stage1_51[17]}
   );
   gpc1_1 gpc641 (
      {stage0_51[24]},
      {stage1_51[18]}
   );
   gpc1_1 gpc642 (
      {stage0_51[25]},
      {stage1_51[19]}
   );
   gpc1_1 gpc643 (
      {stage0_51[26]},
      {stage1_51[20]}
   );
   gpc1_1 gpc644 (
      {stage0_51[27]},
      {stage1_51[21]}
   );
   gpc1_1 gpc645 (
      {stage0_51[28]},
      {stage1_51[22]}
   );
   gpc1_1 gpc646 (
      {stage0_51[29]},
      {stage1_51[23]}
   );
   gpc1_1 gpc647 (
      {stage0_51[30]},
      {stage1_51[24]}
   );
   gpc1_1 gpc648 (
      {stage0_51[31]},
      {stage1_51[25]}
   );
   gpc1_1 gpc649 (
      {stage0_51[32]},
      {stage1_51[26]}
   );
   gpc1_1 gpc650 (
      {stage0_51[33]},
      {stage1_51[27]}
   );
   gpc1_1 gpc651 (
      {stage0_51[34]},
      {stage1_51[28]}
   );
   gpc1_1 gpc652 (
      {stage0_51[35]},
      {stage1_51[29]}
   );
   gpc1_1 gpc653 (
      {stage0_51[36]},
      {stage1_51[30]}
   );
   gpc1_1 gpc654 (
      {stage0_51[37]},
      {stage1_51[31]}
   );
   gpc1_1 gpc655 (
      {stage0_51[38]},
      {stage1_51[32]}
   );
   gpc1_1 gpc656 (
      {stage0_51[39]},
      {stage1_51[33]}
   );
   gpc1_1 gpc657 (
      {stage0_51[40]},
      {stage1_51[34]}
   );
   gpc1_1 gpc658 (
      {stage0_51[41]},
      {stage1_51[35]}
   );
   gpc1_1 gpc659 (
      {stage0_51[42]},
      {stage1_51[36]}
   );
   gpc1_1 gpc660 (
      {stage0_51[43]},
      {stage1_51[37]}
   );
   gpc1_1 gpc661 (
      {stage0_51[44]},
      {stage1_51[38]}
   );
   gpc1_1 gpc662 (
      {stage0_51[45]},
      {stage1_51[39]}
   );
   gpc1_1 gpc663 (
      {stage0_51[46]},
      {stage1_51[40]}
   );
   gpc1_1 gpc664 (
      {stage0_51[47]},
      {stage1_51[41]}
   );
   gpc1_1 gpc665 (
      {stage0_51[48]},
      {stage1_51[42]}
   );
   gpc1_1 gpc666 (
      {stage0_51[49]},
      {stage1_51[43]}
   );
   gpc1_1 gpc667 (
      {stage0_51[50]},
      {stage1_51[44]}
   );
   gpc1_1 gpc668 (
      {stage0_51[51]},
      {stage1_51[45]}
   );
   gpc1_1 gpc669 (
      {stage0_51[52]},
      {stage1_51[46]}
   );
   gpc1_1 gpc670 (
      {stage0_51[53]},
      {stage1_51[47]}
   );
   gpc1_1 gpc671 (
      {stage0_52[47]},
      {stage1_52[15]}
   );
   gpc1_1 gpc672 (
      {stage0_52[48]},
      {stage1_52[16]}
   );
   gpc1_1 gpc673 (
      {stage0_52[49]},
      {stage1_52[17]}
   );
   gpc1_1 gpc674 (
      {stage0_52[50]},
      {stage1_52[18]}
   );
   gpc1_1 gpc675 (
      {stage0_52[51]},
      {stage1_52[19]}
   );
   gpc1_1 gpc676 (
      {stage0_52[52]},
      {stage1_52[20]}
   );
   gpc1_1 gpc677 (
      {stage0_52[53]},
      {stage1_52[21]}
   );
   gpc1_1 gpc678 (
      {stage0_53[28]},
      {stage1_53[15]}
   );
   gpc1_1 gpc679 (
      {stage0_53[29]},
      {stage1_53[16]}
   );
   gpc1_1 gpc680 (
      {stage0_53[30]},
      {stage1_53[17]}
   );
   gpc1_1 gpc681 (
      {stage0_53[31]},
      {stage1_53[18]}
   );
   gpc1_1 gpc682 (
      {stage0_53[32]},
      {stage1_53[19]}
   );
   gpc1_1 gpc683 (
      {stage0_53[33]},
      {stage1_53[20]}
   );
   gpc1_1 gpc684 (
      {stage0_53[34]},
      {stage1_53[21]}
   );
   gpc1_1 gpc685 (
      {stage0_53[35]},
      {stage1_53[22]}
   );
   gpc1_1 gpc686 (
      {stage0_53[36]},
      {stage1_53[23]}
   );
   gpc1_1 gpc687 (
      {stage0_53[37]},
      {stage1_53[24]}
   );
   gpc1_1 gpc688 (
      {stage0_53[38]},
      {stage1_53[25]}
   );
   gpc1_1 gpc689 (
      {stage0_53[39]},
      {stage1_53[26]}
   );
   gpc1_1 gpc690 (
      {stage0_53[40]},
      {stage1_53[27]}
   );
   gpc1_1 gpc691 (
      {stage0_53[41]},
      {stage1_53[28]}
   );
   gpc1_1 gpc692 (
      {stage0_53[42]},
      {stage1_53[29]}
   );
   gpc1_1 gpc693 (
      {stage0_53[43]},
      {stage1_53[30]}
   );
   gpc1_1 gpc694 (
      {stage0_53[44]},
      {stage1_53[31]}
   );
   gpc1_1 gpc695 (
      {stage0_53[45]},
      {stage1_53[32]}
   );
   gpc1_1 gpc696 (
      {stage0_53[46]},
      {stage1_53[33]}
   );
   gpc1_1 gpc697 (
      {stage0_53[47]},
      {stage1_53[34]}
   );
   gpc1_1 gpc698 (
      {stage0_53[48]},
      {stage1_53[35]}
   );
   gpc1_1 gpc699 (
      {stage0_53[49]},
      {stage1_53[36]}
   );
   gpc1_1 gpc700 (
      {stage0_53[50]},
      {stage1_53[37]}
   );
   gpc1_1 gpc701 (
      {stage0_53[51]},
      {stage1_53[38]}
   );
   gpc1_1 gpc702 (
      {stage0_53[52]},
      {stage1_53[39]}
   );
   gpc1_1 gpc703 (
      {stage0_53[53]},
      {stage1_53[40]}
   );
   gpc1_1 gpc704 (
      {stage0_54[51]},
      {stage1_54[14]}
   );
   gpc1_1 gpc705 (
      {stage0_54[52]},
      {stage1_54[15]}
   );
   gpc1_1 gpc706 (
      {stage0_54[53]},
      {stage1_54[16]}
   );
   gpc1_1 gpc707 (
      {stage0_55[30]},
      {stage1_55[14]}
   );
   gpc1_1 gpc708 (
      {stage0_55[31]},
      {stage1_55[15]}
   );
   gpc1_1 gpc709 (
      {stage0_55[32]},
      {stage1_55[16]}
   );
   gpc1_1 gpc710 (
      {stage0_55[33]},
      {stage1_55[17]}
   );
   gpc1_1 gpc711 (
      {stage0_55[34]},
      {stage1_55[18]}
   );
   gpc1_1 gpc712 (
      {stage0_55[35]},
      {stage1_55[19]}
   );
   gpc1_1 gpc713 (
      {stage0_55[36]},
      {stage1_55[20]}
   );
   gpc1_1 gpc714 (
      {stage0_55[37]},
      {stage1_55[21]}
   );
   gpc1_1 gpc715 (
      {stage0_55[38]},
      {stage1_55[22]}
   );
   gpc1_1 gpc716 (
      {stage0_55[39]},
      {stage1_55[23]}
   );
   gpc1_1 gpc717 (
      {stage0_55[40]},
      {stage1_55[24]}
   );
   gpc1_1 gpc718 (
      {stage0_55[41]},
      {stage1_55[25]}
   );
   gpc1_1 gpc719 (
      {stage0_55[42]},
      {stage1_55[26]}
   );
   gpc1_1 gpc720 (
      {stage0_55[43]},
      {stage1_55[27]}
   );
   gpc1_1 gpc721 (
      {stage0_55[44]},
      {stage1_55[28]}
   );
   gpc1_1 gpc722 (
      {stage0_55[45]},
      {stage1_55[29]}
   );
   gpc1_1 gpc723 (
      {stage0_55[46]},
      {stage1_55[30]}
   );
   gpc1_1 gpc724 (
      {stage0_55[47]},
      {stage1_55[31]}
   );
   gpc1_1 gpc725 (
      {stage0_55[48]},
      {stage1_55[32]}
   );
   gpc1_1 gpc726 (
      {stage0_55[49]},
      {stage1_55[33]}
   );
   gpc1_1 gpc727 (
      {stage0_55[50]},
      {stage1_55[34]}
   );
   gpc1_1 gpc728 (
      {stage0_55[51]},
      {stage1_55[35]}
   );
   gpc1_1 gpc729 (
      {stage0_55[52]},
      {stage1_55[36]}
   );
   gpc1_1 gpc730 (
      {stage0_55[53]},
      {stage1_55[37]}
   );
   gpc1_1 gpc731 (
      {stage0_57[30]},
      {stage1_57[17]}
   );
   gpc1_1 gpc732 (
      {stage0_57[31]},
      {stage1_57[18]}
   );
   gpc1_1 gpc733 (
      {stage0_57[32]},
      {stage1_57[19]}
   );
   gpc1_1 gpc734 (
      {stage0_57[33]},
      {stage1_57[20]}
   );
   gpc1_1 gpc735 (
      {stage0_57[34]},
      {stage1_57[21]}
   );
   gpc1_1 gpc736 (
      {stage0_57[35]},
      {stage1_57[22]}
   );
   gpc1_1 gpc737 (
      {stage0_57[36]},
      {stage1_57[23]}
   );
   gpc1_1 gpc738 (
      {stage0_57[37]},
      {stage1_57[24]}
   );
   gpc1_1 gpc739 (
      {stage0_57[38]},
      {stage1_57[25]}
   );
   gpc1_1 gpc740 (
      {stage0_57[39]},
      {stage1_57[26]}
   );
   gpc1_1 gpc741 (
      {stage0_57[40]},
      {stage1_57[27]}
   );
   gpc1_1 gpc742 (
      {stage0_57[41]},
      {stage1_57[28]}
   );
   gpc1_1 gpc743 (
      {stage0_57[42]},
      {stage1_57[29]}
   );
   gpc1_1 gpc744 (
      {stage0_57[43]},
      {stage1_57[30]}
   );
   gpc1_1 gpc745 (
      {stage0_57[44]},
      {stage1_57[31]}
   );
   gpc1_1 gpc746 (
      {stage0_57[45]},
      {stage1_57[32]}
   );
   gpc1_1 gpc747 (
      {stage0_57[46]},
      {stage1_57[33]}
   );
   gpc1_1 gpc748 (
      {stage0_57[47]},
      {stage1_57[34]}
   );
   gpc1_1 gpc749 (
      {stage0_57[48]},
      {stage1_57[35]}
   );
   gpc1_1 gpc750 (
      {stage0_57[49]},
      {stage1_57[36]}
   );
   gpc1_1 gpc751 (
      {stage0_57[50]},
      {stage1_57[37]}
   );
   gpc1_1 gpc752 (
      {stage0_57[51]},
      {stage1_57[38]}
   );
   gpc1_1 gpc753 (
      {stage0_57[52]},
      {stage1_57[39]}
   );
   gpc1_1 gpc754 (
      {stage0_57[53]},
      {stage1_57[40]}
   );
   gpc1_1 gpc755 (
      {stage0_59[36]},
      {stage1_59[17]}
   );
   gpc1_1 gpc756 (
      {stage0_59[37]},
      {stage1_59[18]}
   );
   gpc1_1 gpc757 (
      {stage0_59[38]},
      {stage1_59[19]}
   );
   gpc1_1 gpc758 (
      {stage0_59[39]},
      {stage1_59[20]}
   );
   gpc1_1 gpc759 (
      {stage0_59[40]},
      {stage1_59[21]}
   );
   gpc1_1 gpc760 (
      {stage0_59[41]},
      {stage1_59[22]}
   );
   gpc1_1 gpc761 (
      {stage0_59[42]},
      {stage1_59[23]}
   );
   gpc1_1 gpc762 (
      {stage0_59[43]},
      {stage1_59[24]}
   );
   gpc1_1 gpc763 (
      {stage0_59[44]},
      {stage1_59[25]}
   );
   gpc1_1 gpc764 (
      {stage0_59[45]},
      {stage1_59[26]}
   );
   gpc1_1 gpc765 (
      {stage0_59[46]},
      {stage1_59[27]}
   );
   gpc1_1 gpc766 (
      {stage0_59[47]},
      {stage1_59[28]}
   );
   gpc1_1 gpc767 (
      {stage0_59[48]},
      {stage1_59[29]}
   );
   gpc1_1 gpc768 (
      {stage0_59[49]},
      {stage1_59[30]}
   );
   gpc1_1 gpc769 (
      {stage0_59[50]},
      {stage1_59[31]}
   );
   gpc1_1 gpc770 (
      {stage0_59[51]},
      {stage1_59[32]}
   );
   gpc1_1 gpc771 (
      {stage0_59[52]},
      {stage1_59[33]}
   );
   gpc1_1 gpc772 (
      {stage0_59[53]},
      {stage1_59[34]}
   );
   gpc1_1 gpc773 (
      {stage0_62[48]},
      {stage1_62[18]}
   );
   gpc1_1 gpc774 (
      {stage0_62[49]},
      {stage1_62[19]}
   );
   gpc1_1 gpc775 (
      {stage0_62[50]},
      {stage1_62[20]}
   );
   gpc1_1 gpc776 (
      {stage0_62[51]},
      {stage1_62[21]}
   );
   gpc1_1 gpc777 (
      {stage0_62[52]},
      {stage1_62[22]}
   );
   gpc1_1 gpc778 (
      {stage0_62[53]},
      {stage1_62[23]}
   );
   gpc1_1 gpc779 (
      {stage0_63[36]},
      {stage1_63[17]}
   );
   gpc1_1 gpc780 (
      {stage0_63[37]},
      {stage1_63[18]}
   );
   gpc1_1 gpc781 (
      {stage0_63[38]},
      {stage1_63[19]}
   );
   gpc1_1 gpc782 (
      {stage0_63[39]},
      {stage1_63[20]}
   );
   gpc1_1 gpc783 (
      {stage0_63[40]},
      {stage1_63[21]}
   );
   gpc1_1 gpc784 (
      {stage0_63[41]},
      {stage1_63[22]}
   );
   gpc1_1 gpc785 (
      {stage0_63[42]},
      {stage1_63[23]}
   );
   gpc1_1 gpc786 (
      {stage0_63[43]},
      {stage1_63[24]}
   );
   gpc1_1 gpc787 (
      {stage0_63[44]},
      {stage1_63[25]}
   );
   gpc1_1 gpc788 (
      {stage0_63[45]},
      {stage1_63[26]}
   );
   gpc1_1 gpc789 (
      {stage0_63[46]},
      {stage1_63[27]}
   );
   gpc1_1 gpc790 (
      {stage0_63[47]},
      {stage1_63[28]}
   );
   gpc1_1 gpc791 (
      {stage0_63[48]},
      {stage1_63[29]}
   );
   gpc1_1 gpc792 (
      {stage0_63[49]},
      {stage1_63[30]}
   );
   gpc1_1 gpc793 (
      {stage0_63[50]},
      {stage1_63[31]}
   );
   gpc1_1 gpc794 (
      {stage0_63[51]},
      {stage1_63[32]}
   );
   gpc1_1 gpc795 (
      {stage0_63[52]},
      {stage1_63[33]}
   );
   gpc1_1 gpc796 (
      {stage0_63[53]},
      {stage1_63[34]}
   );
   gpc1163_5 gpc797 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc798 (
      {stage1_0[3], stage1_0[4], stage1_0[5], stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc799 (
      {stage1_0[9], stage1_0[10], stage1_0[11], stage1_0[12], stage1_0[13]},
      {stage1_1[6]},
      {stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc2135_5 gpc800 (
      {stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[13], stage1_2[14], stage1_2[15]},
      {stage1_3[1]},
      {stage1_4[0], stage1_4[1]},
      {stage2_5[0],stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3]}
   );
   gpc606_5 gpc801 (
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6], stage1_3[7]},
      {stage2_5[1],stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4]}
   );
   gpc615_5 gpc802 (
      {stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12]},
      {stage1_4[2]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[0],stage2_5[2],stage2_4[5],stage2_3[5]}
   );
   gpc615_5 gpc803 (
      {stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage1_4[3]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[1],stage2_5[3],stage2_4[6],stage2_3[6]}
   );
   gpc615_5 gpc804 (
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22]},
      {stage1_4[4]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[2],stage2_5[4],stage2_4[7],stage2_3[7]}
   );
   gpc2135_5 gpc805 (
      {stage1_4[5], stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9]},
      {stage1_5[18], stage1_5[19], stage1_5[20]},
      {stage1_6[0]},
      {stage1_7[0], stage1_7[1]},
      {stage2_8[0],stage2_7[3],stage2_6[3],stage2_5[5],stage2_4[8]}
   );
   gpc2135_5 gpc806 (
      {stage1_4[10], stage1_4[11], stage1_4[12], stage1_4[13], stage1_4[14]},
      {stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_6[1]},
      {stage1_7[2], stage1_7[3]},
      {stage2_8[1],stage2_7[4],stage2_6[4],stage2_5[6],stage2_4[9]}
   );
   gpc606_5 gpc807 (
      {stage1_4[15], stage1_4[16], stage1_4[17], stage1_4[18], stage1_4[19], stage1_4[20]},
      {stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6], stage1_6[7]},
      {stage2_8[2],stage2_7[5],stage2_6[5],stage2_5[7],stage2_4[10]}
   );
   gpc606_5 gpc808 (
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage1_7[4], stage1_7[5], stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9]},
      {stage2_9[0],stage2_8[3],stage2_7[6],stage2_6[6],stage2_5[8]}
   );
   gpc606_5 gpc809 (
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage1_7[10], stage1_7[11], stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15]},
      {stage2_9[1],stage2_8[4],stage2_7[7],stage2_6[7],stage2_5[9]}
   );
   gpc615_5 gpc810 (
      {stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage1_7[16]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[2],stage2_8[5],stage2_7[8],stage2_6[8]}
   );
   gpc615_5 gpc811 (
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage1_7[17]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[3],stage2_8[6],stage2_7[9],stage2_6[9]}
   );
   gpc615_5 gpc812 (
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22]},
      {stage1_8[12]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[2],stage2_9[4],stage2_8[7],stage2_7[10]}
   );
   gpc606_5 gpc813 (
      {stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17], stage1_8[18]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[1],stage2_10[3],stage2_9[5],stage2_8[8]}
   );
   gpc606_5 gpc814 (
      {stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23], stage1_8[24]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[2],stage2_10[4],stage2_9[6],stage2_8[9]}
   );
   gpc606_5 gpc815 (
      {stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29], stage1_8[30]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[3],stage2_10[5],stage2_9[7],stage2_8[10]}
   );
   gpc615_5 gpc816 (
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22]},
      {stage1_11[0]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[0],stage2_12[3],stage2_11[4],stage2_10[6]}
   );
   gpc1415_5 gpc817 (
      {stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage1_12[6]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[1],stage2_13[1],stage2_12[4],stage2_11[5]}
   );
   gpc1415_5 gpc818 (
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10]},
      {stage1_12[7]},
      {stage1_13[4], stage1_13[5], stage1_13[6], stage1_13[7]},
      {stage1_14[1]},
      {stage2_15[1],stage2_14[2],stage2_13[2],stage2_12[5],stage2_11[6]}
   );
   gpc1163_5 gpc819 (
      {stage1_11[11], stage1_11[12], stage1_11[13]},
      {stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11], stage1_12[12], stage1_12[13]},
      {stage1_13[8]},
      {stage1_14[2]},
      {stage2_15[2],stage2_14[3],stage2_13[3],stage2_12[6],stage2_11[7]}
   );
   gpc1163_5 gpc820 (
      {stage1_11[14], stage1_11[15], stage1_11[16]},
      {stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17], stage1_12[18], stage1_12[19]},
      {stage1_13[9]},
      {stage1_14[3]},
      {stage2_15[3],stage2_14[4],stage2_13[4],stage2_12[7],stage2_11[8]}
   );
   gpc615_5 gpc821 (
      {stage1_11[17], stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21]},
      {stage1_12[20]},
      {stage1_13[10], stage1_13[11], stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15]},
      {stage2_15[4],stage2_14[5],stage2_13[5],stage2_12[8],stage2_11[9]}
   );
   gpc615_5 gpc822 (
      {stage1_11[22], stage1_11[23], stage1_11[24], stage1_11[25], stage1_11[26]},
      {1'b0},
      {stage1_13[16], stage1_13[17], stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21]},
      {stage2_15[5],stage2_14[6],stage2_13[6],stage2_12[9],stage2_11[10]}
   );
   gpc606_5 gpc823 (
      {stage1_13[22], stage1_13[23], stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[0],stage2_15[6],stage2_14[7],stage2_13[7]}
   );
   gpc1343_5 gpc824 (
      {stage1_14[4], stage1_14[5], stage1_14[6]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9]},
      {stage1_16[0], stage1_16[1], stage1_16[2]},
      {stage1_17[0]},
      {stage2_18[0],stage2_17[1],stage2_16[1],stage2_15[7],stage2_14[8]}
   );
   gpc1343_5 gpc825 (
      {stage1_14[7], stage1_14[8], stage1_14[9]},
      {stage1_15[10], stage1_15[11], stage1_15[12], stage1_15[13]},
      {stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage1_17[1]},
      {stage2_18[1],stage2_17[2],stage2_16[2],stage2_15[8],stage2_14[9]}
   );
   gpc1163_5 gpc826 (
      {stage1_14[10], stage1_14[11], stage1_14[12]},
      {stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17], stage1_15[18], stage1_15[19]},
      {stage1_16[6]},
      {stage1_17[2]},
      {stage2_18[2],stage2_17[3],stage2_16[3],stage2_15[9],stage2_14[10]}
   );
   gpc1163_5 gpc827 (
      {stage1_14[13], stage1_14[14], stage1_14[15]},
      {stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23], stage1_15[24], stage1_15[25]},
      {stage1_16[7]},
      {stage1_17[3]},
      {stage2_18[3],stage2_17[4],stage2_16[4],stage2_15[10],stage2_14[11]}
   );
   gpc1163_5 gpc828 (
      {stage1_14[16], stage1_14[17], stage1_14[18]},
      {stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29], stage1_15[30], stage1_15[31]},
      {stage1_16[8]},
      {stage1_17[4]},
      {stage2_18[4],stage2_17[5],stage2_16[5],stage2_15[11],stage2_14[12]}
   );
   gpc1163_5 gpc829 (
      {stage1_14[19], stage1_14[20], stage1_14[21]},
      {stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37]},
      {stage1_16[9]},
      {stage1_17[5]},
      {stage2_18[5],stage2_17[6],stage2_16[6],stage2_15[12],stage2_14[13]}
   );
   gpc1163_5 gpc830 (
      {stage1_14[22], stage1_14[23], 1'b0},
      {stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41], stage1_15[42], 1'b0},
      {stage1_16[10]},
      {stage1_17[6]},
      {stage2_18[6],stage2_17[7],stage2_16[7],stage2_15[13],stage2_14[14]}
   );
   gpc606_5 gpc831 (
      {stage1_16[11], stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[0],stage2_18[7],stage2_17[8],stage2_16[8]}
   );
   gpc606_5 gpc832 (
      {stage1_16[17], stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[1],stage2_18[8],stage2_17[9],stage2_16[9]}
   );
   gpc606_5 gpc833 (
      {stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11], stage1_17[12]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[2],stage2_19[2],stage2_18[9],stage2_17[10]}
   );
   gpc615_5 gpc834 (
      {stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage1_18[12]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[3],stage2_19[3],stage2_18[10],stage2_17[11]}
   );
   gpc615_5 gpc835 (
      {stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage1_19[12]},
      {stage1_20[0], stage1_20[1], stage1_20[2], stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage2_22[0],stage2_21[2],stage2_20[4],stage2_19[4],stage2_18[11]}
   );
   gpc615_5 gpc836 (
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22]},
      {stage1_19[13]},
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage2_22[1],stage2_21[3],stage2_20[5],stage2_19[5],stage2_18[12]}
   );
   gpc615_5 gpc837 (
      {stage1_18[23], stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27]},
      {stage1_19[14]},
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage2_22[2],stage2_21[4],stage2_20[6],stage2_19[6],stage2_18[13]}
   );
   gpc615_5 gpc838 (
      {stage1_19[15], stage1_19[16], stage1_19[17], stage1_19[18], stage1_19[19]},
      {stage1_20[18]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[3],stage2_21[5],stage2_20[7],stage2_19[7]}
   );
   gpc1343_5 gpc839 (
      {stage1_21[6], stage1_21[7], stage1_21[8]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3]},
      {stage1_23[0], stage1_23[1], stage1_23[2]},
      {stage1_24[0]},
      {stage2_25[0],stage2_24[0],stage2_23[1],stage2_22[4],stage2_21[6]}
   );
   gpc1343_5 gpc840 (
      {stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage1_22[4], stage1_22[5], stage1_22[6], stage1_22[7]},
      {stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage1_24[1]},
      {stage2_25[1],stage2_24[1],stage2_23[2],stage2_22[5],stage2_21[7]}
   );
   gpc606_5 gpc841 (
      {stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11], stage1_22[12], stage1_22[13]},
      {stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5], stage1_24[6], stage1_24[7]},
      {stage2_26[0],stage2_25[2],stage2_24[2],stage2_23[3],stage2_22[6]}
   );
   gpc606_5 gpc842 (
      {stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17], stage1_22[18], stage1_22[19]},
      {stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11], stage1_24[12], stage1_24[13]},
      {stage2_26[1],stage2_25[3],stage2_24[3],stage2_23[4],stage2_22[7]}
   );
   gpc615_5 gpc843 (
      {stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17], stage1_24[18]},
      {stage1_25[0]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[0],stage2_26[2],stage2_25[4],stage2_24[4]}
   );
   gpc615_5 gpc844 (
      {stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage1_25[1]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[1],stage2_26[3],stage2_25[5],stage2_24[5]}
   );
   gpc615_5 gpc845 (
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28]},
      {stage1_25[2]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[2],stage2_26[4],stage2_25[6],stage2_24[6]}
   );
   gpc615_5 gpc846 (
      {stage1_25[3], stage1_25[4], stage1_25[5], stage1_25[6], stage1_25[7]},
      {stage1_26[18]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[3],stage2_27[3],stage2_26[5],stage2_25[7]}
   );
   gpc615_5 gpc847 (
      {stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11], stage1_25[12]},
      {stage1_26[19]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[4],stage2_27[4],stage2_26[6],stage2_25[8]}
   );
   gpc615_5 gpc848 (
      {stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage1_26[20]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[5],stage2_27[5],stage2_26[7],stage2_25[9]}
   );
   gpc615_5 gpc849 (
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22]},
      {stage1_26[21]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[6],stage2_27[6],stage2_26[8],stage2_25[10]}
   );
   gpc1343_5 gpc850 (
      {stage1_28[0], stage1_28[1], stage1_28[2]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3]},
      {stage1_30[0], stage1_30[1], stage1_30[2]},
      {stage1_31[0]},
      {stage2_32[0],stage2_31[0],stage2_30[0],stage2_29[4],stage2_28[7]}
   );
   gpc1343_5 gpc851 (
      {stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage1_29[4], stage1_29[5], stage1_29[6], stage1_29[7]},
      {stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage1_31[1]},
      {stage2_32[1],stage2_31[1],stage2_30[1],stage2_29[5],stage2_28[8]}
   );
   gpc1343_5 gpc852 (
      {stage1_28[6], stage1_28[7], stage1_28[8]},
      {stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage1_30[6], stage1_30[7], stage1_30[8]},
      {stage1_31[2]},
      {stage2_32[2],stage2_31[2],stage2_30[2],stage2_29[6],stage2_28[9]}
   );
   gpc606_5 gpc853 (
      {stage1_28[9], stage1_28[10], stage1_28[11], stage1_28[12], stage1_28[13], stage1_28[14]},
      {stage1_30[9], stage1_30[10], stage1_30[11], stage1_30[12], stage1_30[13], stage1_30[14]},
      {stage2_32[3],stage2_31[3],stage2_30[3],stage2_29[7],stage2_28[10]}
   );
   gpc615_5 gpc854 (
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16]},
      {stage1_30[15]},
      {stage1_31[3], stage1_31[4], stage1_31[5], stage1_31[6], stage1_31[7], stage1_31[8]},
      {stage2_33[0],stage2_32[4],stage2_31[4],stage2_30[4],stage2_29[8]}
   );
   gpc606_5 gpc855 (
      {stage1_30[16], stage1_30[17], stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[1],stage2_32[5],stage2_31[5],stage2_30[5]}
   );
   gpc606_5 gpc856 (
      {stage1_30[22], stage1_30[23], stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27]},
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage2_34[1],stage2_33[2],stage2_32[6],stage2_31[6],stage2_30[6]}
   );
   gpc615_5 gpc857 (
      {stage1_30[28], stage1_30[29], stage1_30[30], stage1_30[31], stage1_30[32]},
      {stage1_31[9]},
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage2_34[2],stage2_33[3],stage2_32[7],stage2_31[7],stage2_30[7]}
   );
   gpc606_5 gpc858 (
      {stage1_31[10], stage1_31[11], stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[3],stage2_33[4],stage2_32[8],stage2_31[8]}
   );
   gpc606_5 gpc859 (
      {stage1_31[16], stage1_31[17], stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[4],stage2_33[5],stage2_32[9],stage2_31[9]}
   );
   gpc606_5 gpc860 (
      {stage1_31[22], stage1_31[23], stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27]},
      {stage1_33[12], stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17]},
      {stage2_35[2],stage2_34[5],stage2_33[6],stage2_32[10],stage2_31[10]}
   );
   gpc606_5 gpc861 (
      {stage1_33[18], stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23]},
      {stage1_35[0], stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5]},
      {stage2_37[0],stage2_36[0],stage2_35[3],stage2_34[6],stage2_33[7]}
   );
   gpc606_5 gpc862 (
      {stage1_33[24], stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29]},
      {stage1_35[6], stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11]},
      {stage2_37[1],stage2_36[1],stage2_35[4],stage2_34[7],stage2_33[8]}
   );
   gpc606_5 gpc863 (
      {stage1_33[30], stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35]},
      {stage1_35[12], stage1_35[13], stage1_35[14], stage1_35[15], stage1_35[16], stage1_35[17]},
      {stage2_37[2],stage2_36[2],stage2_35[5],stage2_34[8],stage2_33[9]}
   );
   gpc615_5 gpc864 (
      {stage1_33[36], stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40]},
      {stage1_34[0]},
      {stage1_35[18], stage1_35[19], stage1_35[20], stage1_35[21], stage1_35[22], stage1_35[23]},
      {stage2_37[3],stage2_36[3],stage2_35[6],stage2_34[9],stage2_33[10]}
   );
   gpc615_5 gpc865 (
      {stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage1_35[24]},
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5]},
      {stage2_38[0],stage2_37[4],stage2_36[4],stage2_35[7],stage2_34[10]}
   );
   gpc615_5 gpc866 (
      {stage1_34[6], stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10]},
      {stage1_35[25]},
      {stage1_36[6], stage1_36[7], stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11]},
      {stage2_38[1],stage2_37[5],stage2_36[5],stage2_35[8],stage2_34[11]}
   );
   gpc615_5 gpc867 (
      {stage1_34[11], stage1_34[12], stage1_34[13], stage1_34[14], stage1_34[15]},
      {stage1_35[26]},
      {stage1_36[12], stage1_36[13], stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17]},
      {stage2_38[2],stage2_37[6],stage2_36[6],stage2_35[9],stage2_34[12]}
   );
   gpc615_5 gpc868 (
      {stage1_36[18], stage1_36[19], stage1_36[20], stage1_36[21], stage1_36[22]},
      {stage1_37[0]},
      {stage1_38[0], stage1_38[1], stage1_38[2], stage1_38[3], stage1_38[4], stage1_38[5]},
      {stage2_40[0],stage2_39[0],stage2_38[3],stage2_37[7],stage2_36[7]}
   );
   gpc606_5 gpc869 (
      {stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5], stage1_37[6]},
      {stage1_39[0], stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5]},
      {stage2_41[0],stage2_40[1],stage2_39[1],stage2_38[4],stage2_37[8]}
   );
   gpc606_5 gpc870 (
      {stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11], stage1_37[12]},
      {stage1_39[6], stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11]},
      {stage2_41[1],stage2_40[2],stage2_39[2],stage2_38[5],stage2_37[9]}
   );
   gpc606_5 gpc871 (
      {stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17], stage1_37[18]},
      {stage1_39[12], stage1_39[13], stage1_39[14], stage1_39[15], stage1_39[16], stage1_39[17]},
      {stage2_41[2],stage2_40[3],stage2_39[3],stage2_38[6],stage2_37[10]}
   );
   gpc615_5 gpc872 (
      {stage1_38[6], stage1_38[7], stage1_38[8], stage1_38[9], stage1_38[10]},
      {stage1_39[18]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3], stage1_40[4], stage1_40[5]},
      {stage2_42[0],stage2_41[3],stage2_40[4],stage2_39[4],stage2_38[7]}
   );
   gpc615_5 gpc873 (
      {stage1_38[11], stage1_38[12], stage1_38[13], stage1_38[14], stage1_38[15]},
      {stage1_39[19]},
      {stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10], stage1_40[11]},
      {stage2_42[1],stage2_41[4],stage2_40[5],stage2_39[5],stage2_38[8]}
   );
   gpc615_5 gpc874 (
      {stage1_38[16], stage1_38[17], stage1_38[18], stage1_38[19], stage1_38[20]},
      {stage1_39[20]},
      {stage1_40[12], stage1_40[13], stage1_40[14], stage1_40[15], stage1_40[16], stage1_40[17]},
      {stage2_42[2],stage2_41[5],stage2_40[6],stage2_39[6],stage2_38[9]}
   );
   gpc1163_5 gpc875 (
      {stage1_40[18], stage1_40[19], stage1_40[20]},
      {stage1_41[0], stage1_41[1], stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5]},
      {stage1_42[0]},
      {stage1_43[0]},
      {stage2_44[0],stage2_43[0],stage2_42[3],stage2_41[6],stage2_40[7]}
   );
   gpc1163_5 gpc876 (
      {stage1_40[21], stage1_40[22], stage1_40[23]},
      {stage1_41[6], stage1_41[7], stage1_41[8], stage1_41[9], stage1_41[10], stage1_41[11]},
      {stage1_42[1]},
      {stage1_43[1]},
      {stage2_44[1],stage2_43[1],stage2_42[4],stage2_41[7],stage2_40[8]}
   );
   gpc1163_5 gpc877 (
      {stage1_40[24], stage1_40[25], stage1_40[26]},
      {stage1_41[12], stage1_41[13], stage1_41[14], stage1_41[15], stage1_41[16], stage1_41[17]},
      {stage1_42[2]},
      {stage1_43[2]},
      {stage2_44[2],stage2_43[2],stage2_42[5],stage2_41[8],stage2_40[9]}
   );
   gpc606_5 gpc878 (
      {stage1_40[27], stage1_40[28], stage1_40[29], stage1_40[30], stage1_40[31], stage1_40[32]},
      {stage1_42[3], stage1_42[4], stage1_42[5], stage1_42[6], stage1_42[7], stage1_42[8]},
      {stage2_44[3],stage2_43[3],stage2_42[6],stage2_41[9],stage2_40[10]}
   );
   gpc606_5 gpc879 (
      {stage1_40[33], stage1_40[34], stage1_40[35], stage1_40[36], stage1_40[37], stage1_40[38]},
      {stage1_42[9], stage1_42[10], stage1_42[11], stage1_42[12], stage1_42[13], stage1_42[14]},
      {stage2_44[4],stage2_43[4],stage2_42[7],stage2_41[10],stage2_40[11]}
   );
   gpc606_5 gpc880 (
      {stage1_43[3], stage1_43[4], stage1_43[5], stage1_43[6], stage1_43[7], stage1_43[8]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5]},
      {stage2_47[0],stage2_46[0],stage2_45[0],stage2_44[5],stage2_43[5]}
   );
   gpc606_5 gpc881 (
      {stage1_43[9], stage1_43[10], stage1_43[11], stage1_43[12], stage1_43[13], stage1_43[14]},
      {stage1_45[6], stage1_45[7], stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage2_47[1],stage2_46[1],stage2_45[1],stage2_44[6],stage2_43[6]}
   );
   gpc606_5 gpc882 (
      {stage1_43[15], stage1_43[16], stage1_43[17], stage1_43[18], stage1_43[19], stage1_43[20]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15], stage1_45[16], stage1_45[17]},
      {stage2_47[2],stage2_46[2],stage2_45[2],stage2_44[7],stage2_43[7]}
   );
   gpc606_5 gpc883 (
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4], stage1_44[5]},
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4], stage1_46[5]},
      {stage2_48[0],stage2_47[3],stage2_46[3],stage2_45[3],stage2_44[8]}
   );
   gpc606_5 gpc884 (
      {stage1_44[6], stage1_44[7], stage1_44[8], stage1_44[9], stage1_44[10], stage1_44[11]},
      {stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9], stage1_46[10], stage1_46[11]},
      {stage2_48[1],stage2_47[4],stage2_46[4],stage2_45[4],stage2_44[9]}
   );
   gpc606_5 gpc885 (
      {stage1_44[12], stage1_44[13], stage1_44[14], stage1_44[15], stage1_44[16], stage1_44[17]},
      {stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15], stage1_46[16], stage1_46[17]},
      {stage2_48[2],stage2_47[5],stage2_46[5],stage2_45[5],stage2_44[10]}
   );
   gpc615_5 gpc886 (
      {stage1_45[18], stage1_45[19], stage1_45[20], stage1_45[21], stage1_45[22]},
      {stage1_46[18]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[3],stage2_47[6],stage2_46[6],stage2_45[6]}
   );
   gpc615_5 gpc887 (
      {stage1_45[23], stage1_45[24], stage1_45[25], stage1_45[26], stage1_45[27]},
      {stage1_46[19]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[4],stage2_47[7],stage2_46[7],stage2_45[7]}
   );
   gpc615_5 gpc888 (
      {stage1_47[12], stage1_47[13], stage1_47[14], stage1_47[15], stage1_47[16]},
      {stage1_48[0]},
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage2_51[0],stage2_50[0],stage2_49[2],stage2_48[5],stage2_47[8]}
   );
   gpc615_5 gpc889 (
      {stage1_47[17], stage1_47[18], stage1_47[19], stage1_47[20], stage1_47[21]},
      {stage1_48[1]},
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10], stage1_49[11]},
      {stage2_51[1],stage2_50[1],stage2_49[3],stage2_48[6],stage2_47[9]}
   );
   gpc606_5 gpc890 (
      {stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5], stage1_48[6], stage1_48[7]},
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4], stage1_50[5]},
      {stage2_52[0],stage2_51[2],stage2_50[2],stage2_49[4],stage2_48[7]}
   );
   gpc606_5 gpc891 (
      {stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11], stage1_48[12], stage1_48[13]},
      {stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9], stage1_50[10], stage1_50[11]},
      {stage2_52[1],stage2_51[3],stage2_50[3],stage2_49[5],stage2_48[8]}
   );
   gpc2135_5 gpc892 (
      {stage1_50[12], stage1_50[13], stage1_50[14], stage1_50[15], stage1_50[16]},
      {stage1_51[0], stage1_51[1], stage1_51[2]},
      {stage1_52[0]},
      {stage1_53[0], stage1_53[1]},
      {stage2_54[0],stage2_53[0],stage2_52[2],stage2_51[4],stage2_50[4]}
   );
   gpc2135_5 gpc893 (
      {stage1_50[17], stage1_50[18], stage1_50[19], stage1_50[20], stage1_50[21]},
      {stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage1_52[1]},
      {stage1_53[2], stage1_53[3]},
      {stage2_54[1],stage2_53[1],stage2_52[3],stage2_51[5],stage2_50[5]}
   );
   gpc2135_5 gpc894 (
      {stage1_50[22], stage1_50[23], stage1_50[24], stage1_50[25], stage1_50[26]},
      {stage1_51[6], stage1_51[7], stage1_51[8]},
      {stage1_52[2]},
      {stage1_53[4], stage1_53[5]},
      {stage2_54[2],stage2_53[2],stage2_52[4],stage2_51[6],stage2_50[6]}
   );
   gpc2135_5 gpc895 (
      {stage1_50[27], stage1_50[28], stage1_50[29], stage1_50[30], stage1_50[31]},
      {stage1_51[9], stage1_51[10], stage1_51[11]},
      {stage1_52[3]},
      {stage1_53[6], stage1_53[7]},
      {stage2_54[3],stage2_53[3],stage2_52[5],stage2_51[7],stage2_50[7]}
   );
   gpc2135_5 gpc896 (
      {stage1_50[32], stage1_50[33], stage1_50[34], stage1_50[35], stage1_50[36]},
      {stage1_51[12], stage1_51[13], stage1_51[14]},
      {stage1_52[4]},
      {stage1_53[8], stage1_53[9]},
      {stage2_54[4],stage2_53[4],stage2_52[6],stage2_51[8],stage2_50[8]}
   );
   gpc615_5 gpc897 (
      {stage1_50[37], stage1_50[38], stage1_50[39], stage1_50[40], stage1_50[41]},
      {stage1_51[15]},
      {stage1_52[5], stage1_52[6], stage1_52[7], stage1_52[8], stage1_52[9], stage1_52[10]},
      {stage2_54[5],stage2_53[5],stage2_52[7],stage2_51[9],stage2_50[9]}
   );
   gpc606_5 gpc898 (
      {stage1_51[16], stage1_51[17], stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21]},
      {stage1_53[10], stage1_53[11], stage1_53[12], stage1_53[13], stage1_53[14], stage1_53[15]},
      {stage2_55[0],stage2_54[6],stage2_53[6],stage2_52[8],stage2_51[10]}
   );
   gpc606_5 gpc899 (
      {stage1_51[22], stage1_51[23], stage1_51[24], stage1_51[25], stage1_51[26], stage1_51[27]},
      {stage1_53[16], stage1_53[17], stage1_53[18], stage1_53[19], stage1_53[20], stage1_53[21]},
      {stage2_55[1],stage2_54[7],stage2_53[7],stage2_52[9],stage2_51[11]}
   );
   gpc606_5 gpc900 (
      {stage1_51[28], stage1_51[29], stage1_51[30], stage1_51[31], stage1_51[32], stage1_51[33]},
      {stage1_53[22], stage1_53[23], stage1_53[24], stage1_53[25], stage1_53[26], stage1_53[27]},
      {stage2_55[2],stage2_54[8],stage2_53[8],stage2_52[10],stage2_51[12]}
   );
   gpc606_5 gpc901 (
      {stage1_51[34], stage1_51[35], stage1_51[36], stage1_51[37], stage1_51[38], stage1_51[39]},
      {stage1_53[28], stage1_53[29], stage1_53[30], stage1_53[31], stage1_53[32], stage1_53[33]},
      {stage2_55[3],stage2_54[9],stage2_53[9],stage2_52[11],stage2_51[13]}
   );
   gpc606_5 gpc902 (
      {stage1_51[40], stage1_51[41], stage1_51[42], stage1_51[43], stage1_51[44], stage1_51[45]},
      {stage1_53[34], stage1_53[35], stage1_53[36], stage1_53[37], stage1_53[38], stage1_53[39]},
      {stage2_55[4],stage2_54[10],stage2_53[10],stage2_52[12],stage2_51[14]}
   );
   gpc606_5 gpc903 (
      {stage1_52[11], stage1_52[12], stage1_52[13], stage1_52[14], stage1_52[15], stage1_52[16]},
      {stage1_54[0], stage1_54[1], stage1_54[2], stage1_54[3], stage1_54[4], stage1_54[5]},
      {stage2_56[0],stage2_55[5],stage2_54[11],stage2_53[11],stage2_52[13]}
   );
   gpc615_5 gpc904 (
      {stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9], stage1_54[10]},
      {stage1_55[0]},
      {stage1_56[0], stage1_56[1], stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage2_58[0],stage2_57[0],stage2_56[1],stage2_55[6],stage2_54[12]}
   );
   gpc615_5 gpc905 (
      {stage1_54[11], stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15]},
      {stage1_55[1]},
      {stage1_56[6], stage1_56[7], stage1_56[8], stage1_56[9], stage1_56[10], stage1_56[11]},
      {stage2_58[1],stage2_57[1],stage2_56[2],stage2_55[7],stage2_54[13]}
   );
   gpc606_5 gpc906 (
      {stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5], stage1_55[6], stage1_55[7]},
      {stage1_57[0], stage1_57[1], stage1_57[2], stage1_57[3], stage1_57[4], stage1_57[5]},
      {stage2_59[0],stage2_58[2],stage2_57[2],stage2_56[3],stage2_55[8]}
   );
   gpc606_5 gpc907 (
      {stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11], stage1_55[12], stage1_55[13]},
      {stage1_57[6], stage1_57[7], stage1_57[8], stage1_57[9], stage1_57[10], stage1_57[11]},
      {stage2_59[1],stage2_58[3],stage2_57[3],stage2_56[4],stage2_55[9]}
   );
   gpc606_5 gpc908 (
      {stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17], stage1_55[18], stage1_55[19]},
      {stage1_57[12], stage1_57[13], stage1_57[14], stage1_57[15], stage1_57[16], stage1_57[17]},
      {stage2_59[2],stage2_58[4],stage2_57[4],stage2_56[5],stage2_55[10]}
   );
   gpc606_5 gpc909 (
      {stage1_55[20], stage1_55[21], stage1_55[22], stage1_55[23], stage1_55[24], stage1_55[25]},
      {stage1_57[18], stage1_57[19], stage1_57[20], stage1_57[21], stage1_57[22], stage1_57[23]},
      {stage2_59[3],stage2_58[5],stage2_57[5],stage2_56[6],stage2_55[11]}
   );
   gpc606_5 gpc910 (
      {stage1_55[26], stage1_55[27], stage1_55[28], stage1_55[29], stage1_55[30], stage1_55[31]},
      {stage1_57[24], stage1_57[25], stage1_57[26], stage1_57[27], stage1_57[28], stage1_57[29]},
      {stage2_59[4],stage2_58[6],stage2_57[6],stage2_56[7],stage2_55[12]}
   );
   gpc615_5 gpc911 (
      {stage1_56[12], stage1_56[13], stage1_56[14], stage1_56[15], stage1_56[16]},
      {stage1_57[30]},
      {stage1_58[0], stage1_58[1], stage1_58[2], stage1_58[3], stage1_58[4], stage1_58[5]},
      {stage2_60[0],stage2_59[5],stage2_58[7],stage2_57[7],stage2_56[8]}
   );
   gpc606_5 gpc912 (
      {stage1_57[31], stage1_57[32], stage1_57[33], stage1_57[34], stage1_57[35], stage1_57[36]},
      {stage1_59[0], stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5]},
      {stage2_61[0],stage2_60[1],stage2_59[6],stage2_58[8],stage2_57[8]}
   );
   gpc135_4 gpc913 (
      {stage1_59[6], stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10]},
      {stage1_60[0], stage1_60[1], stage1_60[2]},
      {stage1_61[0]},
      {stage2_62[0],stage2_61[1],stage2_60[2],stage2_59[7]}
   );
   gpc135_4 gpc914 (
      {stage1_59[11], stage1_59[12], stage1_59[13], stage1_59[14], stage1_59[15]},
      {stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage1_61[1]},
      {stage2_62[1],stage2_61[2],stage2_60[3],stage2_59[8]}
   );
   gpc135_4 gpc915 (
      {stage1_59[16], stage1_59[17], stage1_59[18], stage1_59[19], stage1_59[20]},
      {stage1_60[6], stage1_60[7], stage1_60[8]},
      {stage1_61[2]},
      {stage2_62[2],stage2_61[3],stage2_60[4],stage2_59[9]}
   );
   gpc135_4 gpc916 (
      {stage1_59[21], stage1_59[22], stage1_59[23], stage1_59[24], stage1_59[25]},
      {stage1_60[9], stage1_60[10], stage1_60[11]},
      {stage1_61[3]},
      {stage2_62[3],stage2_61[4],stage2_60[5],stage2_59[10]}
   );
   gpc135_4 gpc917 (
      {stage1_59[26], stage1_59[27], stage1_59[28], stage1_59[29], stage1_59[30]},
      {stage1_60[12], stage1_60[13], stage1_60[14]},
      {stage1_61[4]},
      {stage2_62[4],stage2_61[5],stage2_60[6],stage2_59[11]}
   );
   gpc135_4 gpc918 (
      {stage1_59[31], stage1_59[32], stage1_59[33], stage1_59[34], 1'b0},
      {stage1_60[15], stage1_60[16], stage1_60[17]},
      {stage1_61[5]},
      {stage2_62[5],stage2_61[6],stage2_60[7],stage2_59[12]}
   );
   gpc606_5 gpc919 (
      {stage1_61[6], stage1_61[7], stage1_61[8], stage1_61[9], stage1_61[10], stage1_61[11]},
      {stage1_63[0], stage1_63[1], stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5]},
      {stage2_65[0],stage2_64[0],stage2_63[0],stage2_62[6],stage2_61[7]}
   );
   gpc606_5 gpc920 (
      {stage1_61[12], stage1_61[13], stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17]},
      {stage1_63[6], stage1_63[7], stage1_63[8], stage1_63[9], stage1_63[10], stage1_63[11]},
      {stage2_65[1],stage2_64[1],stage2_63[1],stage2_62[7],stage2_61[8]}
   );
   gpc1163_5 gpc921 (
      {stage1_62[0], stage1_62[1], stage1_62[2]},
      {stage1_63[12], stage1_63[13], stage1_63[14], stage1_63[15], stage1_63[16], stage1_63[17]},
      {stage1_64[0]},
      {stage1_65[0]},
      {stage2_66[0],stage2_65[2],stage2_64[2],stage2_63[2],stage2_62[8]}
   );
   gpc1163_5 gpc922 (
      {stage1_62[3], stage1_62[4], stage1_62[5]},
      {stage1_63[18], stage1_63[19], stage1_63[20], stage1_63[21], stage1_63[22], stage1_63[23]},
      {stage1_64[1]},
      {stage1_65[1]},
      {stage2_66[1],stage2_65[3],stage2_64[3],stage2_63[3],stage2_62[9]}
   );
   gpc606_5 gpc923 (
      {stage1_62[6], stage1_62[7], stage1_62[8], stage1_62[9], stage1_62[10], stage1_62[11]},
      {stage1_64[2], stage1_64[3], stage1_64[4], stage1_64[5], stage1_64[6], stage1_64[7]},
      {stage2_66[2],stage2_65[4],stage2_64[4],stage2_63[4],stage2_62[10]}
   );
   gpc606_5 gpc924 (
      {stage1_62[12], stage1_62[13], stage1_62[14], stage1_62[15], stage1_62[16], stage1_62[17]},
      {stage1_64[8], stage1_64[9], stage1_64[10], stage1_64[11], stage1_64[12], stage1_64[13]},
      {stage2_66[3],stage2_65[5],stage2_64[5],stage2_63[5],stage2_62[11]}
   );
   gpc1_1 gpc925 (
      {stage1_0[14]},
      {stage2_0[3]}
   );
   gpc1_1 gpc926 (
      {stage1_0[15]},
      {stage2_0[4]}
   );
   gpc1_1 gpc927 (
      {stage1_0[16]},
      {stage2_0[5]}
   );
   gpc1_1 gpc928 (
      {stage1_1[18]},
      {stage2_1[5]}
   );
   gpc1_1 gpc929 (
      {stage1_1[19]},
      {stage2_1[6]}
   );
   gpc1_1 gpc930 (
      {stage1_2[16]},
      {stage2_2[5]}
   );
   gpc1_1 gpc931 (
      {stage1_2[17]},
      {stage2_2[6]}
   );
   gpc1_1 gpc932 (
      {stage1_2[18]},
      {stage2_2[7]}
   );
   gpc1_1 gpc933 (
      {stage1_2[19]},
      {stage2_2[8]}
   );
   gpc1_1 gpc934 (
      {stage1_2[20]},
      {stage2_2[9]}
   );
   gpc1_1 gpc935 (
      {stage1_2[21]},
      {stage2_2[10]}
   );
   gpc1_1 gpc936 (
      {stage1_2[22]},
      {stage2_2[11]}
   );
   gpc1_1 gpc937 (
      {stage1_2[23]},
      {stage2_2[12]}
   );
   gpc1_1 gpc938 (
      {stage1_2[24]},
      {stage2_2[13]}
   );
   gpc1_1 gpc939 (
      {stage1_3[23]},
      {stage2_3[8]}
   );
   gpc1_1 gpc940 (
      {stage1_4[21]},
      {stage2_4[11]}
   );
   gpc1_1 gpc941 (
      {stage1_4[22]},
      {stage2_4[12]}
   );
   gpc1_1 gpc942 (
      {stage1_4[23]},
      {stage2_4[13]}
   );
   gpc1_1 gpc943 (
      {stage1_4[24]},
      {stage2_4[14]}
   );
   gpc1_1 gpc944 (
      {stage1_4[25]},
      {stage2_4[15]}
   );
   gpc1_1 gpc945 (
      {stage1_4[26]},
      {stage2_4[16]}
   );
   gpc1_1 gpc946 (
      {stage1_4[27]},
      {stage2_4[17]}
   );
   gpc1_1 gpc947 (
      {stage1_4[28]},
      {stage2_4[18]}
   );
   gpc1_1 gpc948 (
      {stage1_4[29]},
      {stage2_4[19]}
   );
   gpc1_1 gpc949 (
      {stage1_4[30]},
      {stage2_4[20]}
   );
   gpc1_1 gpc950 (
      {stage1_4[31]},
      {stage2_4[21]}
   );
   gpc1_1 gpc951 (
      {stage1_4[32]},
      {stage2_4[22]}
   );
   gpc1_1 gpc952 (
      {stage1_6[18]},
      {stage2_6[10]}
   );
   gpc1_1 gpc953 (
      {stage1_7[23]},
      {stage2_7[11]}
   );
   gpc1_1 gpc954 (
      {stage1_7[24]},
      {stage2_7[12]}
   );
   gpc1_1 gpc955 (
      {stage1_9[6]},
      {stage2_9[8]}
   );
   gpc1_1 gpc956 (
      {stage1_9[7]},
      {stage2_9[9]}
   );
   gpc1_1 gpc957 (
      {stage1_9[8]},
      {stage2_9[10]}
   );
   gpc1_1 gpc958 (
      {stage1_9[9]},
      {stage2_9[11]}
   );
   gpc1_1 gpc959 (
      {stage1_9[10]},
      {stage2_9[12]}
   );
   gpc1_1 gpc960 (
      {stage1_9[11]},
      {stage2_9[13]}
   );
   gpc1_1 gpc961 (
      {stage1_9[12]},
      {stage2_9[14]}
   );
   gpc1_1 gpc962 (
      {stage1_9[13]},
      {stage2_9[15]}
   );
   gpc1_1 gpc963 (
      {stage1_9[14]},
      {stage2_9[16]}
   );
   gpc1_1 gpc964 (
      {stage1_9[15]},
      {stage2_9[17]}
   );
   gpc1_1 gpc965 (
      {stage1_9[16]},
      {stage2_9[18]}
   );
   gpc1_1 gpc966 (
      {stage1_9[17]},
      {stage2_9[19]}
   );
   gpc1_1 gpc967 (
      {stage1_10[23]},
      {stage2_10[7]}
   );
   gpc1_1 gpc968 (
      {stage1_10[24]},
      {stage2_10[8]}
   );
   gpc1_1 gpc969 (
      {stage1_10[25]},
      {stage2_10[9]}
   );
   gpc1_1 gpc970 (
      {stage1_11[27]},
      {stage2_11[11]}
   );
   gpc1_1 gpc971 (
      {stage1_11[28]},
      {stage2_11[12]}
   );
   gpc1_1 gpc972 (
      {stage1_13[28]},
      {stage2_13[8]}
   );
   gpc1_1 gpc973 (
      {stage1_13[29]},
      {stage2_13[9]}
   );
   gpc1_1 gpc974 (
      {stage1_16[23]},
      {stage2_16[10]}
   );
   gpc1_1 gpc975 (
      {stage1_18[28]},
      {stage2_18[14]}
   );
   gpc1_1 gpc976 (
      {stage1_18[29]},
      {stage2_18[15]}
   );
   gpc1_1 gpc977 (
      {stage1_18[30]},
      {stage2_18[16]}
   );
   gpc1_1 gpc978 (
      {stage1_18[31]},
      {stage2_18[17]}
   );
   gpc1_1 gpc979 (
      {stage1_18[32]},
      {stage2_18[18]}
   );
   gpc1_1 gpc980 (
      {stage1_18[33]},
      {stage2_18[19]}
   );
   gpc1_1 gpc981 (
      {stage1_19[20]},
      {stage2_19[8]}
   );
   gpc1_1 gpc982 (
      {stage1_20[19]},
      {stage2_20[8]}
   );
   gpc1_1 gpc983 (
      {stage1_21[12]},
      {stage2_21[8]}
   );
   gpc1_1 gpc984 (
      {stage1_21[13]},
      {stage2_21[9]}
   );
   gpc1_1 gpc985 (
      {stage1_21[14]},
      {stage2_21[10]}
   );
   gpc1_1 gpc986 (
      {stage1_21[15]},
      {stage2_21[11]}
   );
   gpc1_1 gpc987 (
      {stage1_21[16]},
      {stage2_21[12]}
   );
   gpc1_1 gpc988 (
      {stage1_21[17]},
      {stage2_21[13]}
   );
   gpc1_1 gpc989 (
      {stage1_21[18]},
      {stage2_21[14]}
   );
   gpc1_1 gpc990 (
      {stage1_21[19]},
      {stage2_21[15]}
   );
   gpc1_1 gpc991 (
      {stage1_21[20]},
      {stage2_21[16]}
   );
   gpc1_1 gpc992 (
      {stage1_21[21]},
      {stage2_21[17]}
   );
   gpc1_1 gpc993 (
      {stage1_21[22]},
      {stage2_21[18]}
   );
   gpc1_1 gpc994 (
      {stage1_21[23]},
      {stage2_21[19]}
   );
   gpc1_1 gpc995 (
      {stage1_21[24]},
      {stage2_21[20]}
   );
   gpc1_1 gpc996 (
      {stage1_21[25]},
      {stage2_21[21]}
   );
   gpc1_1 gpc997 (
      {stage1_22[20]},
      {stage2_22[8]}
   );
   gpc1_1 gpc998 (
      {stage1_22[21]},
      {stage2_22[9]}
   );
   gpc1_1 gpc999 (
      {stage1_22[22]},
      {stage2_22[10]}
   );
   gpc1_1 gpc1000 (
      {stage1_23[6]},
      {stage2_23[5]}
   );
   gpc1_1 gpc1001 (
      {stage1_23[7]},
      {stage2_23[6]}
   );
   gpc1_1 gpc1002 (
      {stage1_23[8]},
      {stage2_23[7]}
   );
   gpc1_1 gpc1003 (
      {stage1_23[9]},
      {stage2_23[8]}
   );
   gpc1_1 gpc1004 (
      {stage1_23[10]},
      {stage2_23[9]}
   );
   gpc1_1 gpc1005 (
      {stage1_23[11]},
      {stage2_23[10]}
   );
   gpc1_1 gpc1006 (
      {stage1_23[12]},
      {stage2_23[11]}
   );
   gpc1_1 gpc1007 (
      {stage1_23[13]},
      {stage2_23[12]}
   );
   gpc1_1 gpc1008 (
      {stage1_23[14]},
      {stage2_23[13]}
   );
   gpc1_1 gpc1009 (
      {stage1_23[15]},
      {stage2_23[14]}
   );
   gpc1_1 gpc1010 (
      {stage1_23[16]},
      {stage2_23[15]}
   );
   gpc1_1 gpc1011 (
      {stage1_23[17]},
      {stage2_23[16]}
   );
   gpc1_1 gpc1012 (
      {stage1_23[18]},
      {stage2_23[17]}
   );
   gpc1_1 gpc1013 (
      {stage1_23[19]},
      {stage2_23[18]}
   );
   gpc1_1 gpc1014 (
      {stage1_23[20]},
      {stage2_23[19]}
   );
   gpc1_1 gpc1015 (
      {stage1_23[21]},
      {stage2_23[20]}
   );
   gpc1_1 gpc1016 (
      {stage1_24[29]},
      {stage2_24[7]}
   );
   gpc1_1 gpc1017 (
      {stage1_24[30]},
      {stage2_24[8]}
   );
   gpc1_1 gpc1018 (
      {stage1_24[31]},
      {stage2_24[9]}
   );
   gpc1_1 gpc1019 (
      {stage1_25[23]},
      {stage2_25[11]}
   );
   gpc1_1 gpc1020 (
      {stage1_25[24]},
      {stage2_25[12]}
   );
   gpc1_1 gpc1021 (
      {stage1_26[22]},
      {stage2_26[9]}
   );
   gpc1_1 gpc1022 (
      {stage1_26[23]},
      {stage2_26[10]}
   );
   gpc1_1 gpc1023 (
      {stage1_26[24]},
      {stage2_26[11]}
   );
   gpc1_1 gpc1024 (
      {stage1_26[25]},
      {stage2_26[12]}
   );
   gpc1_1 gpc1025 (
      {stage1_26[26]},
      {stage2_26[13]}
   );
   gpc1_1 gpc1026 (
      {stage1_26[27]},
      {stage2_26[14]}
   );
   gpc1_1 gpc1027 (
      {stage1_26[28]},
      {stage2_26[15]}
   );
   gpc1_1 gpc1028 (
      {stage1_26[29]},
      {stage2_26[16]}
   );
   gpc1_1 gpc1029 (
      {stage1_26[30]},
      {stage2_26[17]}
   );
   gpc1_1 gpc1030 (
      {stage1_26[31]},
      {stage2_26[18]}
   );
   gpc1_1 gpc1031 (
      {stage1_28[15]},
      {stage2_28[11]}
   );
   gpc1_1 gpc1032 (
      {stage1_28[16]},
      {stage2_28[12]}
   );
   gpc1_1 gpc1033 (
      {stage1_28[17]},
      {stage2_28[13]}
   );
   gpc1_1 gpc1034 (
      {stage1_29[17]},
      {stage2_29[9]}
   );
   gpc1_1 gpc1035 (
      {stage1_29[18]},
      {stage2_29[10]}
   );
   gpc1_1 gpc1036 (
      {stage1_29[19]},
      {stage2_29[11]}
   );
   gpc1_1 gpc1037 (
      {stage1_29[20]},
      {stage2_29[12]}
   );
   gpc1_1 gpc1038 (
      {stage1_29[21]},
      {stage2_29[13]}
   );
   gpc1_1 gpc1039 (
      {stage1_29[22]},
      {stage2_29[14]}
   );
   gpc1_1 gpc1040 (
      {stage1_29[23]},
      {stage2_29[15]}
   );
   gpc1_1 gpc1041 (
      {stage1_29[24]},
      {stage2_29[16]}
   );
   gpc1_1 gpc1042 (
      {stage1_29[25]},
      {stage2_29[17]}
   );
   gpc1_1 gpc1043 (
      {stage1_30[33]},
      {stage2_30[8]}
   );
   gpc1_1 gpc1044 (
      {stage1_30[34]},
      {stage2_30[9]}
   );
   gpc1_1 gpc1045 (
      {stage1_31[28]},
      {stage2_31[11]}
   );
   gpc1_1 gpc1046 (
      {stage1_31[29]},
      {stage2_31[12]}
   );
   gpc1_1 gpc1047 (
      {stage1_31[30]},
      {stage2_31[13]}
   );
   gpc1_1 gpc1048 (
      {stage1_31[31]},
      {stage2_31[14]}
   );
   gpc1_1 gpc1049 (
      {stage1_31[32]},
      {stage2_31[15]}
   );
   gpc1_1 gpc1050 (
      {stage1_31[33]},
      {stage2_31[16]}
   );
   gpc1_1 gpc1051 (
      {stage1_32[18]},
      {stage2_32[11]}
   );
   gpc1_1 gpc1052 (
      {stage1_33[41]},
      {stage2_33[11]}
   );
   gpc1_1 gpc1053 (
      {stage1_33[42]},
      {stage2_33[12]}
   );
   gpc1_1 gpc1054 (
      {stage1_33[43]},
      {stage2_33[13]}
   );
   gpc1_1 gpc1055 (
      {stage1_33[44]},
      {stage2_33[14]}
   );
   gpc1_1 gpc1056 (
      {stage1_33[45]},
      {stage2_33[15]}
   );
   gpc1_1 gpc1057 (
      {stage1_34[16]},
      {stage2_34[13]}
   );
   gpc1_1 gpc1058 (
      {stage1_34[17]},
      {stage2_34[14]}
   );
   gpc1_1 gpc1059 (
      {stage1_34[18]},
      {stage2_34[15]}
   );
   gpc1_1 gpc1060 (
      {stage1_35[27]},
      {stage2_35[10]}
   );
   gpc1_1 gpc1061 (
      {stage1_36[23]},
      {stage2_36[8]}
   );
   gpc1_1 gpc1062 (
      {stage1_36[24]},
      {stage2_36[9]}
   );
   gpc1_1 gpc1063 (
      {stage1_36[25]},
      {stage2_36[10]}
   );
   gpc1_1 gpc1064 (
      {stage1_36[26]},
      {stage2_36[11]}
   );
   gpc1_1 gpc1065 (
      {stage1_36[27]},
      {stage2_36[12]}
   );
   gpc1_1 gpc1066 (
      {stage1_36[28]},
      {stage2_36[13]}
   );
   gpc1_1 gpc1067 (
      {stage1_36[29]},
      {stage2_36[14]}
   );
   gpc1_1 gpc1068 (
      {stage1_36[30]},
      {stage2_36[15]}
   );
   gpc1_1 gpc1069 (
      {stage1_36[31]},
      {stage2_36[16]}
   );
   gpc1_1 gpc1070 (
      {stage1_36[32]},
      {stage2_36[17]}
   );
   gpc1_1 gpc1071 (
      {stage1_36[33]},
      {stage2_36[18]}
   );
   gpc1_1 gpc1072 (
      {stage1_37[19]},
      {stage2_37[11]}
   );
   gpc1_1 gpc1073 (
      {stage1_37[20]},
      {stage2_37[12]}
   );
   gpc1_1 gpc1074 (
      {stage1_37[21]},
      {stage2_37[13]}
   );
   gpc1_1 gpc1075 (
      {stage1_37[22]},
      {stage2_37[14]}
   );
   gpc1_1 gpc1076 (
      {stage1_37[23]},
      {stage2_37[15]}
   );
   gpc1_1 gpc1077 (
      {stage1_37[24]},
      {stage2_37[16]}
   );
   gpc1_1 gpc1078 (
      {stage1_38[21]},
      {stage2_38[10]}
   );
   gpc1_1 gpc1079 (
      {stage1_38[22]},
      {stage2_38[11]}
   );
   gpc1_1 gpc1080 (
      {stage1_38[23]},
      {stage2_38[12]}
   );
   gpc1_1 gpc1081 (
      {stage1_39[21]},
      {stage2_39[7]}
   );
   gpc1_1 gpc1082 (
      {stage1_39[22]},
      {stage2_39[8]}
   );
   gpc1_1 gpc1083 (
      {stage1_39[23]},
      {stage2_39[9]}
   );
   gpc1_1 gpc1084 (
      {stage1_39[24]},
      {stage2_39[10]}
   );
   gpc1_1 gpc1085 (
      {stage1_39[25]},
      {stage2_39[11]}
   );
   gpc1_1 gpc1086 (
      {stage1_39[26]},
      {stage2_39[12]}
   );
   gpc1_1 gpc1087 (
      {stage1_39[27]},
      {stage2_39[13]}
   );
   gpc1_1 gpc1088 (
      {stage1_39[28]},
      {stage2_39[14]}
   );
   gpc1_1 gpc1089 (
      {stage1_39[29]},
      {stage2_39[15]}
   );
   gpc1_1 gpc1090 (
      {stage1_39[30]},
      {stage2_39[16]}
   );
   gpc1_1 gpc1091 (
      {stage1_41[18]},
      {stage2_41[11]}
   );
   gpc1_1 gpc1092 (
      {stage1_41[19]},
      {stage2_41[12]}
   );
   gpc1_1 gpc1093 (
      {stage1_42[15]},
      {stage2_42[8]}
   );
   gpc1_1 gpc1094 (
      {stage1_42[16]},
      {stage2_42[9]}
   );
   gpc1_1 gpc1095 (
      {stage1_42[17]},
      {stage2_42[10]}
   );
   gpc1_1 gpc1096 (
      {stage1_42[18]},
      {stage2_42[11]}
   );
   gpc1_1 gpc1097 (
      {stage1_42[19]},
      {stage2_42[12]}
   );
   gpc1_1 gpc1098 (
      {stage1_42[20]},
      {stage2_42[13]}
   );
   gpc1_1 gpc1099 (
      {stage1_43[21]},
      {stage2_43[8]}
   );
   gpc1_1 gpc1100 (
      {stage1_43[22]},
      {stage2_43[9]}
   );
   gpc1_1 gpc1101 (
      {stage1_44[18]},
      {stage2_44[11]}
   );
   gpc1_1 gpc1102 (
      {stage1_44[19]},
      {stage2_44[12]}
   );
   gpc1_1 gpc1103 (
      {stage1_44[20]},
      {stage2_44[13]}
   );
   gpc1_1 gpc1104 (
      {stage1_44[21]},
      {stage2_44[14]}
   );
   gpc1_1 gpc1105 (
      {stage1_45[28]},
      {stage2_45[8]}
   );
   gpc1_1 gpc1106 (
      {stage1_45[29]},
      {stage2_45[9]}
   );
   gpc1_1 gpc1107 (
      {stage1_45[30]},
      {stage2_45[10]}
   );
   gpc1_1 gpc1108 (
      {stage1_45[31]},
      {stage2_45[11]}
   );
   gpc1_1 gpc1109 (
      {stage1_46[20]},
      {stage2_46[8]}
   );
   gpc1_1 gpc1110 (
      {stage1_46[21]},
      {stage2_46[9]}
   );
   gpc1_1 gpc1111 (
      {stage1_46[22]},
      {stage2_46[10]}
   );
   gpc1_1 gpc1112 (
      {stage1_46[23]},
      {stage2_46[11]}
   );
   gpc1_1 gpc1113 (
      {stage1_46[24]},
      {stage2_46[12]}
   );
   gpc1_1 gpc1114 (
      {stage1_46[25]},
      {stage2_46[13]}
   );
   gpc1_1 gpc1115 (
      {stage1_46[26]},
      {stage2_46[14]}
   );
   gpc1_1 gpc1116 (
      {stage1_46[27]},
      {stage2_46[15]}
   );
   gpc1_1 gpc1117 (
      {stage1_46[28]},
      {stage2_46[16]}
   );
   gpc1_1 gpc1118 (
      {stage1_46[29]},
      {stage2_46[17]}
   );
   gpc1_1 gpc1119 (
      {stage1_47[22]},
      {stage2_47[10]}
   );
   gpc1_1 gpc1120 (
      {stage1_47[23]},
      {stage2_47[11]}
   );
   gpc1_1 gpc1121 (
      {stage1_47[24]},
      {stage2_47[12]}
   );
   gpc1_1 gpc1122 (
      {stage1_47[25]},
      {stage2_47[13]}
   );
   gpc1_1 gpc1123 (
      {stage1_47[26]},
      {stage2_47[14]}
   );
   gpc1_1 gpc1124 (
      {stage1_47[27]},
      {stage2_47[15]}
   );
   gpc1_1 gpc1125 (
      {stage1_47[28]},
      {stage2_47[16]}
   );
   gpc1_1 gpc1126 (
      {stage1_47[29]},
      {stage2_47[17]}
   );
   gpc1_1 gpc1127 (
      {stage1_47[30]},
      {stage2_47[18]}
   );
   gpc1_1 gpc1128 (
      {stage1_47[31]},
      {stage2_47[19]}
   );
   gpc1_1 gpc1129 (
      {stage1_47[32]},
      {stage2_47[20]}
   );
   gpc1_1 gpc1130 (
      {stage1_47[33]},
      {stage2_47[21]}
   );
   gpc1_1 gpc1131 (
      {stage1_48[14]},
      {stage2_48[9]}
   );
   gpc1_1 gpc1132 (
      {stage1_48[15]},
      {stage2_48[10]}
   );
   gpc1_1 gpc1133 (
      {stage1_48[16]},
      {stage2_48[11]}
   );
   gpc1_1 gpc1134 (
      {stage1_48[17]},
      {stage2_48[12]}
   );
   gpc1_1 gpc1135 (
      {stage1_49[12]},
      {stage2_49[6]}
   );
   gpc1_1 gpc1136 (
      {stage1_49[13]},
      {stage2_49[7]}
   );
   gpc1_1 gpc1137 (
      {stage1_49[14]},
      {stage2_49[8]}
   );
   gpc1_1 gpc1138 (
      {stage1_49[15]},
      {stage2_49[9]}
   );
   gpc1_1 gpc1139 (
      {stage1_49[16]},
      {stage2_49[10]}
   );
   gpc1_1 gpc1140 (
      {stage1_49[17]},
      {stage2_49[11]}
   );
   gpc1_1 gpc1141 (
      {stage1_49[18]},
      {stage2_49[12]}
   );
   gpc1_1 gpc1142 (
      {stage1_49[19]},
      {stage2_49[13]}
   );
   gpc1_1 gpc1143 (
      {stage1_49[20]},
      {stage2_49[14]}
   );
   gpc1_1 gpc1144 (
      {stage1_49[21]},
      {stage2_49[15]}
   );
   gpc1_1 gpc1145 (
      {stage1_49[22]},
      {stage2_49[16]}
   );
   gpc1_1 gpc1146 (
      {stage1_49[23]},
      {stage2_49[17]}
   );
   gpc1_1 gpc1147 (
      {stage1_50[42]},
      {stage2_50[10]}
   );
   gpc1_1 gpc1148 (
      {stage1_51[46]},
      {stage2_51[15]}
   );
   gpc1_1 gpc1149 (
      {stage1_51[47]},
      {stage2_51[16]}
   );
   gpc1_1 gpc1150 (
      {stage1_52[17]},
      {stage2_52[14]}
   );
   gpc1_1 gpc1151 (
      {stage1_52[18]},
      {stage2_52[15]}
   );
   gpc1_1 gpc1152 (
      {stage1_52[19]},
      {stage2_52[16]}
   );
   gpc1_1 gpc1153 (
      {stage1_52[20]},
      {stage2_52[17]}
   );
   gpc1_1 gpc1154 (
      {stage1_52[21]},
      {stage2_52[18]}
   );
   gpc1_1 gpc1155 (
      {stage1_53[40]},
      {stage2_53[12]}
   );
   gpc1_1 gpc1156 (
      {stage1_54[16]},
      {stage2_54[14]}
   );
   gpc1_1 gpc1157 (
      {stage1_55[32]},
      {stage2_55[13]}
   );
   gpc1_1 gpc1158 (
      {stage1_55[33]},
      {stage2_55[14]}
   );
   gpc1_1 gpc1159 (
      {stage1_55[34]},
      {stage2_55[15]}
   );
   gpc1_1 gpc1160 (
      {stage1_55[35]},
      {stage2_55[16]}
   );
   gpc1_1 gpc1161 (
      {stage1_55[36]},
      {stage2_55[17]}
   );
   gpc1_1 gpc1162 (
      {stage1_55[37]},
      {stage2_55[18]}
   );
   gpc1_1 gpc1163 (
      {stage1_56[17]},
      {stage2_56[9]}
   );
   gpc1_1 gpc1164 (
      {stage1_56[18]},
      {stage2_56[10]}
   );
   gpc1_1 gpc1165 (
      {stage1_56[19]},
      {stage2_56[11]}
   );
   gpc1_1 gpc1166 (
      {stage1_56[20]},
      {stage2_56[12]}
   );
   gpc1_1 gpc1167 (
      {stage1_57[37]},
      {stage2_57[9]}
   );
   gpc1_1 gpc1168 (
      {stage1_57[38]},
      {stage2_57[10]}
   );
   gpc1_1 gpc1169 (
      {stage1_57[39]},
      {stage2_57[11]}
   );
   gpc1_1 gpc1170 (
      {stage1_57[40]},
      {stage2_57[12]}
   );
   gpc1_1 gpc1171 (
      {stage1_58[6]},
      {stage2_58[9]}
   );
   gpc1_1 gpc1172 (
      {stage1_58[7]},
      {stage2_58[10]}
   );
   gpc1_1 gpc1173 (
      {stage1_58[8]},
      {stage2_58[11]}
   );
   gpc1_1 gpc1174 (
      {stage1_58[9]},
      {stage2_58[12]}
   );
   gpc1_1 gpc1175 (
      {stage1_58[10]},
      {stage2_58[13]}
   );
   gpc1_1 gpc1176 (
      {stage1_58[11]},
      {stage2_58[14]}
   );
   gpc1_1 gpc1177 (
      {stage1_58[12]},
      {stage2_58[15]}
   );
   gpc1_1 gpc1178 (
      {stage1_58[13]},
      {stage2_58[16]}
   );
   gpc1_1 gpc1179 (
      {stage1_58[14]},
      {stage2_58[17]}
   );
   gpc1_1 gpc1180 (
      {stage1_60[18]},
      {stage2_60[8]}
   );
   gpc1_1 gpc1181 (
      {stage1_60[19]},
      {stage2_60[9]}
   );
   gpc1_1 gpc1182 (
      {stage1_60[20]},
      {stage2_60[10]}
   );
   gpc1_1 gpc1183 (
      {stage1_60[21]},
      {stage2_60[11]}
   );
   gpc1_1 gpc1184 (
      {stage1_60[22]},
      {stage2_60[12]}
   );
   gpc1_1 gpc1185 (
      {stage1_61[18]},
      {stage2_61[9]}
   );
   gpc1_1 gpc1186 (
      {stage1_61[19]},
      {stage2_61[10]}
   );
   gpc1_1 gpc1187 (
      {stage1_61[20]},
      {stage2_61[11]}
   );
   gpc1_1 gpc1188 (
      {stage1_62[18]},
      {stage2_62[12]}
   );
   gpc1_1 gpc1189 (
      {stage1_62[19]},
      {stage2_62[13]}
   );
   gpc1_1 gpc1190 (
      {stage1_62[20]},
      {stage2_62[14]}
   );
   gpc1_1 gpc1191 (
      {stage1_62[21]},
      {stage2_62[15]}
   );
   gpc1_1 gpc1192 (
      {stage1_62[22]},
      {stage2_62[16]}
   );
   gpc1_1 gpc1193 (
      {stage1_62[23]},
      {stage2_62[17]}
   );
   gpc1_1 gpc1194 (
      {stage1_63[24]},
      {stage2_63[6]}
   );
   gpc1_1 gpc1195 (
      {stage1_63[25]},
      {stage2_63[7]}
   );
   gpc1_1 gpc1196 (
      {stage1_63[26]},
      {stage2_63[8]}
   );
   gpc1_1 gpc1197 (
      {stage1_63[27]},
      {stage2_63[9]}
   );
   gpc1_1 gpc1198 (
      {stage1_63[28]},
      {stage2_63[10]}
   );
   gpc1_1 gpc1199 (
      {stage1_63[29]},
      {stage2_63[11]}
   );
   gpc1_1 gpc1200 (
      {stage1_63[30]},
      {stage2_63[12]}
   );
   gpc1_1 gpc1201 (
      {stage1_63[31]},
      {stage2_63[13]}
   );
   gpc1_1 gpc1202 (
      {stage1_63[32]},
      {stage2_63[14]}
   );
   gpc1_1 gpc1203 (
      {stage1_63[33]},
      {stage2_63[15]}
   );
   gpc1_1 gpc1204 (
      {stage1_63[34]},
      {stage2_63[16]}
   );
   gpc1_1 gpc1205 (
      {stage1_65[2]},
      {stage2_65[6]}
   );
   gpc1_1 gpc1206 (
      {stage1_65[3]},
      {stage2_65[7]}
   );
   gpc1_1 gpc1207 (
      {stage1_65[4]},
      {stage2_65[8]}
   );
   gpc1_1 gpc1208 (
      {stage1_65[5]},
      {stage2_65[9]}
   );
   gpc615_5 gpc1209 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc1210 (
      {stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5], stage2_1[6]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1]}
   );
   gpc606_5 gpc1211 (
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[1],stage3_4[2],stage3_3[2],stage3_2[2]}
   );
   gpc606_5 gpc1212 (
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[2],stage3_4[3]}
   );
   gpc2135_5 gpc1213 (
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4]},
      {stage2_6[6], stage2_6[7], stage2_6[8]},
      {stage2_7[0]},
      {stage2_8[0], stage2_8[1]},
      {stage3_9[0],stage3_8[1],stage3_7[1],stage3_6[2],stage3_5[3]}
   );
   gpc615_5 gpc1214 (
      {stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5], stage2_8[6]},
      {stage2_9[0]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[0],stage3_10[0],stage3_9[1],stage3_8[2]}
   );
   gpc606_5 gpc1215 (
      {stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5], stage2_9[6]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[1],stage3_11[1],stage3_10[1],stage3_9[2]}
   );
   gpc606_5 gpc1216 (
      {stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11], stage2_9[12]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[2],stage3_11[2],stage3_10[2],stage3_9[3]}
   );
   gpc615_5 gpc1217 (
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4]},
      {stage2_13[0]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[0],stage3_14[0],stage3_13[2],stage3_12[3]}
   );
   gpc615_5 gpc1218 (
      {stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9]},
      {stage2_13[1]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[1],stage3_14[1],stage3_13[3],stage3_12[4]}
   );
   gpc623_5 gpc1219 (
      {stage2_13[2], stage2_13[3], stage2_13[4]},
      {stage2_14[12], stage2_14[13]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[2],stage3_15[2],stage3_14[2],stage3_13[4]}
   );
   gpc623_5 gpc1220 (
      {stage2_13[5], stage2_13[6], stage2_13[7]},
      {stage2_14[14], 1'b0},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[3],stage3_15[3],stage3_14[3],stage3_13[5]}
   );
   gpc135_4 gpc1221 (
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4]},
      {stage2_17[0], stage2_17[1], stage2_17[2]},
      {stage2_18[0]},
      {stage3_19[0],stage3_18[0],stage3_17[2],stage3_16[4]}
   );
   gpc606_5 gpc1222 (
      {stage2_16[5], stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10]},
      {stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5], stage2_18[6]},
      {stage3_20[0],stage3_19[1],stage3_18[1],stage3_17[3],stage3_16[5]}
   );
   gpc606_5 gpc1223 (
      {stage2_17[3], stage2_17[4], stage2_17[5], stage2_17[6], stage2_17[7], stage2_17[8]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[1],stage3_19[2],stage3_18[2],stage3_17[4]}
   );
   gpc1406_5 gpc1224 (
      {stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11], stage2_18[12]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3]},
      {stage2_21[0]},
      {stage3_22[0],stage3_21[1],stage3_20[2],stage3_19[3],stage3_18[3]}
   );
   gpc1406_5 gpc1225 (
      {stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17], stage2_18[18]},
      {stage2_20[4], stage2_20[5], stage2_20[6], stage2_20[7]},
      {stage2_21[1]},
      {stage3_22[1],stage3_21[2],stage3_20[3],stage3_19[4],stage3_18[4]}
   );
   gpc615_5 gpc1226 (
      {stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5], stage2_21[6]},
      {stage2_22[0]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[0],stage3_23[0],stage3_22[2],stage3_21[3]}
   );
   gpc615_5 gpc1227 (
      {stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage2_22[1]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[1],stage3_23[1],stage3_22[3],stage3_21[4]}
   );
   gpc615_5 gpc1228 (
      {stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15], stage2_21[16]},
      {stage2_22[2]},
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16], stage2_23[17]},
      {stage3_25[2],stage3_24[2],stage3_23[2],stage3_22[4],stage3_21[5]}
   );
   gpc1325_5 gpc1229 (
      {stage2_21[17], stage2_21[18], stage2_21[19], stage2_21[20], stage2_21[21]},
      {stage2_22[3], stage2_22[4]},
      {stage2_23[18], stage2_23[19], stage2_23[20]},
      {stage2_24[0]},
      {stage3_25[3],stage3_24[3],stage3_23[3],stage3_22[5],stage3_21[6]}
   );
   gpc606_5 gpc1230 (
      {stage2_22[5], stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10]},
      {stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5], stage2_24[6]},
      {stage3_26[0],stage3_25[4],stage3_24[4],stage3_23[4],stage3_22[6]}
   );
   gpc1343_5 gpc1231 (
      {stage2_24[7], stage2_24[8], stage2_24[9]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3]},
      {stage2_26[0], stage2_26[1], stage2_26[2]},
      {stage2_27[0]},
      {stage3_28[0],stage3_27[0],stage3_26[1],stage3_25[5],stage3_24[5]}
   );
   gpc1325_5 gpc1232 (
      {stage2_25[4], stage2_25[5], stage2_25[6], stage2_25[7], stage2_25[8]},
      {stage2_26[3], stage2_26[4]},
      {stage2_27[1], stage2_27[2], stage2_27[3]},
      {stage2_28[0]},
      {stage3_29[0],stage3_28[1],stage3_27[1],stage3_26[2],stage3_25[6]}
   );
   gpc1325_5 gpc1233 (
      {stage2_25[9], stage2_25[10], stage2_25[11], stage2_25[12], 1'b0},
      {stage2_26[5], stage2_26[6]},
      {stage2_27[4], stage2_27[5], stage2_27[6]},
      {stage2_28[1]},
      {stage3_29[1],stage3_28[2],stage3_27[2],stage3_26[3],stage3_25[7]}
   );
   gpc606_5 gpc1234 (
      {stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11], stage2_26[12]},
      {stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5], stage2_28[6], stage2_28[7]},
      {stage3_30[0],stage3_29[2],stage3_28[3],stage3_27[3],stage3_26[4]}
   );
   gpc606_5 gpc1235 (
      {stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17], stage2_26[18]},
      {stage2_28[8], stage2_28[9], stage2_28[10], stage2_28[11], stage2_28[12], stage2_28[13]},
      {stage3_30[1],stage3_29[3],stage3_28[4],stage3_27[4],stage3_26[5]}
   );
   gpc606_5 gpc1236 (
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[0],stage3_31[0],stage3_30[2],stage3_29[4]}
   );
   gpc606_5 gpc1237 (
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[1],stage3_32[1],stage3_31[1],stage3_30[3],stage3_29[5]}
   );
   gpc615_5 gpc1238 (
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4]},
      {stage2_31[12]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[2],stage3_32[2],stage3_31[2],stage3_30[4]}
   );
   gpc615_5 gpc1239 (
      {stage2_30[5], stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9]},
      {stage2_31[13]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[3],stage3_32[3],stage3_31[3],stage3_30[5]}
   );
   gpc606_5 gpc1240 (
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[0],stage3_35[0],stage3_34[2],stage3_33[4]}
   );
   gpc606_5 gpc1241 (
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage2_36[0], stage2_36[1], stage2_36[2], stage2_36[3], stage2_36[4], stage2_36[5]},
      {stage3_38[0],stage3_37[1],stage3_36[1],stage3_35[1],stage3_34[3]}
   );
   gpc606_5 gpc1242 (
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10], stage2_34[11]},
      {stage2_36[6], stage2_36[7], stage2_36[8], stage2_36[9], stage2_36[10], stage2_36[11]},
      {stage3_38[1],stage3_37[2],stage3_36[2],stage3_35[2],stage3_34[4]}
   );
   gpc615_5 gpc1243 (
      {stage2_35[6], stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10]},
      {stage2_36[12]},
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5]},
      {stage3_39[0],stage3_38[2],stage3_37[3],stage3_36[3],stage3_35[3]}
   );
   gpc615_5 gpc1244 (
      {stage2_36[13], stage2_36[14], stage2_36[15], stage2_36[16], stage2_36[17]},
      {stage2_37[6]},
      {stage2_38[0], stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4], stage2_38[5]},
      {stage3_40[0],stage3_39[1],stage3_38[3],stage3_37[4],stage3_36[4]}
   );
   gpc615_5 gpc1245 (
      {stage2_37[7], stage2_37[8], stage2_37[9], stage2_37[10], stage2_37[11]},
      {stage2_38[6]},
      {stage2_39[0], stage2_39[1], stage2_39[2], stage2_39[3], stage2_39[4], stage2_39[5]},
      {stage3_41[0],stage3_40[1],stage3_39[2],stage3_38[4],stage3_37[5]}
   );
   gpc615_5 gpc1246 (
      {stage2_37[12], stage2_37[13], stage2_37[14], stage2_37[15], stage2_37[16]},
      {stage2_38[7]},
      {stage2_39[6], stage2_39[7], stage2_39[8], stage2_39[9], stage2_39[10], stage2_39[11]},
      {stage3_41[1],stage3_40[2],stage3_39[3],stage3_38[5],stage3_37[6]}
   );
   gpc207_4 gpc1247 (
      {stage2_38[8], stage2_38[9], stage2_38[10], stage2_38[11], stage2_38[12], 1'b0, 1'b0},
      {stage2_40[0], stage2_40[1]},
      {stage3_41[2],stage3_40[3],stage3_39[4],stage3_38[6]}
   );
   gpc615_5 gpc1248 (
      {stage2_39[12], stage2_39[13], stage2_39[14], stage2_39[15], stage2_39[16]},
      {stage2_40[2]},
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4], stage2_41[5]},
      {stage3_43[0],stage3_42[0],stage3_41[3],stage3_40[4],stage3_39[5]}
   );
   gpc606_5 gpc1249 (
      {stage2_40[3], stage2_40[4], stage2_40[5], stage2_40[6], stage2_40[7], stage2_40[8]},
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4], stage2_42[5]},
      {stage3_44[0],stage3_43[1],stage3_42[1],stage3_41[4],stage3_40[5]}
   );
   gpc623_5 gpc1250 (
      {stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage2_41[6], stage2_41[7]},
      {stage2_42[6], stage2_42[7], stage2_42[8], stage2_42[9], stage2_42[10], stage2_42[11]},
      {stage3_44[1],stage3_43[2],stage3_42[2],stage3_41[5],stage3_40[6]}
   );
   gpc606_5 gpc1251 (
      {stage2_41[8], stage2_41[9], stage2_41[10], stage2_41[11], stage2_41[12], 1'b0},
      {stage2_43[0], stage2_43[1], stage2_43[2], stage2_43[3], stage2_43[4], stage2_43[5]},
      {stage3_45[0],stage3_44[2],stage3_43[3],stage3_42[3],stage3_41[6]}
   );
   gpc606_5 gpc1252 (
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[0],stage3_46[0],stage3_45[1],stage3_44[3]}
   );
   gpc606_5 gpc1253 (
      {stage2_44[6], stage2_44[7], stage2_44[8], stage2_44[9], stage2_44[10], stage2_44[11]},
      {stage2_46[6], stage2_46[7], stage2_46[8], stage2_46[9], stage2_46[10], stage2_46[11]},
      {stage3_48[1],stage3_47[1],stage3_46[1],stage3_45[2],stage3_44[4]}
   );
   gpc606_5 gpc1254 (
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage3_49[0],stage3_48[2],stage3_47[2],stage3_46[2],stage3_45[3]}
   );
   gpc606_5 gpc1255 (
      {stage2_45[6], stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11]},
      {stage2_47[6], stage2_47[7], stage2_47[8], stage2_47[9], stage2_47[10], stage2_47[11]},
      {stage3_49[1],stage3_48[3],stage3_47[3],stage3_46[3],stage3_45[4]}
   );
   gpc615_5 gpc1256 (
      {stage2_46[12], stage2_46[13], stage2_46[14], stage2_46[15], stage2_46[16]},
      {stage2_47[12]},
      {stage2_48[0], stage2_48[1], stage2_48[2], stage2_48[3], stage2_48[4], stage2_48[5]},
      {stage3_50[0],stage3_49[2],stage3_48[4],stage3_47[4],stage3_46[4]}
   );
   gpc606_5 gpc1257 (
      {stage2_47[13], stage2_47[14], stage2_47[15], stage2_47[16], stage2_47[17], stage2_47[18]},
      {stage2_49[0], stage2_49[1], stage2_49[2], stage2_49[3], stage2_49[4], stage2_49[5]},
      {stage3_51[0],stage3_50[1],stage3_49[3],stage3_48[5],stage3_47[5]}
   );
   gpc606_5 gpc1258 (
      {stage2_49[6], stage2_49[7], stage2_49[8], stage2_49[9], stage2_49[10], stage2_49[11]},
      {stage2_51[0], stage2_51[1], stage2_51[2], stage2_51[3], stage2_51[4], stage2_51[5]},
      {stage3_53[0],stage3_52[0],stage3_51[1],stage3_50[2],stage3_49[4]}
   );
   gpc606_5 gpc1259 (
      {stage2_49[12], stage2_49[13], stage2_49[14], stage2_49[15], stage2_49[16], stage2_49[17]},
      {stage2_51[6], stage2_51[7], stage2_51[8], stage2_51[9], stage2_51[10], stage2_51[11]},
      {stage3_53[1],stage3_52[1],stage3_51[2],stage3_50[3],stage3_49[5]}
   );
   gpc615_5 gpc1260 (
      {stage2_50[0], stage2_50[1], stage2_50[2], stage2_50[3], stage2_50[4]},
      {stage2_51[12]},
      {stage2_52[0], stage2_52[1], stage2_52[2], stage2_52[3], stage2_52[4], stage2_52[5]},
      {stage3_54[0],stage3_53[2],stage3_52[2],stage3_51[3],stage3_50[4]}
   );
   gpc606_5 gpc1261 (
      {stage2_52[6], stage2_52[7], stage2_52[8], stage2_52[9], stage2_52[10], stage2_52[11]},
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage3_56[0],stage3_55[0],stage3_54[1],stage3_53[3],stage3_52[3]}
   );
   gpc606_5 gpc1262 (
      {stage2_53[0], stage2_53[1], stage2_53[2], stage2_53[3], stage2_53[4], stage2_53[5]},
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5]},
      {stage3_57[0],stage3_56[1],stage3_55[1],stage3_54[2],stage3_53[4]}
   );
   gpc606_5 gpc1263 (
      {stage2_53[6], stage2_53[7], stage2_53[8], stage2_53[9], stage2_53[10], stage2_53[11]},
      {stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9], stage2_55[10], stage2_55[11]},
      {stage3_57[1],stage3_56[2],stage3_55[2],stage3_54[3],stage3_53[5]}
   );
   gpc135_4 gpc1264 (
      {stage2_54[6], stage2_54[7], stage2_54[8], stage2_54[9], stage2_54[10]},
      {stage2_55[12], stage2_55[13], stage2_55[14]},
      {stage2_56[0]},
      {stage3_57[2],stage3_56[3],stage3_55[3],stage3_54[4]}
   );
   gpc135_4 gpc1265 (
      {stage2_54[11], stage2_54[12], stage2_54[13], stage2_54[14], 1'b0},
      {stage2_55[15], stage2_55[16], stage2_55[17]},
      {stage2_56[1]},
      {stage3_57[3],stage3_56[4],stage3_55[4],stage3_54[5]}
   );
   gpc606_5 gpc1266 (
      {stage2_56[2], stage2_56[3], stage2_56[4], stage2_56[5], stage2_56[6], stage2_56[7]},
      {stage2_58[0], stage2_58[1], stage2_58[2], stage2_58[3], stage2_58[4], stage2_58[5]},
      {stage3_60[0],stage3_59[0],stage3_58[0],stage3_57[4],stage3_56[5]}
   );
   gpc135_4 gpc1267 (
      {stage2_57[0], stage2_57[1], stage2_57[2], stage2_57[3], stage2_57[4]},
      {stage2_58[6], stage2_58[7], stage2_58[8]},
      {stage2_59[0]},
      {stage3_60[1],stage3_59[1],stage3_58[1],stage3_57[5]}
   );
   gpc135_4 gpc1268 (
      {stage2_57[5], stage2_57[6], stage2_57[7], stage2_57[8], stage2_57[9]},
      {stage2_58[9], stage2_58[10], stage2_58[11]},
      {stage2_59[1]},
      {stage3_60[2],stage3_59[2],stage3_58[2],stage3_57[6]}
   );
   gpc1163_5 gpc1269 (
      {stage2_57[10], stage2_57[11], stage2_57[12]},
      {stage2_58[12], stage2_58[13], stage2_58[14], stage2_58[15], stage2_58[16], stage2_58[17]},
      {stage2_59[2]},
      {stage2_60[0]},
      {stage3_61[0],stage3_60[3],stage3_59[3],stage3_58[3],stage3_57[7]}
   );
   gpc606_5 gpc1270 (
      {stage2_60[1], stage2_60[2], stage2_60[3], stage2_60[4], stage2_60[5], stage2_60[6]},
      {stage2_62[0], stage2_62[1], stage2_62[2], stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage3_64[0],stage3_63[0],stage3_62[0],stage3_61[1],stage3_60[4]}
   );
   gpc606_5 gpc1271 (
      {stage2_60[7], stage2_60[8], stage2_60[9], stage2_60[10], stage2_60[11], stage2_60[12]},
      {stage2_62[6], stage2_62[7], stage2_62[8], stage2_62[9], stage2_62[10], stage2_62[11]},
      {stage3_64[1],stage3_63[1],stage3_62[1],stage3_61[2],stage3_60[5]}
   );
   gpc606_5 gpc1272 (
      {stage2_61[0], stage2_61[1], stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5]},
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5]},
      {stage3_65[0],stage3_64[2],stage3_63[2],stage3_62[2],stage3_61[3]}
   );
   gpc606_5 gpc1273 (
      {stage2_62[12], stage2_62[13], stage2_62[14], stage2_62[15], stage2_62[16], stage2_62[17]},
      {stage2_64[0], stage2_64[1], stage2_64[2], stage2_64[3], stage2_64[4], stage2_64[5]},
      {stage3_66[0],stage3_65[1],stage3_64[3],stage3_63[3],stage3_62[3]}
   );
   gpc606_5 gpc1274 (
      {stage2_63[6], stage2_63[7], stage2_63[8], stage2_63[9], stage2_63[10], stage2_63[11]},
      {stage2_65[0], stage2_65[1], stage2_65[2], stage2_65[3], stage2_65[4], stage2_65[5]},
      {stage3_67[0],stage3_66[1],stage3_65[2],stage3_64[4],stage3_63[4]}
   );
   gpc1_1 gpc1275 (
      {stage2_0[5]},
      {stage3_0[1]}
   );
   gpc1_1 gpc1276 (
      {stage2_2[12]},
      {stage3_2[3]}
   );
   gpc1_1 gpc1277 (
      {stage2_2[13]},
      {stage3_2[4]}
   );
   gpc1_1 gpc1278 (
      {stage2_3[6]},
      {stage3_3[3]}
   );
   gpc1_1 gpc1279 (
      {stage2_3[7]},
      {stage3_3[4]}
   );
   gpc1_1 gpc1280 (
      {stage2_3[8]},
      {stage3_3[5]}
   );
   gpc1_1 gpc1281 (
      {stage2_4[12]},
      {stage3_4[4]}
   );
   gpc1_1 gpc1282 (
      {stage2_4[13]},
      {stage3_4[5]}
   );
   gpc1_1 gpc1283 (
      {stage2_4[14]},
      {stage3_4[6]}
   );
   gpc1_1 gpc1284 (
      {stage2_4[15]},
      {stage3_4[7]}
   );
   gpc1_1 gpc1285 (
      {stage2_4[16]},
      {stage3_4[8]}
   );
   gpc1_1 gpc1286 (
      {stage2_4[17]},
      {stage3_4[9]}
   );
   gpc1_1 gpc1287 (
      {stage2_4[18]},
      {stage3_4[10]}
   );
   gpc1_1 gpc1288 (
      {stage2_4[19]},
      {stage3_4[11]}
   );
   gpc1_1 gpc1289 (
      {stage2_4[20]},
      {stage3_4[12]}
   );
   gpc1_1 gpc1290 (
      {stage2_4[21]},
      {stage3_4[13]}
   );
   gpc1_1 gpc1291 (
      {stage2_4[22]},
      {stage3_4[14]}
   );
   gpc1_1 gpc1292 (
      {stage2_5[5]},
      {stage3_5[4]}
   );
   gpc1_1 gpc1293 (
      {stage2_5[6]},
      {stage3_5[5]}
   );
   gpc1_1 gpc1294 (
      {stage2_5[7]},
      {stage3_5[6]}
   );
   gpc1_1 gpc1295 (
      {stage2_5[8]},
      {stage3_5[7]}
   );
   gpc1_1 gpc1296 (
      {stage2_5[9]},
      {stage3_5[8]}
   );
   gpc1_1 gpc1297 (
      {stage2_6[9]},
      {stage3_6[3]}
   );
   gpc1_1 gpc1298 (
      {stage2_6[10]},
      {stage3_6[4]}
   );
   gpc1_1 gpc1299 (
      {stage2_7[1]},
      {stage3_7[2]}
   );
   gpc1_1 gpc1300 (
      {stage2_7[2]},
      {stage3_7[3]}
   );
   gpc1_1 gpc1301 (
      {stage2_7[3]},
      {stage3_7[4]}
   );
   gpc1_1 gpc1302 (
      {stage2_7[4]},
      {stage3_7[5]}
   );
   gpc1_1 gpc1303 (
      {stage2_7[5]},
      {stage3_7[6]}
   );
   gpc1_1 gpc1304 (
      {stage2_7[6]},
      {stage3_7[7]}
   );
   gpc1_1 gpc1305 (
      {stage2_7[7]},
      {stage3_7[8]}
   );
   gpc1_1 gpc1306 (
      {stage2_7[8]},
      {stage3_7[9]}
   );
   gpc1_1 gpc1307 (
      {stage2_7[9]},
      {stage3_7[10]}
   );
   gpc1_1 gpc1308 (
      {stage2_7[10]},
      {stage3_7[11]}
   );
   gpc1_1 gpc1309 (
      {stage2_7[11]},
      {stage3_7[12]}
   );
   gpc1_1 gpc1310 (
      {stage2_7[12]},
      {stage3_7[13]}
   );
   gpc1_1 gpc1311 (
      {stage2_8[7]},
      {stage3_8[3]}
   );
   gpc1_1 gpc1312 (
      {stage2_8[8]},
      {stage3_8[4]}
   );
   gpc1_1 gpc1313 (
      {stage2_8[9]},
      {stage3_8[5]}
   );
   gpc1_1 gpc1314 (
      {stage2_8[10]},
      {stage3_8[6]}
   );
   gpc1_1 gpc1315 (
      {stage2_9[13]},
      {stage3_9[4]}
   );
   gpc1_1 gpc1316 (
      {stage2_9[14]},
      {stage3_9[5]}
   );
   gpc1_1 gpc1317 (
      {stage2_9[15]},
      {stage3_9[6]}
   );
   gpc1_1 gpc1318 (
      {stage2_9[16]},
      {stage3_9[7]}
   );
   gpc1_1 gpc1319 (
      {stage2_9[17]},
      {stage3_9[8]}
   );
   gpc1_1 gpc1320 (
      {stage2_9[18]},
      {stage3_9[9]}
   );
   gpc1_1 gpc1321 (
      {stage2_9[19]},
      {stage3_9[10]}
   );
   gpc1_1 gpc1322 (
      {stage2_10[6]},
      {stage3_10[3]}
   );
   gpc1_1 gpc1323 (
      {stage2_10[7]},
      {stage3_10[4]}
   );
   gpc1_1 gpc1324 (
      {stage2_10[8]},
      {stage3_10[5]}
   );
   gpc1_1 gpc1325 (
      {stage2_10[9]},
      {stage3_10[6]}
   );
   gpc1_1 gpc1326 (
      {stage2_11[12]},
      {stage3_11[3]}
   );
   gpc1_1 gpc1327 (
      {stage2_13[8]},
      {stage3_13[6]}
   );
   gpc1_1 gpc1328 (
      {stage2_13[9]},
      {stage3_13[7]}
   );
   gpc1_1 gpc1329 (
      {stage2_15[12]},
      {stage3_15[4]}
   );
   gpc1_1 gpc1330 (
      {stage2_15[13]},
      {stage3_15[5]}
   );
   gpc1_1 gpc1331 (
      {stage2_17[9]},
      {stage3_17[5]}
   );
   gpc1_1 gpc1332 (
      {stage2_17[10]},
      {stage3_17[6]}
   );
   gpc1_1 gpc1333 (
      {stage2_17[11]},
      {stage3_17[7]}
   );
   gpc1_1 gpc1334 (
      {stage2_18[19]},
      {stage3_18[5]}
   );
   gpc1_1 gpc1335 (
      {stage2_19[6]},
      {stage3_19[5]}
   );
   gpc1_1 gpc1336 (
      {stage2_19[7]},
      {stage3_19[6]}
   );
   gpc1_1 gpc1337 (
      {stage2_19[8]},
      {stage3_19[7]}
   );
   gpc1_1 gpc1338 (
      {stage2_20[8]},
      {stage3_20[4]}
   );
   gpc1_1 gpc1339 (
      {stage2_29[12]},
      {stage3_29[6]}
   );
   gpc1_1 gpc1340 (
      {stage2_29[13]},
      {stage3_29[7]}
   );
   gpc1_1 gpc1341 (
      {stage2_29[14]},
      {stage3_29[8]}
   );
   gpc1_1 gpc1342 (
      {stage2_29[15]},
      {stage3_29[9]}
   );
   gpc1_1 gpc1343 (
      {stage2_29[16]},
      {stage3_29[10]}
   );
   gpc1_1 gpc1344 (
      {stage2_29[17]},
      {stage3_29[11]}
   );
   gpc1_1 gpc1345 (
      {stage2_31[14]},
      {stage3_31[4]}
   );
   gpc1_1 gpc1346 (
      {stage2_31[15]},
      {stage3_31[5]}
   );
   gpc1_1 gpc1347 (
      {stage2_31[16]},
      {stage3_31[6]}
   );
   gpc1_1 gpc1348 (
      {stage2_33[6]},
      {stage3_33[5]}
   );
   gpc1_1 gpc1349 (
      {stage2_33[7]},
      {stage3_33[6]}
   );
   gpc1_1 gpc1350 (
      {stage2_33[8]},
      {stage3_33[7]}
   );
   gpc1_1 gpc1351 (
      {stage2_33[9]},
      {stage3_33[8]}
   );
   gpc1_1 gpc1352 (
      {stage2_33[10]},
      {stage3_33[9]}
   );
   gpc1_1 gpc1353 (
      {stage2_33[11]},
      {stage3_33[10]}
   );
   gpc1_1 gpc1354 (
      {stage2_33[12]},
      {stage3_33[11]}
   );
   gpc1_1 gpc1355 (
      {stage2_33[13]},
      {stage3_33[12]}
   );
   gpc1_1 gpc1356 (
      {stage2_33[14]},
      {stage3_33[13]}
   );
   gpc1_1 gpc1357 (
      {stage2_33[15]},
      {stage3_33[14]}
   );
   gpc1_1 gpc1358 (
      {stage2_34[12]},
      {stage3_34[5]}
   );
   gpc1_1 gpc1359 (
      {stage2_34[13]},
      {stage3_34[6]}
   );
   gpc1_1 gpc1360 (
      {stage2_34[14]},
      {stage3_34[7]}
   );
   gpc1_1 gpc1361 (
      {stage2_34[15]},
      {stage3_34[8]}
   );
   gpc1_1 gpc1362 (
      {stage2_36[18]},
      {stage3_36[5]}
   );
   gpc1_1 gpc1363 (
      {stage2_42[12]},
      {stage3_42[4]}
   );
   gpc1_1 gpc1364 (
      {stage2_42[13]},
      {stage3_42[5]}
   );
   gpc1_1 gpc1365 (
      {stage2_43[6]},
      {stage3_43[4]}
   );
   gpc1_1 gpc1366 (
      {stage2_43[7]},
      {stage3_43[5]}
   );
   gpc1_1 gpc1367 (
      {stage2_43[8]},
      {stage3_43[6]}
   );
   gpc1_1 gpc1368 (
      {stage2_43[9]},
      {stage3_43[7]}
   );
   gpc1_1 gpc1369 (
      {stage2_44[12]},
      {stage3_44[5]}
   );
   gpc1_1 gpc1370 (
      {stage2_44[13]},
      {stage3_44[6]}
   );
   gpc1_1 gpc1371 (
      {stage2_44[14]},
      {stage3_44[7]}
   );
   gpc1_1 gpc1372 (
      {stage2_46[17]},
      {stage3_46[5]}
   );
   gpc1_1 gpc1373 (
      {stage2_47[19]},
      {stage3_47[6]}
   );
   gpc1_1 gpc1374 (
      {stage2_47[20]},
      {stage3_47[7]}
   );
   gpc1_1 gpc1375 (
      {stage2_47[21]},
      {stage3_47[8]}
   );
   gpc1_1 gpc1376 (
      {stage2_48[6]},
      {stage3_48[6]}
   );
   gpc1_1 gpc1377 (
      {stage2_48[7]},
      {stage3_48[7]}
   );
   gpc1_1 gpc1378 (
      {stage2_48[8]},
      {stage3_48[8]}
   );
   gpc1_1 gpc1379 (
      {stage2_48[9]},
      {stage3_48[9]}
   );
   gpc1_1 gpc1380 (
      {stage2_48[10]},
      {stage3_48[10]}
   );
   gpc1_1 gpc1381 (
      {stage2_48[11]},
      {stage3_48[11]}
   );
   gpc1_1 gpc1382 (
      {stage2_48[12]},
      {stage3_48[12]}
   );
   gpc1_1 gpc1383 (
      {stage2_50[5]},
      {stage3_50[5]}
   );
   gpc1_1 gpc1384 (
      {stage2_50[6]},
      {stage3_50[6]}
   );
   gpc1_1 gpc1385 (
      {stage2_50[7]},
      {stage3_50[7]}
   );
   gpc1_1 gpc1386 (
      {stage2_50[8]},
      {stage3_50[8]}
   );
   gpc1_1 gpc1387 (
      {stage2_50[9]},
      {stage3_50[9]}
   );
   gpc1_1 gpc1388 (
      {stage2_50[10]},
      {stage3_50[10]}
   );
   gpc1_1 gpc1389 (
      {stage2_51[13]},
      {stage3_51[4]}
   );
   gpc1_1 gpc1390 (
      {stage2_51[14]},
      {stage3_51[5]}
   );
   gpc1_1 gpc1391 (
      {stage2_51[15]},
      {stage3_51[6]}
   );
   gpc1_1 gpc1392 (
      {stage2_51[16]},
      {stage3_51[7]}
   );
   gpc1_1 gpc1393 (
      {stage2_52[12]},
      {stage3_52[4]}
   );
   gpc1_1 gpc1394 (
      {stage2_52[13]},
      {stage3_52[5]}
   );
   gpc1_1 gpc1395 (
      {stage2_52[14]},
      {stage3_52[6]}
   );
   gpc1_1 gpc1396 (
      {stage2_52[15]},
      {stage3_52[7]}
   );
   gpc1_1 gpc1397 (
      {stage2_52[16]},
      {stage3_52[8]}
   );
   gpc1_1 gpc1398 (
      {stage2_52[17]},
      {stage3_52[9]}
   );
   gpc1_1 gpc1399 (
      {stage2_52[18]},
      {stage3_52[10]}
   );
   gpc1_1 gpc1400 (
      {stage2_53[12]},
      {stage3_53[6]}
   );
   gpc1_1 gpc1401 (
      {stage2_55[18]},
      {stage3_55[5]}
   );
   gpc1_1 gpc1402 (
      {stage2_56[8]},
      {stage3_56[6]}
   );
   gpc1_1 gpc1403 (
      {stage2_56[9]},
      {stage3_56[7]}
   );
   gpc1_1 gpc1404 (
      {stage2_56[10]},
      {stage3_56[8]}
   );
   gpc1_1 gpc1405 (
      {stage2_56[11]},
      {stage3_56[9]}
   );
   gpc1_1 gpc1406 (
      {stage2_56[12]},
      {stage3_56[10]}
   );
   gpc1_1 gpc1407 (
      {stage2_59[3]},
      {stage3_59[4]}
   );
   gpc1_1 gpc1408 (
      {stage2_59[4]},
      {stage3_59[5]}
   );
   gpc1_1 gpc1409 (
      {stage2_59[5]},
      {stage3_59[6]}
   );
   gpc1_1 gpc1410 (
      {stage2_59[6]},
      {stage3_59[7]}
   );
   gpc1_1 gpc1411 (
      {stage2_59[7]},
      {stage3_59[8]}
   );
   gpc1_1 gpc1412 (
      {stage2_59[8]},
      {stage3_59[9]}
   );
   gpc1_1 gpc1413 (
      {stage2_59[9]},
      {stage3_59[10]}
   );
   gpc1_1 gpc1414 (
      {stage2_59[10]},
      {stage3_59[11]}
   );
   gpc1_1 gpc1415 (
      {stage2_59[11]},
      {stage3_59[12]}
   );
   gpc1_1 gpc1416 (
      {stage2_59[12]},
      {stage3_59[13]}
   );
   gpc1_1 gpc1417 (
      {stage2_61[6]},
      {stage3_61[4]}
   );
   gpc1_1 gpc1418 (
      {stage2_61[7]},
      {stage3_61[5]}
   );
   gpc1_1 gpc1419 (
      {stage2_61[8]},
      {stage3_61[6]}
   );
   gpc1_1 gpc1420 (
      {stage2_61[9]},
      {stage3_61[7]}
   );
   gpc1_1 gpc1421 (
      {stage2_61[10]},
      {stage3_61[8]}
   );
   gpc1_1 gpc1422 (
      {stage2_61[11]},
      {stage3_61[9]}
   );
   gpc1_1 gpc1423 (
      {stage2_63[12]},
      {stage3_63[5]}
   );
   gpc1_1 gpc1424 (
      {stage2_63[13]},
      {stage3_63[6]}
   );
   gpc1_1 gpc1425 (
      {stage2_63[14]},
      {stage3_63[7]}
   );
   gpc1_1 gpc1426 (
      {stage2_63[15]},
      {stage3_63[8]}
   );
   gpc1_1 gpc1427 (
      {stage2_63[16]},
      {stage3_63[9]}
   );
   gpc1_1 gpc1428 (
      {stage2_65[6]},
      {stage3_65[3]}
   );
   gpc1_1 gpc1429 (
      {stage2_65[7]},
      {stage3_65[4]}
   );
   gpc1_1 gpc1430 (
      {stage2_65[8]},
      {stage3_65[5]}
   );
   gpc1_1 gpc1431 (
      {stage2_65[9]},
      {stage3_65[6]}
   );
   gpc1_1 gpc1432 (
      {stage2_66[0]},
      {stage3_66[2]}
   );
   gpc1_1 gpc1433 (
      {stage2_66[1]},
      {stage3_66[3]}
   );
   gpc1_1 gpc1434 (
      {stage2_66[2]},
      {stage3_66[4]}
   );
   gpc1_1 gpc1435 (
      {stage2_66[3]},
      {stage3_66[5]}
   );
   gpc615_5 gpc1436 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4]},
      {stage3_3[0]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0]}
   );
   gpc615_5 gpc1437 (
      {stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage3_4[6]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[1],stage4_5[1],stage4_4[1],stage4_3[1]}
   );
   gpc2135_5 gpc1438 (
      {stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage3_5[6], stage3_5[7], stage3_5[8]},
      {stage3_6[0]},
      {stage3_7[0], stage3_7[1]},
      {stage4_8[0],stage4_7[1],stage4_6[2],stage4_5[2],stage4_4[2]}
   );
   gpc615_5 gpc1439 (
      {stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], 1'b0},
      {stage3_7[2]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[2],stage4_6[3]}
   );
   gpc615_5 gpc1440 (
      {stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7]},
      {stage3_8[6]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[1],stage4_9[1],stage4_8[2],stage4_7[3]}
   );
   gpc615_5 gpc1441 (
      {stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11], stage3_7[12]},
      {1'b0},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], 1'b0},
      {stage4_11[1],stage4_10[2],stage4_9[2],stage4_8[3],stage4_7[4]}
   );
   gpc7_3 gpc1442 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5], stage3_10[6]},
      {stage4_12[0],stage4_11[2],stage4_10[3]}
   );
   gpc135_4 gpc1443 (
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], 1'b0},
      {stage3_12[0], stage3_12[1], stage3_12[2]},
      {stage3_13[0]},
      {stage4_14[0],stage4_13[0],stage4_12[1],stage4_11[3]}
   );
   gpc207_4 gpc1444 (
      {stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5], stage3_13[6], stage3_13[7]},
      {stage3_15[0], stage3_15[1]},
      {stage4_16[0],stage4_15[0],stage4_14[1],stage4_13[1]}
   );
   gpc1415_5 gpc1445 (
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], 1'b0},
      {stage3_15[2]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3]},
      {stage3_17[0]},
      {stage4_18[0],stage4_17[0],stage4_16[1],stage4_15[1],stage4_14[2]}
   );
   gpc117_4 gpc1446 (
      {stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5], stage3_17[6], stage3_17[7]},
      {stage3_18[0]},
      {stage3_19[0]},
      {stage4_20[0],stage4_19[0],stage4_18[1],stage4_17[1]}
   );
   gpc1406_5 gpc1447 (
      {stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5], stage3_19[6]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3]},
      {stage3_22[0]},
      {stage4_23[0],stage4_22[0],stage4_21[0],stage4_20[1],stage4_19[1]}
   );
   gpc615_5 gpc1448 (
      {stage3_20[0], stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4]},
      {stage3_21[4]},
      {stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5], stage3_22[6]},
      {stage4_24[0],stage4_23[1],stage4_22[1],stage4_21[1],stage4_20[2]}
   );
   gpc615_5 gpc1449 (
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4]},
      {stage3_24[0]},
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5]},
      {stage4_27[0],stage4_26[0],stage4_25[0],stage4_24[1],stage4_23[2]}
   );
   gpc15_3 gpc1450 (
      {stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage3_25[6]},
      {stage4_26[1],stage4_25[1],stage4_24[2]}
   );
   gpc615_5 gpc1451 (
      {stage3_26[0], stage3_26[1], stage3_26[2], stage3_26[3], stage3_26[4]},
      {stage3_27[0]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], 1'b0},
      {stage4_30[0],stage4_29[0],stage4_28[0],stage4_27[1],stage4_26[2]}
   );
   gpc1163_5 gpc1452 (
      {stage3_29[0], stage3_29[1], stage3_29[2]},
      {stage3_30[0], stage3_30[1], stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5]},
      {stage3_31[0]},
      {stage3_32[0]},
      {stage4_33[0],stage4_32[0],stage4_31[0],stage4_30[1],stage4_29[1]}
   );
   gpc606_5 gpc1453 (
      {stage3_29[3], stage3_29[4], stage3_29[5], stage3_29[6], stage3_29[7], stage3_29[8]},
      {stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5], stage3_31[6]},
      {stage4_33[1],stage4_32[1],stage4_31[1],stage4_30[2],stage4_29[2]}
   );
   gpc3_2 gpc1454 (
      {stage3_32[1], stage3_32[2], stage3_32[3]},
      {stage4_33[2],stage4_32[2]}
   );
   gpc2135_5 gpc1455 (
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4]},
      {stage3_34[0], stage3_34[1], stage3_34[2]},
      {stage3_35[0]},
      {stage3_36[0], stage3_36[1]},
      {stage4_37[0],stage4_36[0],stage4_35[0],stage4_34[0],stage4_33[3]}
   );
   gpc2135_5 gpc1456 (
      {stage3_33[5], stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9]},
      {stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage3_35[1]},
      {stage3_36[2], stage3_36[3]},
      {stage4_37[1],stage4_36[1],stage4_35[1],stage4_34[1],stage4_33[4]}
   );
   gpc2135_5 gpc1457 (
      {stage3_33[10], stage3_33[11], stage3_33[12], stage3_33[13], stage3_33[14]},
      {stage3_34[6], stage3_34[7], stage3_34[8]},
      {stage3_35[2]},
      {stage3_36[4], stage3_36[5]},
      {stage4_37[2],stage4_36[2],stage4_35[2],stage4_34[2],stage4_33[5]}
   );
   gpc615_5 gpc1458 (
      {stage3_37[0], stage3_37[1], stage3_37[2], stage3_37[3], stage3_37[4]},
      {stage3_38[0]},
      {stage3_39[0], stage3_39[1], stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5]},
      {stage4_41[0],stage4_40[0],stage4_39[0],stage4_38[0],stage4_37[3]}
   );
   gpc2116_5 gpc1459 (
      {stage3_40[0], stage3_40[1], stage3_40[2], stage3_40[3], stage3_40[4], stage3_40[5]},
      {stage3_41[0]},
      {stage3_42[0]},
      {stage3_43[0], stage3_43[1]},
      {stage4_44[0],stage4_43[0],stage4_42[0],stage4_41[1],stage4_40[1]}
   );
   gpc207_4 gpc1460 (
      {stage3_41[1], stage3_41[2], stage3_41[3], stage3_41[4], stage3_41[5], stage3_41[6], 1'b0},
      {stage3_43[2], stage3_43[3]},
      {stage4_44[1],stage4_43[1],stage4_42[1],stage4_41[2]}
   );
   gpc2135_5 gpc1461 (
      {stage3_42[1], stage3_42[2], stage3_42[3], stage3_42[4], stage3_42[5]},
      {stage3_43[4], stage3_43[5], stage3_43[6]},
      {stage3_44[0]},
      {stage3_45[0], stage3_45[1]},
      {stage4_46[0],stage4_45[0],stage4_44[2],stage4_43[2],stage4_42[2]}
   );
   gpc2135_5 gpc1462 (
      {stage3_44[1], stage3_44[2], stage3_44[3], stage3_44[4], stage3_44[5]},
      {stage3_45[2], stage3_45[3], stage3_45[4]},
      {stage3_46[0]},
      {stage3_47[0], stage3_47[1]},
      {stage4_48[0],stage4_47[0],stage4_46[1],stage4_45[1],stage4_44[3]}
   );
   gpc615_5 gpc1463 (
      {stage3_46[1], stage3_46[2], stage3_46[3], stage3_46[4], stage3_46[5]},
      {stage3_47[2]},
      {stage3_48[0], stage3_48[1], stage3_48[2], stage3_48[3], stage3_48[4], stage3_48[5]},
      {stage4_50[0],stage4_49[0],stage4_48[1],stage4_47[1],stage4_46[2]}
   );
   gpc615_5 gpc1464 (
      {stage3_47[3], stage3_47[4], stage3_47[5], stage3_47[6], stage3_47[7]},
      {stage3_48[6]},
      {stage3_49[0], stage3_49[1], stage3_49[2], stage3_49[3], stage3_49[4], stage3_49[5]},
      {stage4_51[0],stage4_50[1],stage4_49[1],stage4_48[2],stage4_47[2]}
   );
   gpc606_5 gpc1465 (
      {stage3_48[7], stage3_48[8], stage3_48[9], stage3_48[10], stage3_48[11], stage3_48[12]},
      {stage3_50[0], stage3_50[1], stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5]},
      {stage4_52[0],stage4_51[1],stage4_50[2],stage4_49[2],stage4_48[3]}
   );
   gpc615_5 gpc1466 (
      {stage3_50[6], stage3_50[7], stage3_50[8], stage3_50[9], stage3_50[10]},
      {stage3_51[0]},
      {stage3_52[0], stage3_52[1], stage3_52[2], stage3_52[3], stage3_52[4], stage3_52[5]},
      {stage4_54[0],stage4_53[0],stage4_52[1],stage4_51[2],stage4_50[3]}
   );
   gpc606_5 gpc1467 (
      {stage3_51[1], stage3_51[2], stage3_51[3], stage3_51[4], stage3_51[5], stage3_51[6]},
      {stage3_53[0], stage3_53[1], stage3_53[2], stage3_53[3], stage3_53[4], stage3_53[5]},
      {stage4_55[0],stage4_54[1],stage4_53[1],stage4_52[2],stage4_51[3]}
   );
   gpc615_5 gpc1468 (
      {stage3_52[6], stage3_52[7], stage3_52[8], stage3_52[9], stage3_52[10]},
      {stage3_53[6]},
      {stage3_54[0], stage3_54[1], stage3_54[2], stage3_54[3], stage3_54[4], stage3_54[5]},
      {stage4_56[0],stage4_55[1],stage4_54[2],stage4_53[2],stage4_52[3]}
   );
   gpc1343_5 gpc1469 (
      {stage3_55[0], stage3_55[1], stage3_55[2]},
      {stage3_56[0], stage3_56[1], stage3_56[2], stage3_56[3]},
      {stage3_57[0], stage3_57[1], stage3_57[2]},
      {stage3_58[0]},
      {stage4_59[0],stage4_58[0],stage4_57[0],stage4_56[1],stage4_55[2]}
   );
   gpc1343_5 gpc1470 (
      {stage3_55[3], stage3_55[4], stage3_55[5]},
      {stage3_56[4], stage3_56[5], stage3_56[6], stage3_56[7]},
      {stage3_57[3], stage3_57[4], stage3_57[5]},
      {stage3_58[1]},
      {stage4_59[1],stage4_58[1],stage4_57[1],stage4_56[2],stage4_55[3]}
   );
   gpc623_5 gpc1471 (
      {stage3_57[6], stage3_57[7], 1'b0},
      {stage3_58[2], stage3_58[3]},
      {stage3_59[0], stage3_59[1], stage3_59[2], stage3_59[3], stage3_59[4], stage3_59[5]},
      {stage4_61[0],stage4_60[0],stage4_59[2],stage4_58[2],stage4_57[2]}
   );
   gpc606_5 gpc1472 (
      {stage3_59[6], stage3_59[7], stage3_59[8], stage3_59[9], stage3_59[10], stage3_59[11]},
      {stage3_61[0], stage3_61[1], stage3_61[2], stage3_61[3], stage3_61[4], stage3_61[5]},
      {stage4_63[0],stage4_62[0],stage4_61[1],stage4_60[1],stage4_59[3]}
   );
   gpc117_4 gpc1473 (
      {stage3_60[0], stage3_60[1], stage3_60[2], stage3_60[3], stage3_60[4], stage3_60[5], 1'b0},
      {stage3_61[6]},
      {stage3_62[0]},
      {stage4_63[1],stage4_62[1],stage4_61[2],stage4_60[2]}
   );
   gpc2223_5 gpc1474 (
      {stage3_62[1], stage3_62[2], stage3_62[3]},
      {stage3_63[0], stage3_63[1]},
      {stage3_64[0], stage3_64[1]},
      {stage3_65[0], stage3_65[1]},
      {stage4_66[0],stage4_65[0],stage4_64[0],stage4_63[2],stage4_62[2]}
   );
   gpc606_5 gpc1475 (
      {stage3_63[2], stage3_63[3], stage3_63[4], stage3_63[5], stage3_63[6], stage3_63[7]},
      {stage3_65[2], stage3_65[3], stage3_65[4], stage3_65[5], stage3_65[6], 1'b0},
      {stage4_67[0],stage4_66[1],stage4_65[1],stage4_64[1],stage4_63[3]}
   );
   gpc606_5 gpc1476 (
      {stage3_64[2], stage3_64[3], stage3_64[4], 1'b0, 1'b0, 1'b0},
      {stage3_66[0], stage3_66[1], stage3_66[2], stage3_66[3], stage3_66[4], stage3_66[5]},
      {stage4_68[0],stage4_67[1],stage4_66[2],stage4_65[2],stage4_64[2]}
   );
   gpc1_1 gpc1477 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc1478 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc1479 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc1480 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc1481 (
      {stage3_4[12]},
      {stage4_4[3]}
   );
   gpc1_1 gpc1482 (
      {stage3_4[13]},
      {stage4_4[4]}
   );
   gpc1_1 gpc1483 (
      {stage3_4[14]},
      {stage4_4[5]}
   );
   gpc1_1 gpc1484 (
      {stage3_7[13]},
      {stage4_7[5]}
   );
   gpc1_1 gpc1485 (
      {stage3_12[3]},
      {stage4_12[2]}
   );
   gpc1_1 gpc1486 (
      {stage3_12[4]},
      {stage4_12[3]}
   );
   gpc1_1 gpc1487 (
      {stage3_15[3]},
      {stage4_15[2]}
   );
   gpc1_1 gpc1488 (
      {stage3_15[4]},
      {stage4_15[3]}
   );
   gpc1_1 gpc1489 (
      {stage3_15[5]},
      {stage4_15[4]}
   );
   gpc1_1 gpc1490 (
      {stage3_16[4]},
      {stage4_16[2]}
   );
   gpc1_1 gpc1491 (
      {stage3_16[5]},
      {stage4_16[3]}
   );
   gpc1_1 gpc1492 (
      {stage3_18[1]},
      {stage4_18[2]}
   );
   gpc1_1 gpc1493 (
      {stage3_18[2]},
      {stage4_18[3]}
   );
   gpc1_1 gpc1494 (
      {stage3_18[3]},
      {stage4_18[4]}
   );
   gpc1_1 gpc1495 (
      {stage3_18[4]},
      {stage4_18[5]}
   );
   gpc1_1 gpc1496 (
      {stage3_18[5]},
      {stage4_18[6]}
   );
   gpc1_1 gpc1497 (
      {stage3_19[7]},
      {stage4_19[2]}
   );
   gpc1_1 gpc1498 (
      {stage3_21[5]},
      {stage4_21[2]}
   );
   gpc1_1 gpc1499 (
      {stage3_21[6]},
      {stage4_21[3]}
   );
   gpc1_1 gpc1500 (
      {stage3_25[7]},
      {stage4_25[2]}
   );
   gpc1_1 gpc1501 (
      {stage3_26[5]},
      {stage4_26[3]}
   );
   gpc1_1 gpc1502 (
      {stage3_27[1]},
      {stage4_27[2]}
   );
   gpc1_1 gpc1503 (
      {stage3_27[2]},
      {stage4_27[3]}
   );
   gpc1_1 gpc1504 (
      {stage3_27[3]},
      {stage4_27[4]}
   );
   gpc1_1 gpc1505 (
      {stage3_27[4]},
      {stage4_27[5]}
   );
   gpc1_1 gpc1506 (
      {stage3_29[9]},
      {stage4_29[3]}
   );
   gpc1_1 gpc1507 (
      {stage3_29[10]},
      {stage4_29[4]}
   );
   gpc1_1 gpc1508 (
      {stage3_29[11]},
      {stage4_29[5]}
   );
   gpc1_1 gpc1509 (
      {stage3_35[3]},
      {stage4_35[3]}
   );
   gpc1_1 gpc1510 (
      {stage3_37[5]},
      {stage4_37[4]}
   );
   gpc1_1 gpc1511 (
      {stage3_37[6]},
      {stage4_37[5]}
   );
   gpc1_1 gpc1512 (
      {stage3_38[1]},
      {stage4_38[1]}
   );
   gpc1_1 gpc1513 (
      {stage3_38[2]},
      {stage4_38[2]}
   );
   gpc1_1 gpc1514 (
      {stage3_38[3]},
      {stage4_38[3]}
   );
   gpc1_1 gpc1515 (
      {stage3_38[4]},
      {stage4_38[4]}
   );
   gpc1_1 gpc1516 (
      {stage3_38[5]},
      {stage4_38[5]}
   );
   gpc1_1 gpc1517 (
      {stage3_38[6]},
      {stage4_38[6]}
   );
   gpc1_1 gpc1518 (
      {stage3_40[6]},
      {stage4_40[2]}
   );
   gpc1_1 gpc1519 (
      {stage3_43[7]},
      {stage4_43[3]}
   );
   gpc1_1 gpc1520 (
      {stage3_44[6]},
      {stage4_44[4]}
   );
   gpc1_1 gpc1521 (
      {stage3_44[7]},
      {stage4_44[5]}
   );
   gpc1_1 gpc1522 (
      {stage3_47[8]},
      {stage4_47[3]}
   );
   gpc1_1 gpc1523 (
      {stage3_51[7]},
      {stage4_51[4]}
   );
   gpc1_1 gpc1524 (
      {stage3_56[8]},
      {stage4_56[3]}
   );
   gpc1_1 gpc1525 (
      {stage3_56[9]},
      {stage4_56[4]}
   );
   gpc1_1 gpc1526 (
      {stage3_56[10]},
      {stage4_56[5]}
   );
   gpc1_1 gpc1527 (
      {stage3_59[12]},
      {stage4_59[4]}
   );
   gpc1_1 gpc1528 (
      {stage3_59[13]},
      {stage4_59[5]}
   );
   gpc1_1 gpc1529 (
      {stage3_61[7]},
      {stage4_61[3]}
   );
   gpc1_1 gpc1530 (
      {stage3_61[8]},
      {stage4_61[4]}
   );
   gpc1_1 gpc1531 (
      {stage3_61[9]},
      {stage4_61[5]}
   );
   gpc1_1 gpc1532 (
      {stage3_63[8]},
      {stage4_63[4]}
   );
   gpc1_1 gpc1533 (
      {stage3_63[9]},
      {stage4_63[5]}
   );
   gpc1_1 gpc1534 (
      {stage3_67[0]},
      {stage4_67[2]}
   );
   gpc207_4 gpc1535 (
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5], 1'b0},
      {stage4_6[0], stage4_6[1]},
      {stage5_7[0],stage5_6[0],stage5_5[0],stage5_4[0]}
   );
   gpc623_5 gpc1536 (
      {stage4_5[0], stage4_5[1], stage4_5[2]},
      {stage4_6[2], stage4_6[3]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[0],stage5_7[1],stage5_6[1],stage5_5[1]}
   );
   gpc135_4 gpc1537 (
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], 1'b0},
      {stage4_9[0], stage4_9[1], stage4_9[2]},
      {stage4_10[0]},
      {stage5_11[0],stage5_10[0],stage5_9[1],stage5_8[1]}
   );
   gpc1343_5 gpc1538 (
      {stage4_10[1], stage4_10[2], stage4_10[3]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3]},
      {stage4_12[0], stage4_12[1], stage4_12[2]},
      {stage4_13[0]},
      {stage5_14[0],stage5_13[0],stage5_12[0],stage5_11[1],stage5_10[1]}
   );
   gpc1343_5 gpc1539 (
      {stage4_14[0], stage4_14[1], stage4_14[2]},
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3]},
      {stage4_16[0], stage4_16[1], stage4_16[2]},
      {stage4_17[0]},
      {stage5_18[0],stage5_17[0],stage5_16[0],stage5_15[0],stage5_14[1]}
   );
   gpc7_3 gpc1540 (
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5], stage4_18[6]},
      {stage5_20[0],stage5_19[0],stage5_18[1]}
   );
   gpc1343_5 gpc1541 (
      {stage4_19[0], stage4_19[1], stage4_19[2]},
      {stage4_20[0], stage4_20[1], stage4_20[2], 1'b0},
      {stage4_21[0], stage4_21[1], stage4_21[2]},
      {stage4_22[0]},
      {stage5_23[0],stage5_22[0],stage5_21[0],stage5_20[1],stage5_19[1]}
   );
   gpc23_3 gpc1542 (
      {stage4_23[0], stage4_23[1], stage4_23[2]},
      {stage4_24[0], stage4_24[1]},
      {stage5_25[0],stage5_24[0],stage5_23[1]}
   );
   gpc1343_5 gpc1543 (
      {stage4_24[2], 1'b0, 1'b0},
      {stage4_25[0], stage4_25[1], stage4_25[2], 1'b0},
      {stage4_26[0], stage4_26[1], stage4_26[2]},
      {stage4_27[0]},
      {stage5_28[0],stage5_27[0],stage5_26[0],stage5_25[1],stage5_24[1]}
   );
   gpc615_5 gpc1544 (
      {stage4_27[1], stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5]},
      {stage4_28[0]},
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage5_31[0],stage5_30[0],stage5_29[0],stage5_28[1],stage5_27[1]}
   );
   gpc223_4 gpc1545 (
      {stage4_30[0], stage4_30[1], stage4_30[2]},
      {stage4_31[0], stage4_31[1]},
      {stage4_32[0], stage4_32[1]},
      {stage5_33[0],stage5_32[0],stage5_31[1],stage5_30[1]}
   );
   gpc606_5 gpc1546 (
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], 1'b0, 1'b0},
      {stage5_37[0],stage5_36[0],stage5_35[0],stage5_34[0],stage5_33[1]}
   );
   gpc3_2 gpc1547 (
      {stage4_34[0], stage4_34[1], stage4_34[2]},
      {stage5_35[1],stage5_34[1]}
   );
   gpc1163_5 gpc1548 (
      {stage4_36[0], stage4_36[1], stage4_36[2]},
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], stage4_37[5]},
      {stage4_38[0]},
      {stage4_39[0]},
      {stage5_40[0],stage5_39[0],stage5_38[0],stage5_37[1],stage5_36[1]}
   );
   gpc606_5 gpc1549 (
      {stage4_38[1], stage4_38[2], stage4_38[3], stage4_38[4], stage4_38[5], stage4_38[6]},
      {stage4_40[0], stage4_40[1], stage4_40[2], 1'b0, 1'b0, 1'b0},
      {stage5_42[0],stage5_41[0],stage5_40[1],stage5_39[1],stage5_38[1]}
   );
   gpc1343_5 gpc1550 (
      {stage4_41[0], stage4_41[1], stage4_41[2]},
      {stage4_42[0], stage4_42[1], stage4_42[2], 1'b0},
      {stage4_43[0], stage4_43[1], stage4_43[2]},
      {stage4_44[0]},
      {stage5_45[0],stage5_44[0],stage5_43[0],stage5_42[1],stage5_41[1]}
   );
   gpc135_4 gpc1551 (
      {stage4_44[1], stage4_44[2], stage4_44[3], stage4_44[4], stage4_44[5]},
      {stage4_45[0], stage4_45[1], 1'b0},
      {stage4_46[0]},
      {stage5_47[0],stage5_46[0],stage5_45[1],stage5_44[1]}
   );
   gpc1343_5 gpc1552 (
      {stage4_46[1], stage4_46[2], 1'b0},
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3]},
      {stage4_48[0], stage4_48[1], stage4_48[2]},
      {stage4_49[0]},
      {stage5_50[0],stage5_49[0],stage5_48[0],stage5_47[1],stage5_46[1]}
   );
   gpc1343_5 gpc1553 (
      {stage4_49[1], stage4_49[2], 1'b0},
      {stage4_50[0], stage4_50[1], stage4_50[2], stage4_50[3]},
      {stage4_51[0], stage4_51[1], stage4_51[2]},
      {stage4_52[0]},
      {stage5_53[0],stage5_52[0],stage5_51[0],stage5_50[1],stage5_49[1]}
   );
   gpc1343_5 gpc1554 (
      {stage4_51[3], stage4_51[4], 1'b0},
      {stage4_52[1], stage4_52[2], stage4_52[3], 1'b0},
      {stage4_53[0], stage4_53[1], stage4_53[2]},
      {stage4_54[0]},
      {stage5_55[0],stage5_54[0],stage5_53[1],stage5_52[1],stage5_51[1]}
   );
   gpc1343_5 gpc1555 (
      {stage4_54[1], stage4_54[2], 1'b0},
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3]},
      {stage4_56[0], stage4_56[1], stage4_56[2]},
      {stage4_57[0]},
      {stage5_58[0],stage5_57[0],stage5_56[0],stage5_55[1],stage5_54[1]}
   );
   gpc1343_5 gpc1556 (
      {stage4_56[3], stage4_56[4], stage4_56[5]},
      {stage4_57[1], stage4_57[2], 1'b0, 1'b0},
      {stage4_58[0], stage4_58[1], stage4_58[2]},
      {stage4_59[0]},
      {stage5_60[0],stage5_59[0],stage5_58[1],stage5_57[1],stage5_56[1]}
   );
   gpc135_4 gpc1557 (
      {stage4_59[1], stage4_59[2], stage4_59[3], stage4_59[4], stage4_59[5]},
      {stage4_60[0], stage4_60[1], stage4_60[2]},
      {stage4_61[0]},
      {stage5_62[0],stage5_61[0],stage5_60[1],stage5_59[1]}
   );
   gpc2135_5 gpc1558 (
      {stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4], stage4_61[5]},
      {stage4_62[0], stage4_62[1], stage4_62[2]},
      {stage4_63[0]},
      {stage4_64[0], stage4_64[1]},
      {stage5_65[0],stage5_64[0],stage5_63[0],stage5_62[1],stage5_61[1]}
   );
   gpc615_5 gpc1559 (
      {stage4_63[1], stage4_63[2], stage4_63[3], stage4_63[4], stage4_63[5]},
      {stage4_64[2]},
      {stage4_65[0], stage4_65[1], stage4_65[2], 1'b0, 1'b0, 1'b0},
      {stage5_67[0],stage5_66[0],stage5_65[1],stage5_64[1],stage5_63[1]}
   );
   gpc2135_5 gpc1560 (
      {stage4_66[0], stage4_66[1], stage4_66[2], 1'b0, 1'b0},
      {stage4_67[0], stage4_67[1], stage4_67[2]},
      {stage4_68[0]},
      {1'b0, 1'b0},
      {stage5_69[0],stage5_68[0],stage5_67[1],stage5_66[1]}
   );
   gpc1_1 gpc1561 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc1562 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc1563 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc1564 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc1565 (
      {stage4_2[0]},
      {stage5_2[0]}
   );
   gpc1_1 gpc1566 (
      {stage4_3[0]},
      {stage5_3[0]}
   );
   gpc1_1 gpc1567 (
      {stage4_3[1]},
      {stage5_3[1]}
   );
   gpc1_1 gpc1568 (
      {stage4_12[3]},
      {stage5_12[1]}
   );
   gpc1_1 gpc1569 (
      {stage4_13[1]},
      {stage5_13[1]}
   );
   gpc1_1 gpc1570 (
      {stage4_15[4]},
      {stage5_15[1]}
   );
   gpc1_1 gpc1571 (
      {stage4_16[3]},
      {stage5_16[1]}
   );
   gpc1_1 gpc1572 (
      {stage4_17[1]},
      {stage5_17[1]}
   );
   gpc1_1 gpc1573 (
      {stage4_21[3]},
      {stage5_21[1]}
   );
   gpc1_1 gpc1574 (
      {stage4_22[1]},
      {stage5_22[1]}
   );
   gpc1_1 gpc1575 (
      {stage4_26[3]},
      {stage5_26[1]}
   );
   gpc1_1 gpc1576 (
      {stage4_32[2]},
      {stage5_32[1]}
   );
   gpc1_1 gpc1577 (
      {stage4_43[3]},
      {stage5_43[1]}
   );
   gpc1_1 gpc1578 (
      {stage4_48[3]},
      {stage5_48[1]}
   );
endmodule

module testbench();
    reg [53:0] src0;
    reg [53:0] src1;
    reg [53:0] src2;
    reg [53:0] src3;
    reg [53:0] src4;
    reg [53:0] src5;
    reg [53:0] src6;
    reg [53:0] src7;
    reg [53:0] src8;
    reg [53:0] src9;
    reg [53:0] src10;
    reg [53:0] src11;
    reg [53:0] src12;
    reg [53:0] src13;
    reg [53:0] src14;
    reg [53:0] src15;
    reg [53:0] src16;
    reg [53:0] src17;
    reg [53:0] src18;
    reg [53:0] src19;
    reg [53:0] src20;
    reg [53:0] src21;
    reg [53:0] src22;
    reg [53:0] src23;
    reg [53:0] src24;
    reg [53:0] src25;
    reg [53:0] src26;
    reg [53:0] src27;
    reg [53:0] src28;
    reg [53:0] src29;
    reg [53:0] src30;
    reg [53:0] src31;
    reg [53:0] src32;
    reg [53:0] src33;
    reg [53:0] src34;
    reg [53:0] src35;
    reg [53:0] src36;
    reg [53:0] src37;
    reg [53:0] src38;
    reg [53:0] src39;
    reg [53:0] src40;
    reg [53:0] src41;
    reg [53:0] src42;
    reg [53:0] src43;
    reg [53:0] src44;
    reg [53:0] src45;
    reg [53:0] src46;
    reg [53:0] src47;
    reg [53:0] src48;
    reg [53:0] src49;
    reg [53:0] src50;
    reg [53:0] src51;
    reg [53:0] src52;
    reg [53:0] src53;
    reg [53:0] src54;
    reg [53:0] src55;
    reg [53:0] src56;
    reg [53:0] src57;
    reg [53:0] src58;
    reg [53:0] src59;
    reg [53:0] src60;
    reg [53:0] src61;
    reg [53:0] src62;
    reg [53:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [69:0] srcsum;
    wire [69:0] dstsum;
    wire test;
    compressor_CLA54_64 compressor_CLA54_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h9b15ca35f6a3205889ce64aa9fb12fa967f1c59e9662e7b24ecdc5a59c34a73461aa428f3e0532afb0b6b03636f6ec345d3b19bca0b4c95934e3a3f50f8441a0611719aa1b4cf84eede600f5f0787acf9c5a95009a508aed73495bd9ea00ddcc409b59db46103f2e562285165a4ac6a0638bda699305aadaf06f2bf4bf8d9f5d9feeb8f907c93b2c522c784ea24b78efd53454dea7a302567ec44495f6ed21d7a7d7e1acf9bc6ee03185198d5ffad3b52e05ecf6813563baf0ac95af0ea61c05de22e89201098a389a168e5f5a7288330fd43eac45b76a326fa7e049e44b04e3604212c1d5607e36da6f2702334453abaf797c0573c2a4792e0dc02140a829a208edfa5d3c736977a151e8a8df636ad216a27069e6d23877b071fccc6dd520046564e17ebd9192ef149d4a9e4208942437c67eabc912a5f3a487fdf250690422ffca2ec1c07059729693efcf0ba032aaf26944cb49b71dc9886328c26448da4a3024bd5a0aad6f8915a43b8819613828f74e82a41b35f45370fd0c36104c768833e00fbdda2ce0761c6bba78de2016acd907ad5eb2ce5f952f98cda677cdc735d10bfbfe2cbfbf15279307a4900d9d08;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hf308fd6f8ffb0447d2bd3ff3cbc2ca5619cdead4bd2415f5d7c1b123bf9ba04beff800062e202cb65fb542eb73640368ebb9ac54e19f9c5a44545760d0e4921554491bc0289d110f594a88814350a74a6721bd43a0660f882a624a55e92dae1c6d181b3b444c57ac7d60d96ca1eb8821ccb3d04c446e5f22d661296ff14d68ace2fbdcec7a1fdfc4463d2c474889b40c68c6501529d8965f52625b88168d597e90b054fc1d65a92de58c647af294442d80b3c056d1fe6b7566aebe534c0b0bdeffaa8768ee4375c7eb6c0e14303d296fb6bfeb8a1e7e7b8027bb42de31a34cc76ffd3c82a548cac4ba610ab995988cc5a840705160795ac0fb55a424e7fa9fa8b3dbe6837fd53ad192a6d1a2402e04c04c352099d79b0413ed99ac8881f2c8690c7bb23ba1797204a8652dc3f1edfb6e0b96b3e356fa8a7e260ee03b5279255a89e1ad620b7e1620481c941f610811d97bd86c2c6cce2e1f41be19048d6f5eb71321560388effb60e8690ceac82b33d5449561a7fe3f22d78513e4d1545e00431c10a58c0d5c0e612f29393e47fcc1a13fe023c1aa4178628a189251aff8962f6717c25ed2c9631317b20842ec27bec2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'he19f5d68aab6719a0b99904686001691007efa31d04b0f4b3a5684431ae6d5549eb1dc33b4e1bcfa4a3dfcd03005ba0e5c5aadd475b7c88e90fda49795f865c611cbab6968d0a19ccee4d98b72b2e6f41326e18da3138de26f584531fd5161a04e73caa7006d817ee0816d06c08e68bcf90548005922e5e5ca87d546bf0197739992055fa1a9eb13cff9039d4a26dbc631413d6197cc54066564b3d83d7d33097dfeccf738f20e2c5031906504a73be26868a26eab4a3fd7e6504de75d2294c7214dfb5fbd062fdee7ea5915ec6e3ed5aa5e60ba6fbc4e9e13d6a182a76666e39065ff1bee7ba2eb6f2fce5b0b3ffcccac0a15461d8b2fc2b1c08a0eb36fc6bee596494c5e78c9876294b72fb2ba071abd9b8610dec669e6c42a044992a4efc992eb669ef842aeb8a4bc94aca5767be1ed3f600905bc4b655541b7379c7d4a880baf28540aa5463ea46f58d6cee5d31c55c1d94a0a58fe5e92991b00dfb16c810d512822895728de6aeb405206458cdd272f9262423ca7e5713dd8ef87b1f7f388c2ec7f9cdaadb086c463092ed3b3f8761aaa5d748352ab15d7c44cba94a5615af455e4979420d4ad8c36f350039823;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hf92fada5a75bc2682ae36789dd73fd03462bed194fcae2c4cdf4bf00abd65a1aea9392e8a32ed75542e272cf3810f00b3e60d2556fdbe11b26df6e91f3954aa362cdb3dafabb2cf429f4e5185711f640cacd8aa4965b736885e049483919933f5a0271cf80c164c706bb161b7b8c660519f3acd201827ee0461801685b6525c07a69224dfb5e2a8f28d05d248ff59f9e4b9ecac4d81c803fefa8f1611de195c74b1b0707b6214cb11a2393ed54d1e2a053a5b6bdfb7a3faca6d1e41abdd9bc0c7903c043fed2b47a682bf9dfc2b09a1e504628b0d486e8365371af1db7d47bc44cffe14f725387d9247cb2d107f6b1e4cd39f8c34b7349d5c337fcf75894d6c4151d4c96460c3bd3861b8a339cf004af43e77d5bac00e67ec938b83d111bea817a0ce090d6c6ad06ee0d086a1d0736d5a5bbadc8f3dd1cf3a698d580645972be7ca98bd4b9e7562af089bf26d514547e9e2d14826619f4f472e2057b29a03415d5a6689a6611ec3664d3eca0a158f5d9207d7852cedfbcb92474f559d0a4f563a5b07cfa729e95e5cdd3be4490c996618fe4ca2fa0d39f5dd79e65f67bafc5ad1b9b55433da9d95b8183af6d3d1b3593;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hf4e499461b866abeffe69945366979099190bad867734f6cb1fcfe130f3b87b6a479ccf3a18b3f96ca7eb8d47321c0353757b4ab99a1a4091fc56f73b871dc65cc1d7ca31bc38c37715207963d2fdf7f84389d81a3ccf14247b08ea8210ec92bf7adc5afd25214b971a8f1c6166a610352011c236366bd358e8748a41f2eb6e273a9a47f08f0fdeaa8e1718a88ced40639646336d4887057a9095e165098609a918eed5adc22e05003ebb9e5014e39edee95e7b9227d3ea0ce440102ec9adc0db592e39dc1b77814b336aba58c0267c35dabda2f549f4140024f0f8ecd22a1ee8a211a8de6bc6caf5ec6ccf2d599bb2db32d9352003001e03ee0bd141a68d635ea06733754d66534d0c4a5fb22e9133ab900a2e9e474777c7ec1bf5899022a4e202cdd1a3c6b2a05a21e14c8bd6b9ed25541ae51fce03c262b30cd80cf624361d72db994b84e6338c4b2069ecc4d21940f9ef281ca7b9ced8088b7823c34b118535d37782c3bfe63af978124cbd0779e7634da4cc9d456e865dac3a5e92d8ef0ae72d10e54eb6707cbace02701c6efa9f682949b82bad866bdf6fd2526b57cb1e4450a09abe80d882777e8f37bbdc6bd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hd32b81e47aef9c6deeb7c5e615fde1a143c41212b39ccd71e1e8e68e36f83d6a4950c4b2239d315b879d56a367ebe66529284c316347a892b5316542e321468b82536f9b218ad5eb9a40d80bbb33e7077421327c949fa3cbd00c510852700ffd8e2c055cd352060c23b21e4b090b7d3c70f2ff8f1eb42e9a1430256ea117e7723bb699ee2aa887ac90cdb70ce55991dd42591a0ce72faefaa7e72b2d2c02a8bff59fcd7f0747445624e6627448c367dd079ce7b14e21f4c1d0faaac440a54e280451b489f5ca9fa846e12396cb07aefa3f50952bd63fb1908178b7c2554e09f1edd9f285d4d547ecfbc6d9b7a81df887a17456aa7c5b15cda353210a7fae62eee90457eb57b28952219bac8977f5522438a4bdc45580872cc393cbf6195283cf8824be639d0d3fcca36362b3aa8d9affab47ef60b1e4bd202364b6cb55555b35205df8f5b3047afe531e22ca5c0709df7d99f84a5dc4e2d91b40d976c03a679d24fe1fb1e520b005dcb30735db9344b455cd51eb4eec5a1541367c6af491cb213865b76e2b6fdcb0995786dd280253c81898905d2713e96e6d4cabeec044a1c9bac14587923218f17bd7d44d0bdbbf19;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hc1ea0317c7a59d8298d3de98eba59d6e034328242c483d6fbad3f5f74c7c6799bb9c876d8f13ddc0ac183a02526e81595054302cce2283edfcc9fbdc59ee6158346fa03e694ef98dff24965f98dc8e0f5d81dccee31b1a691aa0c9cd951f8eecb22a86f14aa678511ae1d057130a2b5348b865c42e5a0f3d82f28ce139d1cc4ea9c2ac854bee58d61a1ad15ca8f1649af5950e7f824b47a44a2155ae200403b568a734653fc47f73eefe3c31f1f8f0caa024a9a49a9a8905ccfe5eaabebdb7800ad8f99eb3d304b144c434b74764612f7d5dd2d1831cddb6220a3cc6a638449f9b1737eff25693ce47f07d8557d0eff6af0c16fb3720135501821bab8cb6a9ba489a288f2ae3df5a0849188695cf43e0cfb36c65695d6b68370308f3de6506dc8fe1c81ba14ed7b0a161e207076c1d609f137436d59c1424972f8475a7766621f980bbf41d1a0f3645de0a96ba112457c689f0e5b7559fc3ea858df105ba0e54708dc3af8999bdbb399edb668c104211d76ba4083614d32e1d27cc1f88c72bec2240656d3169a0cc8339f4bb0c1d1949640c530a706c09bd8a27b7df51013b1a7c34c02aa255bf917c5de5f833a8b608;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hb577e6e1740db65e93605306c2b46aa299b5f07175ffe21324cae2fcd91a1c439be00f161cc37c1f1e25b5cf7b43275d6eae154b5cda6a4bf6d783dee11ee30dc5610ed2f465f43c6d3c658d1bb6b05795d9d530a3b5dd19ef72fcb8b87e8758cd776883f2c3fc2e4d6fdad119f732b48b7de3a99c55ac7fb3b89f0305c0f067f1fe37668d6392141d0016fe911312a53ccf4ec5dede2fee82c71b52d039e274a8ee75e7bdeab4a3d7a230aa9f1c29975175a5a61090124f193dc402641b8f0ba58bb0502408348d7bad8646f9b0f11d2110c55f140e4e8ed51923a241b9db64844ae5404a918c0ede93d6c073ba5d9bbce008263ecbe61d304e2c3908bd8a78f6f1427ce7577c2ad84bb06c6c580b425fb0ed2dad532c8b56c9ba60c80e0688fae1e5162fe8b87faa0f6cfe480e598af6c958bb1b2f7824f233120c9d733caf518c53a8c5b6c28c35e8c5697a4d548199a5e4d3624f00159e149f2650f279e4d016fda1758ee9d9fbac8ad34e53bfa20cbf57db1dd7bfb3ccaf386896917994c11f53ce7af4c764b17ba29fe824802b101bbc5061bb8f5ea17efc723eb511e25918a0de9859b7b14f2749f64d933bca;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h4c228157261828f20ff816c17d75a84fd9c0d3a10e6492f8ccdad53dbec208b2e776b81673f3b71201168ee8ad74908fd1aaa37342113fb530c76e9eaec54120bc58c89af56df99cdac9b857df52503a160bf4184a74d1df3b23167bc7f55ec2f1f1804fcbc07634a16405a6362820fba04531aae004d1f1ae3120ddc2e90099e3e6a0cfa4cc522f24cb6ca24faac04ff58dac50356d6a69ec2273393831e9c172e70285fbf706fcf4a8d42ccd547f71a8794daab80e796f1ea509df826f2a1bceb379a5b75764993898aa495820bbd8df33fefb422afb4ba48a99c127834e4b55ef69d2889cbb8f4046e3001f45a4c8fa7912b7ad09505253bec5f962a5cf44a04044b733865e8cc1c42da233a7f3def1f9c822f0a2bd820685d845aeed64acd61bf9cb747db90ae982d464c14fccaeab2484908ac552d2a1c88bb638de69e688d34ef24c97bca940a28ebf9dc1e46612c6facd06803d641a46ef3bcf14ed0e7cb2ac754a6d5472089a4fe1c81cc494240d328cf71f99bc9a478c0088fcddfc79ba9789491d701d434200f70d5a36bdc74dc8873bd54aeaea0610e3f2084084a4abf691389417bf09f661faa37134d3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'ha4d5a160c33c2a9941cc4d932f95eab57506925730e12edc3597ffcf71771dd8b44ffe7ba58be57afdcef60063b1a48e125217695733428316df496a8fb459bb0f0d3444c2be79c73868d3425ac9ce2fd325ae4bc31b5c8263fcb9e27f4378c67f9ff055f214ef150aed263c92f6ebf302387ab4121a509c0643e697fae5fe45f08480e2b9d88debe28e662045e8bef5cab1f14ca073e04acef48641c632847732dcb735f556dac3753676bebc893ce1724c70422c4ebcaabab878dd297534736fab6d3d6403028df5e00ffd797d3cceb21506a5368d07793bf2ed390169d99e55b57dc37e7e50d2d831fc762959fb3837404f46f8f9e958400d7eda56a8e0e8381888f75011b857fb4ef51f388a568bf51b788b773b66bc564f8943a9c1bb950635bb1631173b43e70cc0cbe7902f16139f66bd7f26eeee24309517695d0b56ec803ee225c3a282c49c03f66ffc4fb4626b11998c1c3f11fcff650c3595416e252881afce11f44334004565380d2e40a395a8e8feb0a83cd1270bf628b24cf480169e493fd562322d5f933d7fc169e3ad5fb89e5b9d3d225884e675175c470f2d3801fddcb997134fe2a5a06434e7e0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h382ecdf3919d257d593e5f1eea3e60e78e5c5916483e344049773ce64008fe4ce103732f404500a0c617d8ad925f9aea998c3aa879b1865cc29ce3f1513e1aa0453b30e88aa8defbd33772020b313df58722ca0bdfeb7545a3ed1d9cf8a9c54f8c32c73b149a76d245d3c482ad19e5bed810b58162ac356b62f3936b3093810f0f55cf3f541133e793efaf30bc64845572128bea89c9ab37db2e1121b65a356c9ba69e7b8a4f6c5e1502129fee7c381c24790a3e90d6e4180151c81ece9a5c01465c73f255389dd2d091f6511bf13526c540657f7f6749c348186552323366801b9379e580f43f7d3962c619cfc32ffcd7afcd1a0ad5d3e00e89c6eed6a707ec38d5786a51995e3dbda10710f0e1e6e5a6792b6c3d8618cf171a7e0868a08ae2845ab8d0cdcd3c4bf28ec94a847db9c8ea2750e0c4727e023d445edae900c3deb55c0e538c3c2b166e610fd631ea674a62628e65b9eeaa241e360bd670002dde8ddc3948e1cfdf3ea2cb01508580fa8f8d1ef6f5afcf25b7f15c1f937b4b9f3c01927a2188fa8a0ee7b5d64e646d2161825bb412cc22af19257dbc36a0c114e94d6259e340f5c1a5beb3b492269be1e2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h1207b1018991e6ce107f706d119060bb63eef40ebafd7bf7dbd7dad404e5f1eef69f36a9c286df75049c15d1bb91ff8b6e917e2593a6cc84e2636accd38e4563e912955ec2c68dd5cc929f8c25c7201452d927184a446f64b98cef8a4fd12646bcefa38328fecc748e717b39e4bb028542f5d82f2ce34988addb8de65b0c21895f62c1e9f4b4c3e741a9cc648c502d32f779a1a76ac03f0122a2167c93f70ddc6a6016f07e57afefd922794422b04f62bb2b40d18d73e0742569a0049a6105c3e1c44a59dfcdc4e3e11a6f6ffc3f131149d4ad6b6765db61f7abac023fbe7f234e4a81695f8c94c3636d3e5c8b8e1df5b61b276fb1e14304ecaba8364ce28db6ff4f5e4bf521cf85a1c5bef0511be13ae49f1e7f3794ad6cd684a81a3c77e5ca5419a63951a75d0ba98e4fe80702089820cf6cd223f21362db8a2b2ce7e8eeeb8f499d13b1335e248da378e15e7d77ecb10a7ac84a315b506a815baad55550c0b979906f0367b52df533c462d481f4e6ebdef2d18387e36fd57e84f6948d0bc71002e0c3666c6c289b8be435e6850fad4c1723067da039257dbe92b8ddf3954bbb5ec0d6a248e4e8a0ac61425302e7e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h7430ae39ac8d2c29eb92bcea18723e2f11c48ec9b8cff9d3fcf64b3baac15b69fa15a1e79062fd08fc5a387093cf7071e12d555765bba31a6215086cc99732b1761153ace1c7d03eaa410dc0380e93d1c92ac8b2c89028eb73786409a85cc70cc68e88f2ef439a4e00528e365141d0eeb03a97957596faf52ef27b684e05f684557efb7ce9d763c59c65285d3896e30b0d9265ff9f683ebea98c71869748ff898d0daac198e22ceeccfbdd626ea570f60b12c269581e53ef45d9931669c64f7ca67a6e45cb9ef547a65b970ee3adfcf0469d9241a91600f202fcc2d0991e5d3eff35b059d6434ce4442d94bb762d770b48c698aa39cf750bc22dbd0ab7ac00a8424a4345f1e47986985c3df08fad94f90e1ca1bc1cc5938b1860083be41b95a57c470ea4ad706d33ccfd9e6e960be20bc6695379361e04f37d2b119bc0607f777537704e7689241f447ed1086ff0cc0338ecb1b03b764a22d37ac57cf5d4e4d0f9e0719d7a4d58825da2a7a119f111be6f9c3ae15b0d6e7628e0c70abba77efbb13cd7a1f3e4ac31702d3c2c531e8505a70ea2f0779171927d23582ddc398740f46c7fc681fc49ac4cb5514a6513ca05;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h2ed561aa830d476d30ac47972d3187d2563bf0ca1c24536e83e495dfeeea3229605282de8a8eb685a32e92f8c2bcdde8d58df0d6a0c28ba7b50f1f56682ac17575222c24b8cb049921c257b060fdf51b43b63915550f185660216ad60a598c3a561da6932ad261bec0d15682024bf918b539965f6b5e45b4d89359d036b173bb9c9bc50087cb761d410f32ed4d3c4c9d57e37d110e35735963369672f91c5b4fbae69c2feeb299ed1f24e3c03886e933472e20e5fb8a6f39bc59e90474a190a6c62941017b33f56ce71df6ec767b9cf21cb82ca5618120eb8c4526b86adf958a33ffbef9b87878874f3d75e4fd936dec1c1575ee731b800490d16e4486ed074d35eb661709ad37c44c79c201018eac35e39f0b89799c6224efb84175065d8ed73281fa706cff8d4781b7a7c1fce976f9c9a0dd76978ee25fe473157a2475228644fe8434d175fc51aa47107220f58ce2be0dbe53245ab831d4c486cb0410c7ebe5eb7a81fb5a177b45e421d595f02bad7cf1f718a581a423113b72434a56462dc2f1a7fa1282af1e808445c50480b278354dce50bd60f6f52a92936b60db4f1ad411bb9b5cdd2ed1ade1b384f053eb32;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hc70ab1b96010fa1c3a1864ab434616369d6854f94a2a035d3ffd5e9b1d543e93e0687a15414d11a798353acdc49a8125af9ef0faf58b4ecd348dfd63fa3def40ef275ba595839d20ede57dd359e0515d22f58771af95fd982c911dc90585523f072063e5794e4fd4033c3fba48473caadf0b64e5ce2cbfd790d6f17ae62f4fa0e74ed819ffc75722637981c03e1ce3e8a2a070b77d174ea912f02a004379933739d304a788436b3a349ff98f60214cf4f7acf0ebd9bd281150b0ab95e8de40b0bbfb344e96c54afc52de854d9415492fe6f1bfa1fd98c067102cd0d73462b96b724bf6b88f6b53babbcee67ca16a0bfc99d8461f63d765176578581649004948c7a69a0569747795bde44a8ecd08173cebb0e4172f3e1c5f677736c89d78ec20e494817471937761db230add7bb68a68a6afed7e43445f737050fab4e29784cb07215d69ec7a1623943b284d837d63bfa6f939141363688ac4222d090c6a70363a41497e29abca59f08029d7e1e88b4f1b9716b750dc7fd4f6eaa5ba8d12982ec8c8edc068c4c6b8f685e9eef603c8387a70c39d286b21d3a533cf5cfc505ba087db0f2ec7f3472f4f957f688c73a7fb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h8f8c8264bd37bcc193a959b562f3284613ffd294e5b787a7ee4501a20e9ce2b947d0de649bf8f6842d2996f1f0638e6b42b2b7c1958d4b57e3b3e181f86baf52644f9b88f37ce619f848de40fafe6359168fd7edbb9b7ad3f95d81bb2ff41aac05f86975730596dc3d49085955438cd09749aae6a19afd8aadb59f9909ce627333124733343e09f817a9d2b95a8851a0216ac83e40ec364cf023c7820407e3748383911087ad010a73d19f9c36e06a3df86c5d669b1b8de9754ac2ea60587a001b1d1830318fecbeb001ff71e3bfe73ce45fb7e02a0ee67bf9a96f76fe21dddb466385cef0d581b41296005fdb727186f33ececb90632983782586f95ea560d6cb24ade57cd3a763fa0f3d8aa68316381f434d77715d0799cf278e190f5acf1e9c84d3ccbf8a510a7dfe283c1d7da98890693765aad276adfc99cca4ad62bb11d23ab90f0d33991adafb06560b1592e366c6e6ce4aad74a92d5f6c76d7a8d5b210d027feac0daf05eb4580fe660d6511a65cdc4e4ba83d8ee86e6e1860c5ce8fd0538fe6c55e0c1cd42d4b14266457d28c3ffe9fe926bdc25ca593dc84598563e62e5655224ea6fa4d65f2c611b0ee21;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'ha4bfa768a569e497d21daec146172f9ea442df0e9025d6afe0b88040c3f361c399bdbb52a4b415306e7e74ceb3f3fea64556f67ea9472f94b0ce827fbc92fb6816cd1b3bb4bb140729c16ba16e9d70df53d80611f3bae40ddfe9c09049e5d625aeda8b0b4a12bc45b8c4d59894224d2d1f6f720070bf45c9216719e81769ee9a3c45853e40b7a6020959b33a04cf7026fe52b21a1f8d5690b61d6ee5100c5ccb3f4248152ea515294c12f5ef15e7a5a3347de76dbd066ba9b183f830a5ceb90440f470f36275c2f383b339237dcb3e672763bdd40bb36a0f0edf9fbb8257a391b100f4c7ee2711eff0edd79af7f42f42c4e6e428e0a31a57f9ccb386385e3cde4d496dc6ad12c1f36299667deb9ac9be77fb07ee703a5b55ddc207ba77fde51f5163dcc732f9e3d38760a2d764e16084ad5bc8b904791166da080e686a17ff0f57730b7693ac1f193ecdaf02fb1f43afa2278eb8fbf5fe0a701be690014d7d6be072052fd9189998073f6137ddd5abf9d112fe3108b0b7f581d422a0a29caf1d7de3c3dde9d002caa4c132de9351748590fdeb881e1c5e6308d461617594e84fefd5cc7b6ab32680009cfbabb8fb1445;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h6e972340b13589af818bd34392e1b92eb2a145c0156e68115e5182bb903b20945e48f117f881d146d18b368a40265039659e5ed5bdf36907fec3037afcb02ed9bc089863cd9e0e02fc4c49e5a589eeb8d05d05f664cefcfff8740c3f907f907d9b4dff468385b8ae293b96ce25131ea6262c474bf25b3c25e4b39a706131ec3a90dd0bc888a8e99c322f88c1e1c8f8ad36df6022334e153176cb3fad1b79b0853721ae86ad6889f2708ac492a98c0b0eee351637122c3c94b6d3df985d73c2bc64523900c34abe818737d905e75ba32e1e7be9cf37cfcca5210d44238f0f20654160dd0a860abc5021fb7eea2ae9f9d554a78cdf46c1669a8d4d7550ca383ef0790147d6fb1f641ad58dc0dde92a8501127200a6265265c02bf4e830029cf1ed84450f6e37deba1268a2bd07ab98848e1c9c1d08099857879dab6075fabca5e0fe1e2651e9a10f121e0637ec68f56fa8df95514df6fb766098828f09eada8c8ef0c9fb3c116c34d821920a2282455cb449796b341dd33ab9045a0b9826c77fd05cf96a40cc345fdd6b07666ee6c1488d2b8e8479272d07174314ed48a09534e30d2c729d42f77ef57afbbbfbb964f0d9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h57cb489a45a5dc90f81bb9a4bdc33a216e844865cec4f083573976553afe28445c41d1b9994746887fdfc4c790f8d651cb351574903615ca86dfaf405d0628a9c2f194f2d5996fdc1b1ce2a5469fe95ca5e50a2b7e35597e0822dbaa694a2ca815c71a2d61682e8d777448551fa06979cd3284e45fd2f6e5bf6206ac0c4948799687f03b82ead70485a44025f3af8d7e2bcb1f55afc5124f69717ade7447b67040038aad91947f3e400881ba940f5f91cab0a13086ef417466d14f583bd3605ec9f01fd9ba6cbe927c878fc2801a05c5ff3cda372f842ae083561df802f295acb96f41f88095bb81ad1c0b10c601df19ccf124aa5e7a3a169adc120c1298e3c6e6b927cb96cbd3f29acb42e1c64dacf05dd9f3d54a55329dba11879578bdfa4acfbc9e77c86f773e3fff63af935146dbaf8f708c4d0365e7bbb09cb4640cee7fa0441fc7cdff0b75b7c89571cbaa265e6767a121d911c5b2abf026a57bc46c5a4caf62b014d888adbd3792c62dfb1a685df561bc751e39e347779029cc6896ed2e009b69c3d35c35bca69522adbab200d6fe973c139931ce4a702844c0e9859afc85cc24d40c6eff6637e756b578e724;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h71d430a4f6d69ee1b0f80d983adc24ecbaf3bf0f86346ee9b315c41bbcff38f0aebeaac5e5fcb9312f8f927db082ccf1a87b4d73314a4f39f6eff0a46f879f4610973833155b96016ac8001324d805b26a83617e1985e5b96cd8da9592d4f22ab5b505e9d5bdbb59e157cbaf15c9aae8cdbd6a97b182088408dfe41ad2e507a0bea801fd410f9dad00d2b55c00e337fc5d172aa1eca1493f2d9ddde73a8523c371f7718eaaaf04289030ac475f5cfae13eb0deba8828f70717bd29d85c6dd18eb769af170986a9e38cf087778a0f56ba290224ffd5bd93e2ac07304e44b7c257250a43487f4a197bab882c1c7a0aef3b5efbb1d11c93b5522ffda906cadb9f4be17addd23c24ea561d3c2ab7ae987906e1be4a7784687c55522faf0a3343aaaf2b04dede1d98b8f84a084401d41c7e36061fb587c739fb4213584afeee7b3e14442e8f3fbc84a6d7063c7b45f9b0aee3b2f817dafbf3352f80a5e3275fd77a897c6906a2769ac22a95fec4429b128c33680f3c13a943b5656ce4165428cdd5c0ef0bf393f32f7862d4b1f0e9e69f1beb742b9f6e028e82c26548d24ce095cddbb3e391523160da587403c32dcaf9c10e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hd401c2dc249c5386bd2775a49f43f45e1a400939a0f2330aa169b6ef376af167060d95b4af1e088934248addf534113f750da4bf12d211441764b7f871d12e66217a522d45815d8ed427c56e672886f104280cd1b00bbe5af5aff80b580bb8afcc834f35666ca45f6ba6a7e881603e9ee11bafe1b3a3ae3d218c2787ce0b73e82e2afb5dc85f738ff17f10ec074967e888e54262d18a5906f35cec3774a43c934eff93620a71b76343169a97bd7af566092751baad203a3e1dc18d46680271915493e3d72b950a55ca10138c85478a8134a2d171f0a1f8c76b2b374c07e4a8484d43196cc820405a814ff7616d3c04f39dd59b376fbd2528908a2f8f9cc2cfbcc24a730e5bb3342e521096f6a26b15bc42a5ee9dc7820fdfffcd12359e551c6d67d87a8ad89e81ea596362a44182330cbc81236a162c052c28617cfa0ba062298964caa06b932c3565d761685168551817dd96995d5649c8cc7ab477ca7264cdf6848dcf3b2976a43132097b452586c0889152b7436a71ecf275cf53cc7ad15626b0c19e06b1fdfaabdbc57ccb053e0378816a6692a843bb9ba32267b7985b81b3e37848c5eb992919c8a742cf9fe163;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'ha073bb547ba2bb11757a84e47fefbeab4447a645453ff693b4fae78429923354f3a89369389696d1c5524a9e91c292664585e21a5b6e9563d03206a61dffe05d6bf4654533b47c671be24a5d6d8140f073655ae314b236df52fc446b7409813b71017b614ee319331f87a807fdf6a5bde365e92c59b25ae59441a0bead53b044c208a9a74bc29351b1817a9b5bfb6c2eb3e4fc6e1b15ba0c9e59245cde8016b312c3947ca1de1a9d649545f865412cbad22094ee63c34599c547990dd5c105778f85d19c33c33bef00c5cd7dc7e1526dd003278eddeee3fe1a8b893883054d1a76306aba784c067ffb027132a26261e492d4ac891bafacbb9bcd252c18caebb34ba58ae9071a03bafdf6a986e37a7ed08f24e875f10e8b5aef5f22399da91eb5f9e418cf63e5098635977907aab0f871114fc0bdc0d00d1214cd1db48c7a3b414ad3398f945bcc45dd6a68679a880efd55f7f3b07a28dce166d0938cca4f4208bc60324b94d55d602597faff33f48051c995c9b273a1cc4c8285093274f7ef94d0a94ff8f9a69ea0cc88ed3e9b6cd34ee1ef0e69f2ad0458af78098e6dc513dbdffcdc5ade3b07fa5e7ca228ab844257;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h49595e92c1d2349d682ab26ebc5fb0fc8e3689207e2be22ed8c13c660bd34a7130c20386ca3ec0f753dc7f0b032d5498660e0156f90d4c9b17c25c9388f4c7a0c6042361ac396df1261a6fc014b4a2e284be7b4abd6b5cc0bda5e2b21b4ad94c8ae783fb702600b1ff81947512de942ecbf8a67eec14ccfd85890894ad876f3369c5a746bcf1750dff1a07706336d43b50b5eaf7c6f1fa7c70bf72992d598ad2b5fc8cd2de74e25ad328c8be9c7df800cb736c27cd94af1fdccbbe0ff547aa0dc03c505beb459f8e8172ff7665ed72c5d13034bdf5f3f1c78b5ce4a39dbc950d15720f4aea85f08bc0f1848c092acb864cfa654336b2b71c15a0c2c03bdc9c22afb13a33d137522659ede3d3cb0963b5d81367c8da8a12ac322c553255d6ef5db3364d2e0573bb34af4130a91cc15f168b807763fe3cad3c7558aad6a7d5288119d51d8adfed86cec0feab73fb4c6a7b203a3b8c6969c527bf1cc72d91b9dabfd747d8d23869ee2215004c54a9387228de06195301aa5cc9c2615a6450c2c38dad7b406658287284f49dc1f406361a25a70acd8e991dcfe488378eebb54092aff4ef4e05bde744caa76367279f8ff6a2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h8b110a0b13a8ec5edae4eb7b962382ec425fde503c769bb98abadfefd20e8ce377c3cc64e0abb1233d0659f5d12d72979a327401414aa2d9974e3e4f5671ef4342e9e3f64b323f83eb603aabc5619e4bd8e004b29daef257aaaccc3af8ce2b7d0aed61af806f821cd0070f0c611eef8ea00f06ca83c23f4ab9b1337f0e85081b6707f3969a8b93575c14b3915a9cfc735466aed365f9c220c960c58430241c9e71c38e69639a33733b60c1c085e8c9c8b64f185e350341f7d88372a99850983c5ac2b879de8f2a234930315106d29e86000f0c5260fb812d775651604a37ffb04e7b0760109b91f652f4e7004073d880d2ef32095607c2a138e1edfe2f81e8fd45a73ea253d2bd78a1f19d920d72e01073c255ea67a5cdfc23d1f082578e1c9064b0be7af3ec823381e3d32a333315a2483c9de5c7a906ee004bfc4434201732b9077350e83e35ea1af1a99d3181979218aa7bb68974a48d9c8035e7ee2c7a56abb758ac1b9d9c32a8d13823e9dc92e9ba56beb5aea6b0f729fd21160650f5ddcea1ac2d98e7680ad829e5c7c044c166d2d7c6eaf498a6b5f3002b071c54bc76d8f20eba068ee5655e016b5d512bd550;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h9806c6820e6fe40f095ce8c3e9f7c4ecff46be15264a1abfa582806998c004b329793eecc4c1b6abb746240f1beedbe7a6d461612f68606ecbe862c2f992ccb2c37f47d512b611c2182286c623333f6318852895175bc601fc5769a71af8a19dd005161fe8253ebcdf8f83ca19dff1fb64e80c943fb6099d2d2fa18ee9e087d03e79ac3e9cdd6d63197f555826e0b1c4e992da4ab1e782a3b9d2e5bc26fca2534af609a0a02cf70d6e2cf6d237dea82cfc9a556da3783d090343a56af108f06ab87bf4b7b4b510203e2d4b5d84c7c9422edf4fda8aa7def7b82aecf661cb242781a97e171d16be7a9d26005e4906129bb3ddd90c152cb9aae294a54cbbee2847ad40e23db57955d87595308cad5e6bd4257352a8cf79338b640712ae727d8cebf7dfac818f89bf271e115a5b25a5c8b5a9b30f29c32efcc972c3226f4eb1033da0838a51fe62e743d2b0842fcafa81073d2ddba67e10c31e51521096178f9cb4f3251d2a3ebfc124442c949f9b576bf49d31e522143e4c29b1d9e63d1f6f85169b63703b3f9c8736f31aa7753352d2124d1897d4d94d3c2c308f25a8b8648239002787c62937011ea957f85af58092cc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h3b3522c36b5ce75375523b776371bd3e402b1f92003c4ed48a2841f3f5b418993985ff3643c1a15b83919fe06612368cc5880694f841fd030006ae25bec1e08c44e840683376114f381f5428d327b100771548a9128c48a64247f042f7cd9d18fbefdf49c9871c6cc2802acf8ca1fd353f35a7737c2103fe6466f7a72596fc168a72e4c01994f32e3ee418c988bb8d2bdfc6f8fd51e11c5f4110c1477ad6e84bb9c9f973200596a6f5ce09769d98b7cfb0511c738b18f2de8a9c603483fa9f26be4f79f75dc1498c182a024238fb9fcdea5d5480868a40b6bd695b815d56a581b3b189e20ac51798a75b1ce0b60c27e17c2ac6aea98471fe5dff38cbfa99e8aae746a76eb46572df05273bbf8f6567c2a984a38be9e252128d3988f7bf368c982f7c574a26913d0e2cbe671b5f70e5a9f1e2329200a7cd2d577c468cb7a0879e63b7055ee24529c309e3777e2f32f11e4def1cbee812f9987d92adfb3a57a4f8fd03a39440c1db4f1d33b28fb55dc532153f97f9494d5c03a38fe552fc238460f7953856bf7155cc7086524370eddc7f35ce8b1ac423a8561fe9ffd51c7a827052c9a4bce62925c87d54059a2c3fe5d2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h5aae6a12bc8a05ff91c0ce3bc96fc88e71b84e73b7243d407d33e023b8ab6a698568eedc22be69dec05df05d3fd90f84c266edc222dc105c649beca985088974df80024e1d4050a5d79a79c3b5e0a5c5dec404fdd3d446b3035d037fb1f01381451b9706104781768a2fcf080a0719fc6774d0efa1b5ba761c63dcb17371e0a87989ebb8917442fb1ca416881acb2c54bcd094ca86f6b74430475c4cc702efb7c19f5f3b26e1a039e04082a34141bcf7a19513027edcf71afbcab570d00b6ac88ea0a6bb8661c9a0ca5567657c85b37d3fef58efcba0a1535cfa6c10f90ae629441b514b9f08f81423a450fe9d0373386c0cf95881febf08c31b20e1738f11df312c0a4af5efa5655178a3d08fa29035af34c86e4dabeba876e2009d8d336a43da607b93a522614c63200cc7b094c6abce6b509ce4fac748ce6f92e77dcaf836d71ce17e33c75d3b4407f0ea0ce9f647330f34f0669c377d11f51d73f50b6c5b907dd98cb1cd101422534b9d67fa229fdaab8a54fb0d697ed5f45c1491d881115df2787dc525a5c49e4cbd40b74f74749eec74c10d415e1b4351ca06f67a46f6af6e9ae62c31b16fae4b1d3d33ca1afc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h808b1487ffd085e6927a63db16c058b64603c1d6d2a5557687e06b83a9d0803d778d3fe3a61324efc5a8e4446417f591d8b8a61a3ecaac240120a695d963eeab3bbfadd5f0e9830942f6fb7f35d37c618d0a5176355fbfa67e34300467963b5fa1489c2bc949dc67d34025a82d5c2a360ba4088c65d4111e95746bb124fe6ad6f543e67203f3446b11192625ffd2efec568d90cd285b31ec22fece05ab246e385fb824c691fffd00aec8592ec24b78e1db26bff7553428e4a637dd48717fd28720abdba761752163373b8f6c173b9877504e41d7bebd2604b61f5a7b78b87a1c5ef65adc7ab4381d272931bc3b34c53a46fdb1aa2c10697fe8ecfb14db9ee802e609bc7926f955b6b11792ef051a28fa12c176bab00941276f72c948c1850480cbdb842e6fcaeb0ea0466456df50fcd6ebf1fbd1f2953227f17432fbff8e976c8197a2df55a2a8b678775b840433d2fd2cfd19a23ef724d04dd7d1cfd7fead93c49f8c805429137ccaa12bf0befa1202e8e1e0b127fbbab9497f545206794c0c5dc2f630dbc05f7f2cc893d76175c6d28eb8c70b41a2b7f578f36f564c17872ad868d80dd522ca9bf1af6edb64ab9ade;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h27e85c5c3928e92184419b57d1da991c8d36da38854e0e8b6e955a30f53e44034309ccf44abe5df8bbc4a508a934f4a881b62a83e7ef3cf5dc4607886f9d6f5a2f76e0198ff1116600988f359cbb84dffc83a041565e05010b3b4b4988e23ef9b160f8bdb9e01fb1c9fbeb47c1ef76df8dbc3650f8c7d541fabbfb7b4d34887a933238c2803aafd6ce483d4ef1bf698a0f92f747099d4abc144ba6bbb606673bb0a9093a3ae67206fe5925c5c51f9b5afa88dad8453b6950974eb0a3a38764b152063d2f6d23f7e88afbe07572925f95aa3d8a67fba330ed411f474643daec068975579865e407f10b3d159a20655618b73ac6e46a835144c3d4dab5ca63c7b8ccda573e6285cbd49685ef75aeef99ecfa855be7dea4cc0e56d89d91f5be4bc9374e922fcbb21fb980f462a568b23892585556eac9efe38bcd94dec73509751976397f2552a8d42550dce3278c7d020790b87fcaa4c4230f0a63fae58cff93e94100f86024c005c2da8696b27434be9ea1ee5e6066067760e72fe0df3e41b211a8974d7c3389783be0d00c6020e517068f54af5e0987964b078995830dc8ff8da06253aa4ba6d22783a266b3334de292;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h38b137b23e270de42954c0cab85c5c4c0b16023b80fda407b4f3ad6136827980a20bf952a06c58f129655924bb1c48e527bf199c1a44c8a407412bd7fc679147fc8d2c4f7df3daa7fa04921233c0fda3cbd844b1d79e6ae95e99d6fcf50d5271b97ef62d44688ddbee73b1086bd5bdae86567506ceeda6f344b45ab26711f242095b1506f302b4c801077fb8cd607e9a013dab8e2f162da9cc79a97ad200742f40403f624a3d78f38a4285db1f950ddde45cdf39e4f0247a57d0680dc8d7c1e5f6e683a5d59f300d8ae4d69b03a8c66339449f3c6024733a985422fd817e210a88c8c22199ff3325a4d1e2c4d9f3163c06786b98edc44ab1b90fa8491cdc72d9ecf61af4874a75c4a8d252126165bad93bededc622c8dc4eccfc8cfe7a332bb2a509cb0ac768db2782c647ff91d3775c66e9225e58ac0abe1afdb8e6310d2283ef531d6bec8d13648a8034212d056650371c718e8b4c3af480ec1e27a5771e22b388525913bd0aaaaba9083e6f2458c2299b445b221a34fc6582e52dd33cdc33b02a3d213ea2fe037913f1aae1ffe0ec12449de4937f7b23cafdd0e74609b52bcdfef74064e2049941491238fd73dbc7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h28ec648061afc3fb0970ddeb4dba629a63893c16c3ec1b391b18fc6a3ba8151944f2c0d0fbae7f93f6e565b3aa59b3614bbeec615bc7c2a2ef364b32b6580f9d3bdfeef59e513380f385891fdcaecd9454175a2ed90e4aca25f1a47f4d70c6994061bf2957b409abdc28fed856b03ac30f9ce72f6d6a931727ed34065ab7f71c25d4a42deed424ffd1272bed2b018776e7bf83a6dc5539046c2652930fc49d2a88615c1afe830f9fcf5d7a85521532dec292e773767605bbf0e863db19438a3e6968de909a477eeecc06fe6432ec40961bbe6b02a801d6e0390d6451157fcd9afeb89db55bb7f2dda32b21f3fa1433f3e77f1b8b6a907a466559aaeb036376af99cf52ac586e8e2b464628bec56b4eb40ede77f8a85d24da43bc9d1598352776d44eedbc8be4edc0f3309edb06e55db95ac58aab8af56036ac49ea2ff322250a1cd444e4cf203e811c07c7da0d15ec9cfbee44968aca5d4c3cae4d00e3fa1cef2ab84b3c61f0b1c4993433de62243c7902f2bb590a621f79b45d98f9d8abfd6308969af1124f8be8368016e1fa1ecc8c1b70c679d494d2cbb860abb56281b38caf290d917649a836b0ba953f9f9496c5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hadd513f5dea46a3c84bc91a5b5ea6dc7166a3a915243f0a473fc55ab79b753c7dc65ba013e4aa3efc976fb727af8a5ac0eb519c23539c3e9aae25e8f5d24417dc12e58023e4f22c1221f94ba3347542b683feab2bf0cd351805b21a9c62ae88f884013bea969e2bc0a27c70a503fdd3ea2135b1567f826d347eb0a3f0e9f554e2ebe83629dbf5b5d594c87fec0d1892c891555902c889cd68142b0937e87e47213571efb722b825b61a841d7b03b0b20e77865526564bf97b0e53fb5bbc125ae1275ea6b501783d177ee8e8b73cca63265340d697cfe9c46cded3b8927a89dda68df022df6147b1bb3b721a985e36ca3f28498a790023f2e2e6964b92cf626f638aed71ba2b39893859ae13f0056ec3fa178d8d35bd8e817a3efa80ce9c7a8288c4a1b87c24c03256c04fa4649d94f568307a8b3fc14fe73d020c81b2c3a05b02601b41b17c1d5e1df8b365d7355ec30bd6d3cfd6a65a95690052fadf1466870fd5b10bdfdb4f9335ec6aa025b47cabce575903e83634611ba093888fc6471012dd9ea2e76edad35dea198afbb6b8b705fde5231ed57d238589e9775cd1187d8447bcc402a141d45d1b8e1420466e0c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h877ec144791e5f8357d0221fdbadb36fefaea8b10b1b1f373f0124b3e7ed223be4ca01d729bab143fbe07040fb58c7a4dac00a0afce689385f04da9f38a360d8437857af83965ec00f3f2e97f1e29191315a326978f4bb770e24674577bb0b74a42fbcae47f2ff8119cbd9ba99c4fb3b0f05c9fe7eda5a143dbfadd32420c35147c4115a45262f7f41ffc3fb3c9ec86d394f3aff10f0829020ea21890002aacf4e0eee7303416a8cbf5f5801c460c520fb6624a29f4dcb9ed38c2100e9d25641f87722b74c0a3b05d01cd04def42504649de840e3492ea7abc6d8767b35cf41a8afb8956d1efe1e6b888b4a1bc48d76b1dfc2b869a77147048cbd8742645b819e6d1297f1bec45cfdb02e9ef2c19e3d75bc66d83eb60d5054e2e363fcd673fd3c1fff1fdfd1e13e305620e37aeb61c011cdfcb50b2d86404a5279855769b6a570f4d208bd1ddf62aa10fd2a8105dfad7179eb21b1d96b1c7e6a686eb6e5e46765c89d8b65d7e5c036d6164b357e284cf9ba99aa4dae45ec0559b65f02e5b73e93e4b7bbae571ccc2f75fd3903238795aaa72d0ffee54bd5f953edf251d1562d97ac2e816170d31e19baddb952ef9154;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h2a40bca3d594f6c86b23e7a210c33dc6622ee49869bd60216cd2b2c653ef6a3892ec4f3b8a7424f2b8b6281bdc8c2889b1af1c935a26bec98ecf748f0db453772ea3911e841100731e06d9acb08980a1901caef777922241cf066e4eed38d66e4e1de818b6853dc83bbcc2528f63e75bfb5ce2a4b128f44d820ab011385760003f98bfe78405df273e20b7c9b933075bb1a135457c2124b26ce7967e7f2b1d3125abaec299f2964da2e6f521b597f55ed0d9f0005dee5a4833b7b802bd95438e57d2dab18293a73d0f48eecc89b5213bda268c8d814a9e3cae4c4c109c0107e7d46c9310428a0e31293054559592f868568c627f2a6b6c58d3c1d888d82678d3e509f1193b46df586fc9ce4da9f0f7073275509a9b0eba2467a5aab416be187e8d7a83cbec80ddcbbf0d0607adf64263324aa61575a27bd38c97324e80369a84b0602aef21f0c4bd2f78011e8decabf20eecce5bde991f58bc2fd211b5f13646f0c66ee82ae77538cf657d8e060ad5c0b71598bc457a948e5a50bf3c531394cb8aac979141e5084717d2b701d756a57d243b7a1057dd6365628dac3ab13bed20723123b0d88c31754a64bfd165bd4348;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h7caa504dad2da7e6b6688cdff282c6991da64dd82254eada60f9e94ec0c73de4723c782adb123eb7551743b89b4d5b331db6fbc98c6a24c947f4d4c38b29ced25874b26ca5f156211096ee2ba94edcf6f6501489eb198d9b0cd05242f3d0535f6219f8c9e7240c5b6860a0e34cec46c8ce28850d5397ae9df1e0405503b11239f6af46ee405abced882d47cfb32462e114121cf3e4dd66d4f091832bff3857636fa9d23a8b879adc7695acc0fa94cc6ccdf4645d9df64411aeb095d19a6e91db7284d24cdac1d61dcb25af06fc802d5fe77a4c3395d063f91bd9f7467d0ddc2200bb74c3c51c23eeb37e858fc9b882d303e0235ef90f4647b590a6f4ef392c50886c4c15c872e523dcc4f643ca7737c06423126cf68e6ed88e60c89858fea1cd6268547bcac7bf7b36e431519f4589485602ec6d0f3f3e1e914654b088a152a475a71c7c4686bf7df2100762dfec18077c330d8a589e5461d9ba6807c31ec5c8fdbfbd2fda54930db1d62a6526a419165cade81486e4d426ffd413d449822bfac8c981d7abe17892f1c351f84d9d413b1be057d363edc11b381b1d04d92066f825b3a2fecacd10450b2eff02d76c56fd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h85e681df479d3256e31640ce204ac73d1c92b0849d1a3ff71e5504c6d7bc64ab1aa5c5e7f3f41aaa34b294db43db6a1eaed5e46c19da6d4ed6504a7976140b78ff171fc5e519775a2b5784835f89b08315d7ec2db48fe4bbc8a479e534f6aeaf741b9d8ea8e11968a3a780b1b5036d8ce0d2f4843f30f9544851b50660fda6364354807e0969c0432b9dcc1c62051568c2ec2a39c79872ab636300397b4750b545a2cb3252bb87fa65b46c47918e20bb06fed65bc6bcf3c86f8bf40e8435b53b9dde0decadd6c473f4218e7d15f85fa001fafba14f772203de00cbc73ea20ce0e1b78a6fb89a5103e3810a75ef74b7097b7100649da180e134c5fdc00f03e2286a29b49aeec66b39ec0b64d0aac1368b0b59ce5aa5593b9de8d0d705a0754795d0cbeeb6ac72cf7f56c9fa93e8b51279ae38f6d8d0a0a9f6e031b6ff016241b3289928325a05239ecd33f7d8418a661614a2b6006915902c95e395517887de01e7d5b55f755d7b930b70aa4f2814c089e430630d15c5fc4fbed56ce84b5969a95f61c8e33300835f936580cbcf952ed356d60e278653426acbdfdaafd6e1a90a171691f782e15001c0d125c44c808437;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h898d3e8c15c8378a770f9b6392b8e72d9f5e20385c7665718fcf4108fc0e7ed140a4f9855058ac41638c66e0b76a4a316fe439686d6597527e00c318e1ea5cb9e04cc4bb5865faa8d43854a0de95857308999748acafef37359e7c667c2d65689695dab2362418990e3fd58af35bb3e44c6984d1c697baeddaa6990898f95bed4aa3364fc1dfd8ee870afab406abc894b6c887df7fd345e6121a17180f52cae6d7f88b6968aa3f292b2a85e49481c6b4e61391f165abb2107ae15178602bd7478962564722e9984072b5f46ef5e426b58bfa2d4aa09dde006a24f75c105546a3fecbe76c42ca4b53af99b3bc7a54fc84661872e4dd56413488aa596ebb114d6a61f75d02a3cb4d3945504fc5afce12d54f912e9f111a3423ea04c1e49d37fd74186be2a1e2f1f87e0e8d3ce1acbedd0637f0e502a88f14e68da4cb243cdf2c9b3714722ac5eebd97f6c4102df6d7ac267a8c5f067203b262918b5745156d44444a40f1ab2ba714fd8399150d36699c91a59b93b7ee526f03bd689721f128da61b53d1025e240122d69716080c4012a90f39406ff9fc168b88c492ce63b1fbfbbab53d15f17c739de335260eea65830bb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h73d451db566a279654b342441f384731651ef13f085e6138379d14aed3daf8fd6a3ae14b77c1b2506bea790c0ba7a14b1d5f110a70a968b42b1ce2fbd32d219ae943c45992008ac8cfa1e9216a5ee9a0784b96d762750b12344130963fc86aac391a2fde53291eadefac439cd4d333a22549a8adae6a955e0dca049eddc7c81b53a58886844a51a00d0cf2ef23584be968718f0bcef5068b9a91ed230c76852b3995cd67fa8f2b858f35b3a0143a965cdc999ff7e38eff6f5fecc259ad90973f708b110fb140a37bdd03d8a0ca4a656488cac4d6f1b1373c106bbaaa627675fbf337d42e545fb17ee635b6124bffd258b9da0818652b9057b02389752c5b7a57c7faeb78bdb5f8040669d640de93488f1415ab7be9305cb16d5d2cdd7ac1ae7df18000976b59b3d836fd291a3086043177a42659ef1324980ff6d4ab26619561b4da1787991577744474f238a44ae88137a9f415e36e3f61f78e595d595dfbee46298770175e214c705e4fd9236cbeb10674e3cf295310b442352ce54ec04e246c80220c974b6574611a355b301ebb98283e350767830440996c003af25c43728c0373cdc797a3d4dc08f3426030b76e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hd2c8b3746fc32f4e5788dcb75647b07ce965acff1a768392e1a77f5c03ed95ce2cc559a76de773b7199dea45221394db6042c88aae32ef16e2cbbc7f3a8cf6da9839647aa62de78cddcc91ddd629ea5f3ec9643448b85a63519ecda210d9bc9d69b2679097fb0b6929263c56f2c8f845a66c8fe085d691969d3bb89e01c6ad7736a5806a39fcaaa183a528b29072ee844c02c4f50937fffa7836f37828adbfba9a013f86c8e3d35fffacc917d2450c0382f05b29b029abbebfc34128851f5d2dc398cd58a96a1d1c5f0955b8bcf8c04cec702e3ed9b657a1d274e8e6b036bc874381393e72883881d84d99959687c307db6dd7de9c1f6ea863058ae21fb881dcee6f161cb129ddb712453a20b385dea6d76cffec3203af674b7d147f666d014ff439d2ab1d1bd8997b82915bcdbab73e0c55d4da1429cf8dc385eb7007e95dbe0fbebb92a5392472624ac7b05efa4d93a10f0bee0ba7bfe343161c2b750958c4f1dd861127758afaeb81efec85c7cb91abc46b80a7a1600a0fbc31243167935866a974f72639ebedf611891f8223f01b749181ffbbc229887eacbe72fab6c31ea9704e9fbca9ae7bcb63832fc90b836f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h6000b9506e34d507d3ee0353629f24fc6e2a7d179f44e9d730dc08f296f326c145494f4e605a2acfe479f1b555c41fd6e88b7924a14851925ada7ea8d88fa6a42646d71814d068752392586630197abf062bbc8e32d01d0a6cc5585ba169784ae01ba8989fbde1d3af372e6b48aae66800a9c3e4263b390bf344470966e2d6dc298597c427dcde0b3b0ce72eb626d6b3d3502f4ae23ed3a52c028fa869e2273b33f8442388c0581ab2690d71460f2cb33d62c10cd0b0a31889441113c891332822d2ede2e651fbb54202a8f4721b989a2d00550f7d2f4ffcc43f1f59f7e7933d1adbdde6a61389869e2299ea4825d3d746aa2f4e8b3ab5ec749997c613eb3611decc0fb9f0e9c2f65e10214c09fe02cae4b91ecd9cab88be5e5f19e26dbc3073d34b18c78f34c9e75a4be9916c2005a3d1dc8050f0b343783c6056e2225734d0b50566a54b23484243d8d67dcee2bf81a8f3325b60024106102d46d66d0bf810accbaa779835abf84a77ea158f2632301c6205e7ca7b9078ce337645b9669e6827d4e20a44b3efcf0f6bf7051c90dd39d0332c94e2fbf6abf46abf8877fd1b024a795e10b650df24fbcb7046d330a17d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hfe16122d2f431f24667d36be31b176c984f0432106f3dc3162fb895572eab13f6abed1b2773f7e2e1e65c511d50a01877e1c95fffbda4f766f0dbf09b4f1aa0227ae92c8324db410b18bfbe99f6b99bfdbdedb338e0d559b4bdd733551576e32ae78a0f33e8f8246fb09495fe4ad8c409c40e03ae796640fe68930e5d323541d540129ff95edcf429c1cc48b0abe9fa3d19d66820fb5985cd7d0303cb2b3613503cd115e8400a7087120a307c00c968d3bc516a1496fa896151983f2718aa5bcae8478c5d70148ed63ec80e472385d2727dec094ea7cfc5aae1f98fcbd6d37d12fcae2eefaa7157d1a3ab0e60c145623da001f626bae5e0b35b63fb4ef4441a8188b1cb160186800790591ec53c63bb6b67b62b6ff96704434d9ef404f06075822c99924acc88605f01e850fddf106238b0f12735058960e347e8f0232d4a75e9d6d927f8d3387f3efc31cb699e64f2760e7bcb4b3d751dd43bede4a999292b8c1f784ccdffc1f6e811956f6f580d7ae081296f88d45b3f96020b8062bdd6875996aaf4f96804f3e30a2ca912632edce9287256371bbe1f3033455289c417ee475cfbffaf48f14953b5743ff81260220;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hc22869d4a153a325701417468f32bdcd7fdf4f1039267626f7e68cae4e8150da5db118c74d24841fc2bba52438534d8a29a2784e34d04c14f8e949ae2f01f0ca3d60a5be1062231b0fe7f4905a0c1d880d8388cfc6d534bbf700097c4b7016e199a39c0e6438be0c752ec748936fe1cd23d8432b226c3f675be3a8951f815bad79ededb96a5ca8882b736e739e475c7000407dde7c245082bc8f6994253f18efd9f64dd92ffe9abeb7fa1b36dc410ef18663530e41673416146d773bfad0f7321179f4f1613e6e1454ca2c8540170119d5413ea5b80ab424e7a74addcbb703675bc3f1cbb259afce3e46cf09ddc23078fa8da35f7eed86463165eae2cd386be6baa7a43ee64c6129246c5d52f938e7edceede55c155137fd7b06c16c7dd82d7fafaf1edbb7f1c61b682a9acc43745d6f0eca28da08da629cea4d0731bfc95258b5d673c10b4a61a92958615b74039265b6ecfa9e51db054d890bcea4fd535f26705e92d3512a5864978c73cebb5d0b3356e0f918c5d5ff4b540beda97d1bf4d9b8dba6cf80069a864acb16bc4d131c8f106c3e52c8744d9a238fa8f931a0f18250bed5a10d3b1ccc2d002ad4c77ab673;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hb33d2aca5e6807c03dd4a50e89d2251f40f78e2f30c31c677b9f3da28ac0b2cc6d61c44a12eb657d27d84fce9055118c59d2965dd0056cb7b4d6e8ce0440c17ad09418bd6967cec3cb6c707a5e39f0b71d5c4688aac4d02c7a2dcbb05a3f41e555efb0c13cbe76785d2e09d3a637963fed6029587d3fa39b63650f34adfb649fd940b775107826f4082834cb9df97eedec9a194fae5391c16e8cdc449ee6310c0ba1ded2bf030eb9c0bd3d23f026145d85f87eee40e22ad3dd4a7cac52a3eaa0e92d5279ccb2272d8ca7d2e465276d77744bb3fd1144b276d65f0bb4d9227d83827256e71ae48f0a7db1aed848f2b6711ae661e53e6d94d61f160b7a67b0c66e0a490c59c48f15a8487874a824fcae8bf43d4309e21763f592420b3d0dbc1c4812001af2cbe2a6845ba7e7b248fa4d038288f500c15b1ef5b944058a08c1f5e540eb83449a2d67d01bf50ede63e9acfdd7809cfb3c93e06c3b0c37d6921e32605d4821ce14f4b585f88fbe2b9a799c754d4c3dd656dfa0fc7b6d796eb673974c6c6522401f5c088b6e2cba65ef9b46ad540cfb28ef1b14412f7754e6e39072bbe3035dbbd63d41925253a61203460677;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h65f36e8ba931b7d79324426bfc48cdb3d86b213a6a76a16b0df205cd790ef72d6d927e7d520c57d882b87f2602cb4e562a502aba162ac45afb73aafe1da35e5de88b8c5e73a18638c87fd21f7a25c421eaaa1b4e0fccca6287663071f9a9d2e8df3ecde146c4b6f4a65d1f9081f972a451a3aa5583849d04d2809fb1cb40481188865fa489c68c42a7d8071007d34955580cc4681538cdcefd0e8044cc6590d3784f1f032ac203a25deb55df2e0c63a12a1f62b58cbcd8cd2acb547b13eea7aff62238a48baab02818fd2f8864253861661c728821abcf4cf191813e47c7c85eb6e275d6266b3d2816f92c0d38a3ea452f9a8143b88564672f21751bddc7700725ecc4a295592c6f39a22a6e4b07fca20e199da56cb6fc78bc748724ff759600af0dc172bdc011b613bdf831a600f74d46eb0b237a6b1c9fb260b42e8aff41ed93f9df34e3218ff9d4d21f3bdcb0d3d4d4a71c39ac6bcc0a464150d0ecab383196511f18fc70364ef3082e7a52a84798b6299db32046b7b172dcd251b0fe1a3c8b52ccad72337c673c007a09a45c9f366dd62e9fe06041df11422d698f979d74612ce781c958bb3d37de5bb4c87df05c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h4c8dd94afeb4c5a054aa51a32620453efe79b23ebf43dd9cf3d3b439fb9780a6144cf88430313a5d43329c0ccb0a2d6fd77b2174905fbc2d29e7651837bb7e19729182ccfb181a583344d01cb25e0b3af4dca891e1b7fb3beca86b9475a9d616827b509a799c6c5de219accaabf19f781eefe18995d1730e1a604a24f551082941b2dd32d9a5d0ea469681da63fb962482d94adb1ed0792d7240ed05d90ed99026d2ef1c6a35727e874f8c821ca93df625cdcc527369608f5b6942a8fd3aa45c8d168f7ac418ed6eb9b12a7496721affcb11bbfa4c6f30dc19e95983ed152aa6152b964897e00154eaa0b4b0b45be9df85833aca47353ac4fc8af8e0980109b195fbfd80f505bff1f455f612a096ab35325f2d2ac906e044a694809b05f18c1eee6a97f7d06aaecb6a6f64926b3cd577a44f9f6a1ac53d607e2029f463c6a0f747f5854fef5c78925c9cf0fa4cf3e4fd965f5c195179b7aad3f0d184fd671ebf76e04428f3a8bb6c99a7e55dda0738d7dc5dfc70c0527c1b42cb5c8fda1159d705785ff53c5f6e89b6f5caa884aa706056e26a5d857714dfaaf15a4b06d0d33f87e762478b36ba7a2f06ccdabd63e4e9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h8c1195ead8da01b042c5e2e7229f05f3f79067d38749989e84ed72fc8843b90a7db5c983224552d65995dfaadb24de3ae4e3ac59df063895457ff13f3e7984d9ce1dded781023183796dd6a89b2766f552ecd6977d216dfa1e8e9fb046aa7ea643e6cab1547dc8dddb3d80ba432ad59e9180a1ace07a21a5cc08a4e5ca7b159fe2c2e8424ca6fe2290628f50f12201d0d1cfc8186d0d93c95ccab4bb4707a4259dd71b688f141048401663957c17615d9b153f11370f599661666912c3fd8641515c775fdf5ad978c1a5a8542b34a1dae047cc5f12d675851ee23436e2ec78c8f1b3b0eb439baa9ffdaf8f3b80970ec8c7f48dd7537f2db789a4f572df2f0ee71ec0f202164757e68db17a0d8601128bcb7158d15f4623e0f65ab7f4d94e69ae0a6189ea0e43c123ae4b24d28f8145817bbf91ffcf010b0e50b287a3eff6b77d7e6ab267f3aa988b1c94d97b13b14b478b382f0c98c9a59769ee80a8514a386968586b89576bb1f8e9a6a35716da24cb553b1a9e7a21f9c430d70ee0821cc677b11bd4bc9aa57ec7ed448b592f031c3177ec0431072f56d3081fc720012f60ac597d605535d234d7d45716b79e4c10dc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h387623ff764c2d9f8ac67d9a009e2b6b8ed5b84d7c0dbee4e0f130d827816e9613d10cc7ba3d90fc6d6fdd256a9fad1d3c42fed6a533494bfd975a65ca84db806549fecdbf4a76d3ef0b99ad4b9ef7d39690aa95d91a49b92cf3e3ac5a1374bcdcdac8c7bcc1ca943b5d370dcb39fe40198d0953844f158dfb33197b9bf7b343cb3a53e73a24ccd10765943c9152df5fb3e60b6877c8f03e73bb7a936c46f3d83aa05060184f9934d9bed7a26760069a3233319d4f03b7f03a833a2c65f20fac0b53ff83997fa794f4f5491eff999e7cfbb049a0e07ccfd7b0c584303f054e53e541d6eea3d2a7d6b7c29f4ab86779693aef396e2a16365a3c80f557cf6e76982d83e89b78f261f473a8f991d6a7c6eb2a1fd2989c1e483aba63f58696780552d1620348213a35bd498541e304828efb5e94d16a78626a9b176d7ba3728af45d2cdb2ad50dbc0d298c7241886d8d5ae4535058038a6a7b9d035810aa28c9a48dfacc9ea10cd0e4e3293bc2023c4997b90b87648df75bf513fea7f8a84f1a1879ba7a1a045d299334cc677f729cee7b7b18122cbc01d8ffd4036d6fdec6296f3c9cf1f144fb0c6e5e608c5f0e7a23890b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'he9a6fd7ea2bd8dd03dcbfe173870f9ae017da1953574f48680beae17a851ec4b64abc2f2fe01a415abf63fa842e86c688ac07291617ae0c46e02e79547a18189a660a00ded93f03992400dc24da0b7a53519d083e77e23f76dd731e5c9351ea0bb2ab319f479803488f30a789e87eaef0a321a7725bc9a39f9e1838e615be7543ce77b2a168dd4666391daa0b0b49feb7304c1533413cb7f06f2cf228fad667de8c09188bae22c8fdad80137003734d1339775170c3b66ce440887f547f547683b4af3406a508b8c1c68061f38cd32c10d74b5ebb56b54a587921dec23f2f3ccba659f328ae006d8278376b1d140402ac1c5abf061c748ef69ab8448769831671352990640ecbfc392f885a31b26735d979b67154c5b69edf8092bfcc6bce23867315fcd42be5642636f0f7e2d78a825e311e2f63684a104cfaf829f9e1352bf984edb472ec9603eb6ec47d240306bce20e02bdc3c67639b9b888ee6c8fe77c5a45d6e4bf57d7871a743d4c0bce60306be3d22e5052302db441f02c99298cf113fe1d4b052acec6c6f2e1f42193cf5d041fc9cb33085325d961959d2669fad1d3845e0295978b7e6b5f424cb1f5c40fe;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hf6a8d66c3a278cbcf96530d5e4bced56a05889f26180bbc179133c044e7636fa6c213416ee518e1a10d042a25c5929c8dec2e9858994af0a37cac452e878cf687fb648b3d1ad8d0382b75eb9ed572fcb5bec7ae0cfb11f857813f347441b6c921130e86c159898705046429a73baf689b6f27408c3bcee9e3754fdfd15f697d7682d0dd3e584f4271b6986a470809220b083ae76ddcb15a1e019e7d6578bf9ce9a9fe68eee213143163a1d728edd9c2b496e71afe70a397075f9be688b6c6fe117c6f6b3316f95ba5678cac096e04fcf0b446fd191f6bb0a31b84c5e0b7ff7f34afd18e57dda8916e6490aea3284e73cf14530f584abf8e42867afbd87c6243fd83b88a2ab47816c017dde6d14d6d6c563a71a3c7f5470e595f2bda915e408c407a9253a810ac1e5868830540216ed3bd513e908921bdabe2853a06ec4b9589bf5e0b9c7805848fbb869466e4137a8869c04a8c37a6892bba4b7004f45014657bd3d4fe980a6253ce176e17b93ff5f836aaa88b864cf1a316351d8b68c2e56f14320abdc8810e973fdd53a95c2f912f62d3a1652e00dca71b718b01a9cbd01b853d4deff5b9dd6960244a5fae62c7684;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h6c2b2b3e5e825222b2c139c44912cdfead777e0f30b088ed5e318a0883f0342a2ddd3254982c066269fb2d07fb946ca071a68a880120039dc8d044dce1451178f5f98d46c8c289e9c678665d6560f8062283d4d5959fe940848411a489f762d2c70882e70a6da171e5944c79f323824299d9b8b78fbfb7eb660cc5bf2ef42cd4ea10ee7c39140d548690bc6e569e5ebdce56c33de12954f85cdd1995f014df32f78d01c75ca9edfcab5c328710ee2b4ffa7ea83c5f74ec6ea225a6dd4084225f5c3c65956aa21aa30e0d999342d71e0538976eb9adba871b0999cb2d3c1f3b7c662ee6aa83949af4acd2bb07f0d3f4ff6688ec8577ba557e35349e16c868a8c68d00155668b8ee87c0c395ba09ba280cc9e3b9602a5aa70a99a6fb5939ee6ac705a58cf666e4ea71dc346962bd18c6af935af7a7f9aa026ca44182e930a9b516326daad447db6fd1e9ba8ca746c710c0f71be4263cbac57d2b97f9b5fca9a2a1d5ef7dc7a17b123b24a0d985fba83b034981bd57eb9daf70368343e9feb641467f392faaaeb48354ba62b14ff9baa2da2a6a47f7eb4fd2d6f7d4461bf9fb0fb2adf7c3c74bc7a0ad2955058ddee5bf5a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hb307dab6aee7c4c7cdaa459c45457f3401b52080707769c676f5fee466a92724e296f91ca20a49102bd258826bc9537bbab58f024d4cec8cd0a320b2fc994056140d3470a5548937bd9b61035cd9c7b2d05ac5ac5a5128cdb239f989d9644808fca0a11104697083a06579d73c669ab9c37ec08781495c48d8d056e08f03291d3870b93b63fa4664d7d013b1fd63014d1f4c43166fd11669cb380c4d2a2448d625e0efe91f05a1c0ad17a64458d38ee2e91e146ae4f52178d2a1667827e866c71e0517b8ffc98eb39d667ca1ba3133fb37fb7934401d64867df6a1bb0d6aa406a2df00c696e3c01b9b4a4953e8e31cb5c9b6468d3ad8705b310bf19e5c91cd103371e27b03987f7ac0333a76bb2358fdc217b8c3c945f11d6350a8e595c74d90eae39e5abd94fd21817239e13c77af56c929b823f3e14022af926c1cea11c3973f66727a9a4a618b8f604f49852827f68ce60a9bf2c39f146bef4cfbebb798195c3131cc689d112ee75ab2beef981384f09bcad9b0c0c5e7eab9d800ce79425bf2cb856385f0de4f9dc594947a31591d40e87849e606003baaca5b1fd4f4ffeffd477261508326626c3f13f3041145f9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'haf2cd672a331883542926f681cd275b1c0926673b02255121d8018a8f2660ac89423dbc0af242557ae8cde3a55b8a2216ec01c110f8ea0bc3bb4232bd2855842e40a3990536736f042ef54029fcf2de903a512822f3894046da6123911a8fb1b84ec6381df40c3f1910591d13cf72a53a70792908e944e87f3af743855a54bf7b365a370e70d4d54d4344afd4f710a774a8009ecea50fb475df7da8a474a6a9cfe4dc9a65ec3d68b427227c4b055557294e05fbd21e200dc618327ad6ff25fbdfcda9f9171f0e556a08c27be517769e07b9c2e42c68c96c12436f538217aae8f9ce7a83a66558c0d949b3eda6a563e90dff74ec8575d2518d6d955163137bfd68e01f122c1b241cbd42a58e160adf58bb1084eedebea536c0cf4fab52f06202f6130bb2ca4584171a23b6f15d57bb97b3449824e7720e583558782de58aba4244df493c644f7aa24ddc57581c53db271da207156615b15544c93d12eb4b2296b77a892c539ecbe63660c4047f89281d6cea21daad8dc55e54f07732e225376f05c9d80a962a5cf6b5875e7bcffbc7fa6ccafa08313bc01010138b715cdd36525c50524c1ea57a0dfad81575809725267;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hf457637da5bc59ef0fb70806ab4de6f00e48d9c5bd32ffed4db9dffed4cbcb68f6b86067f77144c46d0284d1c42e841f8acc87a683ef560d51feeab4818f25c46342281857b2afaef874c93ff936245ad122e25f09be5b68dd6f713202e8475c8e3bb8de07adfa9627660ea5f8acbc530db0316631def7ef366aec271f7874552e333a85f4e5b2cb5e948c2e68e61f7464ad534e4aa2efbaaa6d7a4dcc2e022a0d584f2adc078b052665d9c552a83350fea01f8388be9f9dfc45b1d07b9837c21604e98e7e91de4dc3b1e607c750964ee0fc8901ec68dfc4f4049bebc05b3b2aa6feff568ae4574d5c609ee843f1479acf3b3b807bf6189bf4a53e3c2a702d4b38956ce0bc6008c0d8792211b682f79d0813e407ff1102a495e9157b703423f57359932444c065897bd052f2cc868c5b63278a744e4d42f009b0a427c6d4dff1a683d72598e5b110b4d27b475ce2a1c021a28ac5941753ce6a3d18fe3b7ea0de080c84785950c168da8a8596375aa3bfdc7d0eed22bb9127804847e7f38a6f59afcf6ba56586a3d83b9192e1652c95cb05a0ea096ddf680b9dd7560efbc146eb89bebc3b6945c1215e0b45c8e858a46b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h17ea3e0453643f4e34252285f7e0d1598448548e6a21d38ee2b29a999833f0c2299d3a9e21e4d1d3faa0ff97fec2b857e1204f9401f06ca5a1726da29939ab4b5c2a40a8e8a89da67afad7c896dbb0d6f3fd5660af40e244bbd02831bfba812566493b56d1ff3dc54a6bb580e370336521a9b8b857ef95604e1db31ca789d14e12c000f3937079bb9e6f9dc8d6d75ef7b73c0bfaab460db0abda14f266a8008440d40cea77ae0b3e40767aa83b32857a124587426df77a6f0ec139f802c34a17f6127256770be712ee86d20e9dc58bf6a8c82011edf0658ab21e6f3263e7165278962e0e6aca6a362562f6138944e1c03596d3d82261a4e71bd3d33a61b5d5c41063b3a922f859267a26979a8e27ffa8e15f18c5fab06e4899ff73d27e76cbc766ee4488c88337d93c5c3757567f1048e0da1517a7d2609bca33ca758876e2aa48f31e6b55c513e90ef1880f7804a4186f205e6c8ed804e46661b2f2d4e3ec2ee990d13fd8b910e3124a0a8023e647684280a30328ac3a20536dca0f9399c8b91d580bff9a8b809f9a392083be5e57c8ddb7bd18a446dd795f34064547d01f798e92e2d59b8ae984d20a9eda06e7166e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'heed9a9e2948f872c6927c91a61c6051cd8c5669ba334f76bee522e7ce31479aa275e16e6fc57ef9f3b5e8575fab2f670dde2cf702b311f08cc79a30047206a5b81ec333f5a36a415e8700ec347f70743f3003b34144230d431fe513b73f5203ec012f12f08f2714f2f876eb4ef69d6e87c9763a1a919bbbed1800265f1678d71f487029c026e3b800b6aa9173bbff8328e1e0e952a67bdfbb49b4c5c993155106a9936a1d3a40d7e79241cc04cdbe7115131c56e1f27281f53c5e31906047c1fd82d70f8f3a2f5703ba08a1d2bf56b1d4a513f0ca586afadbebdadbaaca44c07c73534274f0c7f284fd7991d5355a269fa8720e029865932baf0ab6e098e365b61b252fbb6f19ca0357bb966187ff0b948a8f2dd80d2d23bbd403df85c0ecfa93467fea99d427ff06888701ed2bcdd8e59b2541c760bf9993ceb8708d15c2bf706104db793424f626603d55d6d91e8121587b32b657401b5f0e7ab5f848fd8d5d6162585e799ce8aa7f52a1804cc11fd14577169ea59b7d7129faa7d5d6e6408db74646548ef1b4ae8303de9a01cd3ee6567a6a59083c63a945d66ece150dd45edb89648dec019bba32bb0e4ba306aec;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h9d1bcd5b1e0cabac74522baac085131a454d55967ee9ba776b849c13f2b4ce67a9db2f98f0a7fbaefa45634e9678490a7f4d18a27e84e16a03e898051c74cd28d8a467845035aa6a5c5b44a4d82e7b3137f3f953fc46b11799198b18f736059979a1060c3e45a22f2d02117305229726938c43e90d3f7ae234f3d83ec7ccfd176e4cdec7dcbd77502080808c0ed5faceeb2d62eaf1f8c66cc1c0dac63c664988758a84d7ceb9e7bc2dc5de1b5993f3f45c2b1a354eb36f811d2318b6937674e402d9c82ade592f3f0087b11d32a17d4353a6096d3bf804b7bfb21aff032b9756f154a6899e67c6bafca0a95e7b858d8555a4ebdd2389e12432d30eee2ffe06e35473565fc5ba7f995ede1fa37673ce971bba0ae59dd4ec1fe90905951bd6b3e603ff801370318881682a99788f0544566d534c736c36f3954e66eada47d48f57bc7ee626d591f9c10aa768a85d95056dc64fec1a52f591df1ad3f1c843112311721dbdd146dda8c2be653312effe407b381941c34d542b1eb1d521c03ce5497bf73001e54887cff8860aaccf12ca5032271e9b806bc01bd75e1c550147b8818a9777cd81ed702da7456f3a8c23302aff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h2147edae94271679bb8b809c313c530b8d07bf9cfd4dd6012806ef09485b93329f6c1876e7fea42b455906858c75a6cfc8a90467d2bb0a62eaf5176f228b240505d47d25b22c8a3125e7ea5fc4f066afdd8bd195b7ffc75c930b6d9058839ee021538ec2aca986e1bacd11df00bfc647f9531d53209a623e7975144cd4a862669cce881e605ab46372d5db01bb61205b81e4364277193d93e178643318c8af17fe9fc633e25b303d3b81bc75386ace072a05f08d743b96a535ee1981f3290b9fc377370d6d399aca8a5799622f2b6e6557ed23275886546603ba77ed7c042bf559e5d486ca2d7b866c0ab871bc0cfdf7270925fc0186868d3713094340ae75e2ebd3a1544ca01f9630329ee301049cb66c75fac5bf2cec3d75599d3ed5542a0c5f7d97fc5ad8d6e998ea85a492438dad36f3f2349d3a08d146ba5577010cccfa482cc1d58115b8cf2d2b80b4b8bbd7f60609b024726553d9d023b9b2d9d65daa95d5656d8a24df98f607c5eb30df7745dee7d3989e34ca2e7720624d9aad7fd257214af8a1a77fecfc0219e0bdff6689d3b52baf0658abd0b0643b27487fb6ca3499e1dfd533b30ca8e99e80f0fb993d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h3b47a0cc5236a29c9d4cf0bf708f7de42b19a46fde0c93fffc67777d8ff242edb95a47828ae7fdebf4ea307439fe1a0a8c37ee71e7487beda9a3af475003ae19e55808f8967fdcefdd35195ce50b302e277e973b262298504e59b555b43558908bb85910e112298a99fd3c21d078e0633999d97b955a3b73357422ba601f34848d64a7404ae431157d7984de65224bb9f44731761a58b07bae31741b06334d2c0176c9e8f62554a3dd9689f4f884b802ad36032812ee6ed76c842b7f433e1c0b6bb51c412a22a5c530dfd8aa75255372fdb10229598dd352187699ed2166eb78b02c5fe83c904574e7e5a36ee3ad0d404870c8b21243efca461971c356c7a7bc2e551d22cb748d0fc4b4b39b0747bde58a05a1e90200e7c1ec5435e9917bf6c8b1ebfef5322b5e91f5db07259eb6ba44754db971cfb949b6d18bab24e6facb817ade6eaadc62c3cda9578652c7b886b39a5cd96e0f6f62f48efcea68bd3cf6faa143eccb08c65550dfe393b944d5342550182b972834d3ec2aefe1020b55a8580b2058ff1a8a0d3cf489d941e9854de6653f4f20d056a0c5607f60a848e098458528af5ce918e9c05617020f1074eeeb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h9583c61ce40091a5be21370fa619d6c9f6e6d18863a8d71d5f7d155edb31ec57ce8201d025ce7424160292325e26f8f252027c81d1481bbb12bacee40036cad6cca7f1b0e7ec931b265551e48b742052a6e466db3357a57ec061d13d2a8fa1e47d00fb582f81b4e1539416dca194b99b5f9f3c9434fdcee017ed7ee95d056a4939693405dae8295978101dcea07b52a08506e770d0fbe0bc8ca1a73d7f21d9366b5e353b4b728e0ebec5fd0f2bd5d692076a1f54b9628929daccb60198a9685eb18c45f2fca74c6ec2c830ffb40e6c733ed760e021765849d924e4f47fd2b97bc868cb82aea3d1e9b28d9f75e512d70664d48c526287474381e1f221b7c5d50b35272b56a8e99bed5149cf63fb817880f2d2d41246ba946188c2c1cd13f42674f621796db944a70ec4236dbb25b4f8e5cd76b22828ab56c95ff1973750cf77a8942bb374602f18531989438de923a7b06d49e9a84b489d2bc25a1965e0783c905cd913482f7f1c12a299d182539bacea696322227be90e4097dfb34ca4692633bcef4dcf28c30e339fedfd20e51ad7fac938ecb75dfaa5d44693a1adbc2186b5444020a74cbe0674132119e33b2394d6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hef0921838da0ef2eac16628d423cd83a4de878aa7ec4f79a2add1c27a931b8a44dd32adb4c6348bd0f31d59b1f6d004299e946c37d9139b1f4d2a6148a9c6b4d07864591492e48c615fa8ae19d31b81968bcf1df8eddf6c3e86fc33a6e84b0ebe55afd4acb99f7f31dfccc7a873d810e334fc7e2affd37a83d531531c5fecc3ede1410fdf415c4367a80b47a5ecaf857b2033d3b761f5d39a12009d0e6d226bebe64a15cb6f3ebbd20b3a2ac86e4fb4f06e77760cb9c24e0d454b633d4777909a20bfd71132a24e52be2bd88e8de91ec19de57cb36dcfdd8c64869449aa706a6bfd308028c4ebf5dff6abd839d40116d5cd854476f651dc75ae45f56262061ec3fbd3d6ccef49fc085d492119cb68df5f796015ec5440c5f6c7deaa56be0e564aa1e70f937d1add215bf79461558156080c817808c9c4be7e61d209c206b2dfd5a70b9127bf62b7e34f7041d9ab3cedc2a7c38560f3d38f5e144d30d944c851f8153614e76aa86bc0c631c4962fd82c02c06ab73d1eae0d57bb6650349f45290b3e1fa5925d70f8e9f1ff0a852220816333a69ec2aa09d66dc53b93bfe19dc7115227e786d109a8f394f64468b12a7c0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h614352b21dec01b6a093c06c78550e04493c163baa17837c616104c224b32d2fc8bbf8d3c594ee1cb6c996c223c6bf53985284a8c695f660025754e2ff324d20ec5c281d31a8392765741c8c9bfab1d085d05982a13a41676fb0d23e72852e8f1bc6e0cc6c8f23e2fc8d0d2bf435a8d2a6fa9344a5572165c4dac248c1346482f73f0343ce712f04ecb7efa53656d3473feb5e573f5d261daaf65b13ceb7e90f82bcee7907ecdcc67aaaec226acbca1fb4a24e0ff4d6ec7fe209c4bba686dbeb0ab97e0c3974f79c7b72ed3f668668fb4d20613e251f61cf41857acf5e378cd36bc80fc772beb9878fa59b2883c63c170dafef1b89a27c8cda8c346bfdcc197ab1f5a73f682dfe638699ba83aef57267862c34dd8a8a3b85efeab2820f996b2d10b3f464a764ff6ebef4ea41896e46ff282bfc29d600ba3f9f35feaa5e9bd13a41bd79f67572ba477081a518e86ac132bd540e569bb4bab9e1b956ad68873b07a18609149cf6387212059e025ad0a3b696735be30d99844a5834d9818c08c40fecd757bce2b3f19d2a6916cf738013823438bbbe79b11a3b6374fdbd36382d6d1dd2460f32c2401f1f2906ab3573078e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h7d19ce527bec41d6fa011478d6ac2d2a87470da77c3780da135de5d78ab76209d4be8a643f2705e2aa2dc3271bb9012497c40874641cd613e489ee235fe74904fdcf739712140729a21bc2fb8029e7e735f96ede24928a8aa95d18fb8fe1eb2b11fa8dd8b3ea0ca651ae2856cbbaba491eac15062979ad921cc1ec5b6b2d1a6291c0685ae358b400d791c3ed494c17ef949a66abaff6284cc9174791ac58a160d1014e13862fcf4dc442c52bc38cd2c78258d66b41a9e680ea64a37de5651a37eb573589ab35a84452af2389fb070f7254e4b82ab3bad0d2176db075279bca89a2241250ab8c085bf69df8ca7aa90881bfa5e9f4afe09d5cc48df2e80729a2cf65a2fd0ea49061ce38345a4858bee517ad6d5778b58428fd3706083684c92f0029dfe6f3d79f560842e82ad1a68d4a94bfad69408b6ec7310201f27a83465e04bcc1ec0dd0955096861ddc9b2b6f05a02c57a5106ca27e921a97f3c7f49c052ca005999e7796bf9064fa5b50012271f80b70999afbe4bee6faa59be32667cbe1a5b5f44c8445c5cd0af193500ba913a018a409c30b4dbd9e69b34cfc650bdd591f51ce069b5a3be61a69acf8cc0f3ce3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h63001707c421f8e0d841e7652b5fb37e01a1344bea865f5c38079501f66d6ac314d74ea09156edef4b9f9ffcf4705153b07acf6bf2a4064a6996520bad720627c256021d091f04e7866825475a1da6ebb9d17015e0c389057d30b99034ed30c43136ad968b1998187b969b0b628ef00a863cc46baaf642af25879bf843c87782b7da306c52c3927883291654ca95767c8d2953a3e801f9cbe5d8d8192f05a2a8743653cac275cf423f7c71ca67e77a19c70731bbb9f3bf3013e897d5b03b501f46f5f7a7d99e13974d76af6e13fd6aad1b6fa8b1427aa77f6f563e73395367104bea0a6b28ba2dab47e087da8311262afaf41b8f5018edadca94e48ca8b7f585b4effffd546fb9288027cc7cbf2ef30f575a07d2c79176be29b24b0d0c043c9f79b940211f440b264ed9b038233a38175e928955544f7fb7ed3938a4192c3a409f5366579026323d07031744972f44cde6af507ee13e0d49dec0507dc6b682ed2ddb7086444c65c564df967a0db765bec806204994f9812df103aabed3cfd1196756350902a9e5b1c1dfbcc447628a657504425f233103574503d5db5813dc48c753f08364fc67bcd82f29f6173c0c34;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'he2af6462dbc0a8ec070f4849f13fe8771a5d79a1f711403ece886e98bd3493a640266441d9eaebb491d42caaf2eec9f4c51498b8d0af5dbf83844aa852db3ffbc2088c9af82c7c6a4d5f4dfac6cb5c8e9a4220a1899a3a877b5fdbb67fc060c8bede56860c5d3d3869b802ca82bb7fd0f512d3368e08a64dcbcb79d9cea8c00d274954e7ccdd09e6ba71f12f2e4a9f49f76c250b45b22d0b072459e50cf730308a1ce3e52814bd94c2f84c29b238ebb16a972b6ea09d08119577106cd5bd13c6f309e208a9d2be59a4be952ba8a406e304d49a6dae9ebc17c4003ec4f9605ed93b19f076926d19656bb00608d6cc7b26b0a705d1d41f155df4ced90472bf0d5c1f289b64a1c7ea1279c4001a707746f1533a26fc7c0abd6dd887452f0c6a14bb0ff7d6898ec0c074348de997cfff204fff3ef543b91494d26a120ace900ae9cb7e9787ed791543f9d81651fbb04c7b858df6c69937d757a9e8d2bb50584ad4b599659ce5e7dec02812d7a95671641ebf7c59474b1702bc6ce28f0a9405ed59ad282ecabfd573ff5acaf95a29e380112b74aa8d7203a1bdf944a2d6c734b26e3e45d9749afd93905f8cefcea7d4653d88;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hdcd1ee87ee2a612a780dab216b05ce25e2b52fea6e93b2cad2e8dcb5508f261c47e53073dcfcad47c884bead92e9c12aed8a2de41751a987e011e3412243e9727adfa358c3a5a3b015d244be100bd6a294e24021dd13c1f895498b9ae7458e32ed5a4f2a533990cd7af182d17a4e02b6d9dbc90e50b232cbaeb1e621bbaeb03b01c6b31a999e2e828193eeb1d0502d0f379d7472de7b6fe429cbe51506e15c69ee0130429ded673b6a5ed33dfc6117ff7bc70ac7878b342c427cda53668dae01dfded69dfaf96579983260ebd81dccc2463def24d100ed0beea557b07f620ac53148766f70081af60bbf79c0d8fe814389cae4a8f53db6ce3d34d4343380b515e34691a2e18ada0e9ef7608256a23d6b3f3148009b310606af400233697b638426bec833debba3c790cd7bfa738eeb60f8f6c4cbb50d08880524d4f5d7686cb1191f90afbff67672769928a8f7679a2d9e69bbccb3efc896b373f9b32a4fa3c62f50d119db80fbcffb80206d8b7bdf9c39fdbed7cca539b1c37ba029ba9573d4436112ebb56fa504813250369dd5a4ed81964af1c97ae30ae3609841f0be6da27bd1990549f9687de511b91602075141;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hdbc19057d5ec75445ed16242a65b25ebf4ec80f257b65489c2e126bd3503d1aabf0599b5b58c107011f9c4322d21b2b4155a6288944fe71c2ab63386ba05f714ef42dd3dca63f3194394c71c192b889cc4690de00efdf792dd2fb08d1b95fc4f52ec1955021c2833e2f910627be1541e8468b250a6e34ee6cd5f334c06a56d410c7627136bc6cf1ab7db338039f3b40c98d64961897672a5add851c4fca4ce86b59b149e9ca306fa609f12c1a315e41f163865fdb8f37f71c924e0f623c2bc7b17c98593a81afe9cffc1cbd39673d5b44f10ce806e594ff7ee19dadcc8995692932036ccd8841b143efecd894a4d20b70baf02624e1a38b4eddca4c2c54dcab2cca4764fbafac407cd6c4f35d6c29fba31d42e3311a30e811d499220435101753cc1946ff5db0c55c8bb1daaa7507f472ad446554b6c7304662ec652d7495dc0664c2148d0404ae2330bda3d12c2bbeda8ff35c4476090b8115e11bf128d1872e01e1a14f7091bea231b579143c293afdc40f85308bc74e5e7803f79a1f12623a1b99ba0716b3fed008e3d2ee7b055678dc6d71602f647ae40491cc7813b32c6f8670f52dc80af8aabd62c5277acf1a7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h22f1bce9cb1217510b94e78346039ba9d23d76804d0b8a6d516d3b43207c0e3356280805eeac5ccf4b41413a857a449096e3f8bc1434ae53224870e0588e0d05ac4fb7db772139bad087206468ed09f7626b03c26822a2f27c21096a3e1f6b437e0e6d63508115f361d9dd1e927ae9f143404b97f9f3e22133668f081b3869815728beec2cbc9956cfefee1e1afd644f1f329da7d4f020c10d68e220bf4d40b21ea6202df69439a58d9f06d1b2df83f47e1a62cc7cb566747b285b536fd3c98aef11c10d5fb14a6c36747603c9f4eb4e17d21581f331312cf76d3f8febf04d459104d56d5be7415690ce64a7280c92888dc2d058a41d7d763710093b3a27f48d33863607d7e7b019b8c044ec865e4d3f34f0e8b0fd3602542b96a1cbaa198550c89138df9b9ba05357117c8d0d3292cf4629464fcde84acbb17cf46cc2242d5a1eed7f702ec1dba37d5699f37aec7a98b2ce8fa842bb3bd7a82952e662b9d54cf2592399309c5a2a8db83ccefe12f74f914fa629f7ea9f5de48fa425e8c1dd9cb0ca4db43da50171577d575ee518d277153fabec2901f85160505430a9f440c13c5a11323127aaf01ff11f5cf8a70fb6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hbab824ba4b6ec07cdbc6417dfb79bc821f2a97c9f3c22a5d3ca5982e797fcacfaf0e6eb306483fb6e3dcaf4a190d558dd8222666f4d0fd23800ecf499eb26cad0d56f63a9cf42887c975388a560f2b2ae1e46709b15230679be07095482d7475ec9fcd9be6d8742d0b9b891b20cb50e32d5ede8f5d35ab136cf6e52de666e5fd5d3ad40fb264eac8d0c6899ae7babc1902f12ae42ee34b68caf2b3cab95082725a66397f0d68d941ff2ae136f47493936d122ba720498ff219e4d043881369f23ddabf1901a92f0abc554077d628144cf214f1a3bef2e8274e8ad682a7898b9572ac22f2de8008124974c97b365f64bb151f8f63ccb7e7af0d8c08c53cecd94e172fc9599939d8b6e5d461750be3ac9160f7a570c99adcf788fed2ad5cd64c5c22c43ce6461ba17b23aa906714cf037e325dcbb2f46d215f9a62e5618e8a471e5c2b2355e0fa67f360746064dec0acc3c07b5266c5a9647c5763862a446eaac6d5563e2693c35d3275cc523504b41774fd5be71c7e4087aa5e286cd7cd1a14a4ed89eb4b083ce34f2aed28d212f67a402e25822130d6bbd37922d414a6a9d83fdc032ff9e9f33abe3f30ab98ab176053;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h2e67e082db616d160d0c5029036156f1c64053b9f7a92487e26c2c6a1f4d6ff7002dbeba6b264fb57155c29e61dec4af32d8ca8f7afd9159c7a0f07f459cfc90786f006bcdba1373c9a4117252fdcd55636b4013843f3e804ff2bfd89d73d8d0deeaf2853a76354c4fa867fa38c49f999286f395d4d4917926c76e8d8d61291ce77b1abd07c6173dae9e86abe8e74998bd3aa7655827f64af31480735e8abc24c33b396776fe076dab612b161217b10c0a1e5eaa80cd69060b6793cd6916d8161c56c28d0cdab19327f12f46afdce258985a7b7fbbe50f2fec57cde3d3e32dd7e48c82710d7b2600ee9c46215018a9adb791dbdba5afb110db06387e1f60866537ba58e1e94e6307e5ac0d8407703c6c6963f0be08286287d08811b8055df334c8d8b7e368301cc0ebe70b4862a9fa7e99b878b42360209eaebe0194ca4e4f4e956bed0326d03fd6fa8ff0ff74aa3aee703afef6e4f44bf512e271fd1dc817ac172031254b225e8123e943cbc4669045755ae2e0388d77d19f0ac33ff242521ce3804203370e571d5a83a114ed0412e62240059791a4f80a44c637abe10ebe827af1791feef02fe41106987efab2ccbe;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h25af364b0f9bff34a7334cc6c0051fbde59ed123d096d48afd4489f0d4e624d2e2b41193219daa3cde72928ccf9db76bf6ea616f8bce7be07c030657f394b6e40648d38e53f4158314f87ce74a14ac64aa3200004c0dba39b55a53f2ae6875221fd857fd01d36dd6b6a7d0bdc99064c0826a5e7b1944300d48021563988e2f071df6cd44006d38c4467aae6e62472de88c4c5a60fe93d1896d33cea69eba6f3ed7348709c58dc02838f03bf36571074e28a507a1b703677a824475d487dc8d5ebe395481c6e9428fdd75d65071829770c5f4450b7f1b487b8c6ba9b7e7e0cc82e922ee8a4b090ea1230d696aee30a35ada98714605e0b07139136f8e94c16b9ad3ac794d85c3e4cf7011febdf7bb452609c2374dc8d75b66da9d27106abb84af7deeccaeef14561dc8cb6d387a1e32a54081e3148b2e7a91db3fededf94063ff958678806df21d76bb0f59f7e2e8b126aa177ff07d6415b9c773629ca12dc915235895806d6f509cd160fcf6a51b8fd31d004375a09810ca9bf870476f2ffbf268eefc5ae6b2e751d0c8f1ee0fcf75ab47d0ff7f11223edbd29d6ae87397c055bc47a4273fbfd13beb82062c0580c4cf;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h5edd57e70d6a3b5f7e720602b129dc9425b41074b4dbf8a4785c25d9c79c76af63fede646fc44e1c9cedd42116acc97fc874a005091232b4e10daa5664e13456e5445f60fda4393c4b4cf2dfe7e9ff43353c8ce8f55309573ba8a7818d7cc80ac77f1f67e8396cabce8e14c9969219042e9814a328152c87d7cbeb925715740cdd5a2d14ed487c84da88da56fcd965e0c2b448c646ebc5d6a2b5ffd8fe39cf795fff4afac5bff7f2556756654f21ca2efbbe55c502ab54852f3f27241621309127afb7567d56b823ff38c04386ec41b7ce2b8eed6cc202d1adc4b798f9a48b002c8b35c369666b164f5f11b6fe361369ddd5cc9200cf049364cb7580723ff89b15751a59a5fee4237c366217cc44e93b879048052f963079527af7bac5e95888df40b5a03c4cc25245db307f7a44a883dba229dc4714bf5e790c9ec18a5ff772bab5ba98827c03041ec506613d5454baa500b5784da838685a5031a2febc9a38b06df9225e76ae650cced98239df1e6c76c893327286e466054ef9eb7e4705f77eb34ccbc416cf426fd67937445e96a2f66ba4fb902884119e45c226003a0059531e39bdab5f523769ba1ea968e98103;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h6f3f3057fae988a6fab603b04d5ecee170ac507e1bf814d5132e2d9a01f2edc24062943f41b76d13a544cfef8eeb55b1fd33c16a6d4556c71a628e2f4eb030e1075460f467e48cf7c5ecae47c9f3084964022304cd9c2e7768ee9366ef7b98ae12073fc960a728d31393c22ef4b24264fbb5addb93ba486d159ae97a837a30d64d841d59714d72b8358a015d4343e887f499e628869e5835cb931acb66eb5af76f0fde8759e07ae60f0c03b24034427cf349dbf614bf8bd11a2c0853f4900d6b942186d557ecf1a4349b1bc9a12dc8684d0478efef2a4b4e9d08de10556a9586dcd1c63a4d15a9a4882dcdd48c38fcd67f0127bbdcf23e02f590c65fd1918726ffced10141fbd07fbbab92187499f4e09baafe305d4a00edf027e1b4fa650d4d79a4e8f3f474f1952b4ac846d8f19e7980b8a96857b561da48b90266ee517502347b179b27b819b2cfc05c9818f798fc182ec1ed7687d53216c55cc0020ce6bc85c89326e307aa6a1355a479d409fcb0924c2c5db0c0dfa98869b60403a93025591a7538d3fbf42d9cf3fb0cda61946926ef5ccb1541f84e8e95d57b4adc0b8a311057b1b464178e770eedd559e1e5aa;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h650bd08ba511197dab5d1a44075bc43939f0e3c9d2675ec5f6cd99981eb47f66d39e51369497122474c9f1d5efca664c5c64d4a0b3bad91ad8feaded4914e60106edd427fd7de7fe2aaf39fd5f3bf416919a558ae5bc2d1cd66b1e60b3edb11b4ac49c1282de93b34d7cdf2513974b50286a2b8bee5de499627c956bf5ccbcca75b021368ac3c5be535b5432dd42c21d8e1cb20afb33ac24ba7952d50a200714ea635993a5f44af03d624db6f579373e5220d6be9a711aa737872f21b53596951058a3b18c1cb48c3466b52a7237665ecf32e7e7e29d45d8be51e42fc64d11f7ccb27746e78472285edd21621e67e9bb68c071f52970088592854644642722c2bcac6611bda82f550ef496eb88ed95175f9c4aeaaa6895f2a14e50cf167c282d4a4296c12e2618de2083061f12e8e6d075407f942bf9cd7756d0736cd61a7b98b5e1081a0667fffa04c9334805168086bbf18b7ca7d7d58595fab97c661f998fc3f194f50515ecf3e010b2208827907b14c84ccc4411c686ebd23ec30bc30cd574fda20a31f03097a7021e870b185db3feb339ce9f2e6b88bfd2bfd843ec23dc10c5692b8f1ba6a7828bffc8eccb62e2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hafa9346ab3b8f3b3ddb1b06dacfd50dd95a2c06f2babd0f64c719511d37db087cf8e7ca1c49eb05fc23c8e7fb6fc0ebcfa6e5beca1eec35cc45fe3676b4bd8cdc8e3023ef33351bd8f011d7e4e4c3910ff4e7802051291d365f9db828e320753bacdb7a7cef8e1d21163abdb3ad98ee6cda76ea6f0aa7d4bd2586714b28e2ec940459b975c3be9e6943f37c921eca281f6d08fc6104d9ffdecebf3464bec0798bd501e20eefbebc9f56e14e205bb4d00ca37bec3b77ddf67c67edecc771446f72cd4a3df8fd5b16f8410f573c71f53110d09bb5a2f2345587829f062aa320da38b8d80ce8973fc3f1e1e86fbe9c309bfdd85ee8141119fe8ddcefa65fd2da6bb20e74d058ac867f74d7cbc9781504665bda2ce9e023025e7a95381f1040a3eeba0253064f47836b34bcd0643016b0d864fd4b91be918fdb8ba84852c7736be9370c42af5890043ab7fdf49ca102eea86dbdab5c470324e0f29b6f3f58b85cfad23827d6c9935a87a62b868a9200aaa53daf9d0ad68c6c58d2746cdfc687cb987705baad97fd16fdacf9b0fa374cdf63985437206c1fa6bb911bb2443044554d67e379071828dc24c89f781ecf13b4623;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hf12be42b759cdf79fdb3e6a6e842989626154fde90bbbc28d258711f5689c9e2f9cba556f73005bdb08bf1cb59ee6e608bea8c72349e2702394a5b1fe8ac4867b9500941ef2546acd9f8aa326de5574f3c675366460bb8ee50578436bc699c25dd2111cccd8d2da59512d7da6f40b6bc7e1b6ab6d052fac18eb924c8158b893a5d6dd497ce722b36730f87fd49ba9cb5cd347cfe5b894e8cf873d879c494fde07f475e084ca8ef3c236123afb8c7534e63806042bf8bec18d18ab52cf7155dba327b31c3d68cff445ae705565618637b4d839e38b353d360fe30ebe860a8719ad2530af984dc05b3b092f00614a74e3e069f2cb79ec677d8a958c69880557d5edc220dba908eae485baa5defcfa57c01103c15cff32795b68780f19516fe1402d9bea05190de161e51776e3d435c4f1ada68858872cf9a8c4a6af478d2fd25af0ed60e879da968054458463d4f3f32f6f766a00ef466156a1f0b2e58ed88cd21f1e4d36b4765c76112a7181bf4256a4b11e9505c4573bce02cdd12521c66c5c04882515c31e1f0c076df30954d985b0e96a658eeb8260c33a81cd3641e32f5412ba1f4fa833cfdcbc10f6da602ffaec6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hcb7c0dc231ce265c0bc16593b6ac919b9d215d99c60974ee9944e6dd280dcf2ef0320fe8ec5f675f5525ab3b12a2c38c0bbf32d8d7a06072f2f503b4e3fe4073a8b91b3379f797f89796ef1aa2895b275f9d6618323a5912a01a3fefcc30e621fea5b35c2da0e005ae8e5775d89e162d1ea13dba8b27c90d5bbcef933166bc4c106ef34a77a54d5094388e6347d97a3e2527eb66bc8bce84b1bc820684bb77a0ff1fc3565408583298a5cb11147eab9d0d09eaf476c6804edc76eb027af97803fbd8c43ca743f76cd55e1b53c58ad539e499f68e1e070fe87fd31a4e4c34315288b6d9f2213c45e679f1eb790a83977bcf977952ab655cebfc5cf3e7c0e578523d0292dcc96d63e45d85540eeec0f1ec1f66d9afa57072690a09c37442e0ae2811a98d83725da28dceb6d2a5d864c41565e6cbf50f23193eaa0e206e08f96982ecfeaa689303aac5074c5b099c082f7304d86081abb8ceeb7f46a866330423f3b9fec2beed016104e1826be42b70d766e2985383a8b2c21254926ec838176ea76569041e0904bd5d9ff00ce60e901cdeda7eba4992ab8d2081be4b84a2fcd9d9c405470bea83a4f64bada4cdc2dd7485;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h32899125cc53894929f9e7386c4f4311eccae8f68be6bebf0660a144fcf7d2a8c4a2a061d9f08e6c2676f49757708ef8e1b0a17a8a3c8547e92038acc3d66b9778a2be13b6a464b39be5191dd2876a6de9797ef80aa04ed1e18da1140d688828cc760fbb13fc81f80555d06324300394a9638b3f9ba20cf739c7c14e5530656fff8b83b01e3c4cbbe5dbb045b5f090bc679d5a58031202d760f7f6748ccb169faedcc9992ba0e2d817171f4fa23159204651ef353819aa09697fc418fb7b4636d681ed75b3eead0eb73a03bffa8e4f6ccedf8fa2c6ca5c936dd83c8ad7f0267c7790bf5585906c13a9be08e896bde28176a29109a738d65963189316d3efa0755aa2bf09cac616993f9a31383a708cdfba3eecc14e03270b62c7c066fa5d3652b230b9077dc80b74dbf4c374f86b76a6560f28ec8f3a3dd6f829fa8895c947ac065b259ecd23b67430ad0d42743c75429aacee50913a38d88052b5c53b19505c705cc615a089b992916709af34eb129b039e9a7055d236a471a7b5fbc179f06642005db316fa94d60cbb5f20a16af736775d84f0ba358e7b9524b9f08ced036cbb28d55ffaabf8e93c61439ed3f43e7c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h40b0c07ec4f7325981b6a488d50acca28ecd1653a0ae1b30bfa24166142733305df90e3cc103a31f76886ae9520c6a6ecb5736089c00e633b9161fca7fe6d21866045c3ded17f77c035b992233958ef415550db635a4b7ae8c49801e909f8691e1bb4ccb3ee5b7be772b01f0225e2070477c9ab973c3177c4f7a67e1c33ebf124081160b464bbc123a1e4fcdca78711799ecf064964abc5b37f8af0f654d08c52bebcd1c88099865de9244c943c7e49ed89278b15663d153ab8354842ff3e93f1dc68c779401af57bd212bbab9dcd570e58aab054fa7a5f076e2cb768d303a87be20320b0fe2fc6a0543172cd22cb80f9d08d9d4672e50255fdb5f3718b6480e7af4ff96193e5136e5a716fe4f8e533d7dd2ace8ede46603f6969f84b38a0f1daa7da6c8de575dba20ab543c4dd19176bea97a50f9e144258f05f9b092e8998832a51d3479aff14b41d7694848ac26545fb30ca0d13dd09484a3bc98dabb73390c6b6f12c9477cfa298d8f8394fd6e1ad6989569a8747fcc155761436c35cea3af404aebdff83c2634acce51e53b0c9513ab84cb4aeca40685f1d4e22bad03ad0736378aa6dbca82cbd9d4ddf223401b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hdd34255f510079a1da56c3b8ff114575e909700cad828edccd8446f1056360d89943e59b7f40501b434eadcbe4159322e2394c394f7df92d6930aa2502e3931505ef9d7e6003fb23bcd9354280b78ac6a17965718759175132795523838c0f10e45eb0158debf1e21d1f65f79b06172820a535104677f1c4d19a93dc2b5604df84d185268088571816c89cfb652f345906e98616ef1c4127cf95b901b43e1231e2dcfb32f67347d92229e80fac9cecdd2ee8fbbfcc513948805726b0f1ad8e27de310556c77811dd44dadd62b2068f1f4df58b1e69044655cf21e03ab95ec5be59f8ba576b47df62ccf3a0867ab32c8ae3a9b2f8a7711d9ef8dd4690210c2c55133b9c89db2864470957ced2ad41726c4b65da3533a565b19c4a9c3976850aaacde7a420d12962000f1c7c3d20a0f5308222e9178b4024b699fb7325489428a3002ef8ca29da0353efb536af2f9834b06dc5a912030fc5e510173fefe40d7fd3a90c99dac9dd7cc0aeb937729b3981a4eba007a32ac44550a7842fc1a2257a901266986f93ecc6b623181bc434dea8d70b98472715294e1c53473e355f4ba7cfec8dd54efb453d4ee336fb0c705d6268;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hc8c3321ca2714842246b2fdf1a67ae4bdbf16f5935cdf6712f157e42af65fce38c65b95a36037108e812132458ba3d3e8a38eef7219ee6881e912808d5ac457f348b085bef35fa944f9b8042f6bfb3088344833ea5327c84b0cbc26036d5a7594c0d15b29035fde5b7c8c82d3a034b02a5d56a492da61fc9b540619a65d96996d3fc4360c036c5a277295a053dcee4b0f805567f5b3b2b4e0b058a6818284b011b005a5af452f71ca20ca19772867a7d1e3c7810cb3d482fca91d673635a0d4373ea94a71d35d594e7a5a7efc68e6ec2bbca255fef68da12b68a096a67df27709f71c40bffecb9eaf62404ae932bd6ab0a4499cb375210e166dc619c0c34ecae974c5d478a0ebc43782d2943e806874d8f2c03182267c8f813f6f3a1cbc76b5e4a53f9248b56a77b9b4cba7f40d07535cf69fc95f6a1c05ea1b92a7b72966175df0bba6db8c93afb42008277bbf9d0d26054fe910837239e8f0ba344d9ad637a270adff77838a9b44feffb895947a85c4cc107bd00d054d8434cde2393181525639141d2bd97f3ca718f14b57be365a622b0a1231ceaa2b3d525378f114c4b2b05f3b70f80cef5064212f96b547763ec;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hbd8fe8b2b7430efa0fda31a064f6108484cc93ab2d478f7cf260342e66ee7ab6e9fc474de5322775c13b02044b3437662e4aef701819061dc94d0c679d4835e0516f51bc282d53950e08a1a6ca9946c44ce00efd9f33cae557dd7017496aeead3087e794c006a02ee73d0c88367dbfc2008a60f688b947d11e2999319be6efe9fac471ac57646c92a0f4dec5d700a874c9778c65856075130fa91da03398980c5fd82ecacc5087e1bb6710be3167fead05fb000ed3926bf74b6550ec6d24ae0a54379e170ff267ba44107e4e3f594b0c745f466de506d626ba4d0a41cececd824a7a1d6c19b4744dd9c60f06489f51b70f6bb9dba2f517f9b77f68d187a48702e875eda865a0bdc8f52e7f439710dd411d69cda0c0120e2c0fb82cc5434c10096e70a31373c126e83dcceae758f454fa61b9d7b271d82b4cb235f5cc426cdbf43e8bab47bc1eff91a976a0ee33b79650a4ebee0d79339859a7c5141c106c8c936548a88adf509a16ab0c6d8ddc8098b45c0cc52feba5a740f3186be0a13cf3ad12295473e30b191ae9f7db410025ed8e78e6080b5660f2ffbde3638875638fc017dc09b20c3c5de7e52c247b0217b4ea;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h3283fe259d4371811a1bf4c55247145b9ef6fde5748d164ccd75d392b7e807d6efd0bfed44501ac6c6efc54e7f5fbacb6ec7fd963a4a1699adea9672a2efa1fded4bd6201322ef1ce7f0c061ac56609e5ea91cbe91c53c43fc7c3a912f7a583fb7b54caf1ecaaecaa103c01c205cd359523da468b6622f88609a7aba6ae8601f31535a287cf98f84c3c554b20e134c86a43942b2058fcbbe70903c33983a0460afb2199ca2ec850f6792d5aa729bf38a629e5e53e80569b0685eb8de149b46798ca4e2deac079ce518e3b92fd276392ef37bf29128eae734b7bcbcafe7c8273da32c7d73cd5334004624a3f3ea0318e91742552378c3c5d4f02d21f6210e1eb40264a59b4c29eaaa3636f7b02df7e6d77c8e9c7546e8399846bf9df23e12b7a48e28eb3db119347327dd191a5738deac5d8dcb1b2af31974e03f2a5076405cbae321b003f68bbcccce8519dcb047b1ebba0b778cda37c3b595b9d6a2da887a756214273e5fd656f1d8c62eb9dfd31d84f0a9041348cde60350404e94c98e5ae3b7939fb02d754c3ccd70a0ba3bcf639a49a7ead4edd22fa0fad73c5e75188c35b12eb348d658e03451c6dacae56abb08;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hc0f46c7b54681be0be3649fbdfd5d9c33cb3e2b7dc66fd52b85c50473177cc62cda9c790c19b545642c9b279fdc4eb53213284349f927dcae2cee507e4b1d69977eeef68b728769be772363f732dd273f9dfc8c3fe7f131e34bae69dc3724ba0088a4fb2ebd6e03a8430f4361a54ef6137adba7a741bc6b870ebdfca3b8b6e902f3aeb9a107cd84ec623dc619fa8c8d3cc8c53e4bf183266ae15f275ab81b55ba1414c09b9f9c2c251a47328673f78665d6eb81a346358e4c429c9b8fb83014d9d5e91443377cf5ac2fcbeec87dc4d47dcced607929f901df81ab4ae34c6a099b585a9bff345f3a81f3484609c02bee615eaf9006c6738c94a2b9673b8ccc4329b13c5acac6d757fad267555b4816f1110fd45f5e45dd3dce28e9a531fb2ea3d8f678895529111ac57e9664b791cc3bd870a1be7a45d226ce665826f137a7013f158b833774281a9fb6e8ce1d65fdad7b798d82ba3240df1be9adbb5e8b5477f178b5fb4a27638e55c700c99418c776cb02929445080a7d05312097dffe852ed2679c7925967d6f8ae001828cef1a9b1664f8a70f83204e294eb3ccb03d97dd2d1f08009a2d066b4539fc5723d93d296;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h1eb0a93978fa7207092728ce04caf20b6dc87e011b115426ffa2661cd5aa25a5daec089b3136c57d792b8f917888f89e38be6ed441547244c1c6091cb7997fd46684480e79f598149a7eb68202f7f00fe0f9cf1961b744ad6a901090c8bb648827e637ff1d0175fb277d397d3b93d11a9192c1e750f6f413a6814dcd2df47ced39336cec83e66ddfccfe1761141c497a314c7084b97f9ddc4654eb69493738d581bb78634f5ae8a067727522e15bb53ab7d5ce63e9236b9caf517028a78de6d9ebeaf57204a75d8f08ead1f66279333b5f2bab8a2cfa9300c5147e0644c6909807dd3d753fbd30c5d8928d35f133640d6ae76d0ce0f87760776f1eacb3f9601dc3841f52c447c5bcd17a6eaa6d9f5c1c0b5d2083ca0d1fd2349b4d0b5c21f9cf417e52433e4d15e0b9b6a7ca99d115d79610f32b27f36555441a1a1467e67f8163555a9d5b43306de3468bb2b2f49aba11b98ebe3ffa7ca42660c724cece164347ba20c7ba095a5a1836e8763c1069dba2fb4f7bbf646347ffe80e11130abf90a483e514e9d4c596c16e5e2892c751bb90eb124bb2e5bfb740cd1f1cf7b25ff730a098932b2ce65e01ca87d4f97d7901;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h976ad4af78cdae6bd8cadff989ac473c2dbad9185fad92889245a9e82e5ab038145c7783dfa259de1a57009fbb86e298af44ba585b46dceb024f896620b6c810cb10b7ab8f762a1ea07a715b6b0fdcccf1473db8e870c72f65d20e75d8533f93ef683596982e3e665867e5cf2172f26b1242bf39f0f5c23cd6c09c73b6e8c21fd1acc34148cda72f728ed953bfafb1312931b0ce2989ad0c3a7b9162734aa14374a062d2a9bf7006398b7fd29cc6d180df35de77fdbde2364a1eb6f72c0c19fbc8ccc456d3bfd7ecc62fcb7b63bc30f811cbd5f86da1d2ef069b2efe0dc741111a2a46b9b9224a962094a330b12ade3dad24e927d55663ac3364c296618ccdf84c2a90557bc8d02945460128e90d3ff0ea0b4cceb51b6cb89be5e73d70b60ffb85f195b210b1c4f5bdca5d0f175f86f6a7f511ee02df4251e5b3e3b430d0695903be82dd70fb40293ed0ff8635029bb83f044d2ce7baaeec425c2dd4d0df5633f816f0f661cdc232adb34ee730731264159c58cb873418ace6201026c910d52c7d7b5cd2edc59dd34779fecbb83036bc16e89ba13be67f5657e44762a2a69b18d95542c2fb8de362f3c0a74a69ac48ba;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hd69ce2ef40724f141af702cdc304f75003b871e9b22750d7e58c1f60b3a422a9eba6a70dc4d08a1e7df81f1ea2272f2bf37b646990c41fab92217ef3be799faf3c9ad6881eaf1ef9ded48c2c6ea54a28df99e8dbb547c0fea2a09f2c39946142c61a4f0d10f94e8adeb33f41dfa8e2698b90092a4e32c0823999fbc892cb23ee3ed87fff31dec1567022bf78a8073941eb07af5f54e28a8e8e05a48c47b3060a849d9c5c0a19b72d3900e7b3c8c0d03d25b6b69fec0135a94cbfe2cdc181e116b7d76d4d3ba1eaa09f7b07bb03cc2adf324bce6c70420e6596f52c0c0062ea5d3d85d0bfef4e11dee78f76e5febc2059ab3482efdebb7985e4bff3ec02b2d2abad3c9f49e452a484c335534992503f6cd192887f31930855b3c11fbbf99f2574eb6be4baafb5cb8b9bb8c6d7b7923e6b64f31b27dbcb85e0ef71ad4a44c23803dc8e2fcf7c867c410782a13c14fde40e31b2ac0957eeccc935506fe416d2e9872e75babb103b4731de4af27ce455d45c5160ca5f8fc258c21e3dd62fa04e8e00b192f7d8acece46d737de041c3457ba83fc4fdcdf041da87500fa5394d1f06e2f6455f3b29333717bb77a1b8d1b1c7a6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hfd84100b7400e715e50a5a8d69e8099ad0972ece502234b0afb36ab5fa245f43670f9f865e0fc2e29c77d3017f269bd1acb28d7efbddafdce4c761fdb050841932fad3760e47d71ca2c1c3600f280f35d2d4390b20bdd2cdce2293acef5416d29e74d1a2aea0485c27135c19881911dbb4de98d22071ac77410f59eeeabcb87754c44e2e77cedabb2f5d1341ebaee25db14fa256d28fee69d9d72adcaed078b845f04b2c83c0147946c98c4694eb68b155cff6d8698ac540e5babcf8a3395fd04bd461103fdc1fc08424f5a30e5e7def2f26d3e2eba31c7bc59483dcc8dfc4f90a6ae3ad3659480f15e2c233b5400ec32b518eba3530a3fff2868b0b6843a15a97324a8be0a4a3ed826028cbc1cc13cbf375e91f167d03f19ddb58110b2a9c4ac0e25d4f24c73f440bda1b5393287606b67223505a0aa4eba92fc5a77f2ed12402ce36c619d5653b430a329aee2d0d5fe4c66197f6a2815c6f2856440f92fafe42f7915e0ae6f6b1f49f432d75c78df021c60b0eaa9e45a1e1ccaddf887ce901351e862e82e4509b2162a38318e6869db61e3957a489214b8a1a3cac3bbcef1e25f2198e36f2a80e438d8fe7e244b76d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hf98e8be5f65092885f398ec98ff977e79d6266622a3093b657d0656e61f6b656ae84ca685c8d0b5416f9f51e628a3ce507ac75f30358cbe50d8e5e296ffffee60291991842993b0dcd259744f610d055282fe08005ecd878738af896937831cbd507f78f468b14c1deb89fbaae5c74922769fed8ca2c44e4d1bb31220eb6c3cdc236371b7cce3429c6882f270e697de817bb708a76259b307845edbc64486a367dc1703a95aa2e35d43669b71151fe894085a8611df9c6a36d38dda95530b23c5f2dc8a1cbd2662e8ee3409e182405e526eb97199421df9ff479bd3d66a9232dd894732483d5214d2cc07982d301614031249acd07d23211bd3df78d59abe8f78c5d1ed8c24e1f52ae78b93efe5566a40584e4079772d3c9ac3469892c9e2b9b60f0328e246f83cc145bc4a2191d9c6ab67d1432e187c4192c79a553b69e5a6b60bf355449ca6e19e13d9b36d43b1e73aed83e45f50ccf2825ec67790398223ff977f7e53ff52ff8462fef6e28c4cda386c0cb049a5644a73c3d1996354731ec7170b69ff7dd71528caecffad51c0127d78c0043b1292f5d8f2314521db931b83e5f1a2066a8bdae3f932dbf7dfd73a8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'heb60c86437d15044577604ecca7f2f372d93707028dccba58b007be20d90bac1001536f6b13d07d262d4b13eed68c8c71300c6b41a15b15c42349e12b9309d9b100254fa9763fa05d0126bdf5968d373d2424c79a7802019e5f6584a5edc33e3b825910e53aec9fcab23cd6f67f486f4ebbad7eccd429cd117939ba996d14f04017f12650e817b3fde555f6a4aadde50a1c88697a3b381be165943f88a26e1a9474baadaed9f0e8d9c497e8229d6491bfc74ac171fd11e6dd8c894a2ecfa9001ec8c6ebaabe9d0e34ef851b05db88c172213fc71b94c9d5114613e8665e23291c5c22bc7f386222a1f94db466427e9fbdbb5caf1661e5f22caf12c92f2562532c0bbf03e3c0f05069d1c4687fdb7fb01902a5245a344e12b60bd756bbc814126c297d9baafc389187b5397f82c0c86ad70f474bac74f11e9b73def239a38ad44975d41da21b637f0554de30a3fe56d08f3422ea82561092446ab416e903e575c9636bb8e72d3c0af23fbad2c5f6f5acc3fa9ee88a1659c6dcf2b2b11cb20c659431ac76fc7ac27ccfe1f9d490671884a72733bc044fb7ac91e3bcd636c41e317d3dbda314f42371695a4cde0cb1f3e8d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h221684fd381efd7c6961ee99463f98c047ece76e2d1b81f3f66b671942e64e47e0cfb1e9c02310005f2aad3af9e72655015197bff1fcbe27abaa660e1e1c93069d7a5a792beefe638e95a6d93865cca18c450d9434a22c46d16b8beee2aa56ac6b33b746c43db3dd2db3f6126e5e51ff51b21fa18b324b577a4dd1e5c27cf3102e2c73317888e587f6672a55f52142829462ef20fb0eb5c9f6ed3f16b06c4c0ae53833da5a3bf8f35a66f2022eb073fc1a849f9f3bd96c9b33ee81ff31aab6b34ab64c879921494d725045cc3e56261f843ebfe50933d578f8ca1524717e773b7947bdfa7c93ad9ad485a319062f9c61a4b101e3af07d89b545044f52b8d71359216aefd1c8a652600d51fcdebb1b336164c49ae4ecba0fad328527770acd14c8d3efdb920159c910dc541342706a568a9c756cc952382b64ff9a653a37e98cf84ce260a9a3a14a9c868018501daa389d31ae13488e345cd503a615f8237a2c3c441d3d0254c4685b254ba246f1adbaf65a9d1c3fa2ca8d9f73d13c3a793c70ec81e1eca9b09fbff8e81559a45e02290c6808ce26468579083715eadb55eaecdac65f6778e9aa7a675228945e08d62a9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h590ae60ec78d9764937816e6029d1df900ccedff158aca29e3984e869788df2cf28621797d30910b4516fb8825ab417aaa5111af54d5cffc16904f3c8a85f365fc10307437ad0242132e2dd1eb97d647ccb8fa2347324e5cd649f265aabf738810c9862754f64f7ce1ca68d5ccfe48cfed93633e60692ad60440cb3f75119305232a81b543e5e38d224933fad9a255f96889b1b82cb30b7f390595b68e54d2104f3a0b8737385214acabfc9b13d0d07292743344ab7571f1bb59f6918db3dc4fbf0187c5ae6bb2f11662ed0d238fa657c1d9720ecb5d0c1715a01bb9127851544fca03cc7e497bb4455fbb4ce4fc1a825f686936f0c7d140fa4969febb34c6d33ad62889e330a5d301180942e876b43df07438a44350f3dd06130546228b2b586efb8c7393ec9cee90c48b045a3ef81fcc8e2b2ef5e4df646cd9cc9d73762a403d921fc4e1be4f954a9e1d5b62e9a47d8ca226e5fb2bdcc998b61222bb22c0c9e4d848dea0fa85c21f02757ffb01d122012568352fcb48deac4ad18e9c8444936c89e461bdbbba232ccd02efe84a639386935d2dfcdd149ec2472225636d0ce12dad2fe170695490d9c88b113fe74882;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h6d23367fe864b58c3840857a12ba1c8259765b699bfb126b82a6745dec580e467e8da7108bd13fa8b5848018cf5502d4c18bb765608cb1950906c476da3b995747d9dec04437927bec4b52ee4faaefbd9c7b7b2becb59079765fcdff7bae8e6a4591c3bef5bb2228cb1fabaeb732c41706512bd3a23f69ce5ed7d57f3994f6fede6afe92da6da3c9f8f58e050edc4b7dc76db28af4ef54e2854eb4e78accd7420e28fa4b2b182359e3fcd67e25004f5027750365a63f76f85952f0de8b4c06e91248315834f0d3002082bfd0f8879f1a75b7d2c48e5c2c11b5900c1b7859bfe1021bf0ccbb9ca06cdc29607f1a68684884f942f6318c8417da933edf22080e49e72ac1841bbbb1d97da603b517a5b6b9248c5f40046eed947d37bdbf244b8ae682a9aacd7c700275de92472753aa6c42a77e1cec4bb72445a6c44edae2fcd8887d001a2c40fab00b72113fe9eb178d36cd82a02bda39a0a3448add735b9b9389053e6ddfa194a906ce2deff7a1de60180787b69c781f3306f742f54b6ab1f5e1a9cec1007b939a647819d05702e82bd00be269d760807d97a4eaea7d6f7b2531770281ed4e2b40af5636c5d17fce983b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h2f78ca37a707f2350feb000d4b1a38a9b4c827288602fc7126cba54c5cacc669b1c5a16f00d8647db4e69bae6cfe7bc326121d40cfdaa1d9329eee954c89d9837accc5c68fdf410bf025387a805d718f5731859907e35cef8ae0ce72c25ea694b02cf6d8e40a3bbeff488847ff773590796007058e44915c69c42a3965875576a5616113f48c8e4a6fcafce907bd3bf58e5f7cf2f51c5458c8e70dc12c6f24a7b545b1fd8e42df0014b9425dd0640a5bb65b9cfa596a9f4dfaa5674832b0dd264967ccd1fb373ab26960333162f34264a1b648e9a177226affc8058f08b79a52fc08a9567a50ad835221602584ccc6c20873f6950769fb7e0e526c7f4417d61c664ccd40aa912c2ecaa1f3ccd96160673d4cb82e1433bd5945dd0e7a669d94835f1e5701c90b203fa64438287e6fc61a14e52fb6bcce6e74093f015874a2024c81b78194c5b8b61fbde3f16616b18aeab492a240f092ebbe48df3c314d87ecb9a50576e0ddca8d76e30270f1c8e960f4ce6b3221777489febea57e80d94cf6d12cfde7f74ef13b76db858aac6e05f55d70655d5584cce0a3d0eda330d8932e24139d1b06a2192fa5953e509be6ef52c6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h4cf58c9c8c66ee3a96ee697a9d929578bedc73ff8c400b77b1f0452afaba484255a03f600ce7b525cefabb755775fdb52aba7d657c8940e36049f1625e300414f8ce9ce8b98f25a8472cd09ee56dd94258e1776d530053e7dd1f5dc9967acf26f8395a2d79d8998ec16ea25be9b36477d38e0583d495ae8b52e56abc971f141165e047b384416c06ce7fd4eeb5c0031e0ecfff37f46fb93220393d9d2c18c929503c0f36ea36dcfed32e4b5575dd5d8890cfe73dfa1deb3c86918974d619fb57347b7f6f0c8035054baa53037abf2390d1490be6840bdc1180b5f6593727d0790af62db593061324ce71d67f6a76fab06b14329a81837def3c928c11495de8a8b6f980884ae6cbd9efc0bd3e66c8a4cb5021f0615adb992032156a763b8a31db7a17ffd57b3f4a9d1e09183fd96c487062549043bd7015b8b3876546abb9464347514a17595d5b3b037160f682e098e5c90fde55e321e7ad3b86fa57288183d64038173bec678828070c66e95a8a3dcade8bb864bda7141ba6717df8b1387df56d7ae7e772888083efb613e4e02a777e74fe674c1111af100236fe17bbd07d4d40c0f8e1e03dd6e6b541a3348c0010cc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hcb328f2e5e8fd0431074d3268743c262a175cf431d5c0baa6b0170e215a74202cc367bef5de5cee517958561e4be4a5612fee5ebd2efa4851c2f434e194b8b7fd07f9bba90b4d298244500badbb0e44bdbc7df5786a4ddec7d97eeffdb4f47f71230af5a78620316bac75e3c27a3ff4c389bf13aa2c827b61a510c68000ff6c7533a6247c0a146c4d48b592a9aede438ec15094f29b49c0bc13fc6bf5ffee6818fa417292683c38b5a6d26da626ec904301f91c386068a6caae6cf50e520d3f34244ab0ac5a0bf3b5c743bfcf2263cf5592a55c7973f3556fd8aae5c5a2e175d91c1040784fe6c327e77c3cb6e195348e1672aa0ee6080069f869b13da7a9662ddde9798c00038f0af6b1935b56fa6363ab965050edd7ca5aca66813e67750413965cc3409fe68653898b9da9f149f2c04fc2a581471d0536c0e4ff98d963e5d23bed168bb31f05bc9ca553f396e4596075c47373715ac96ba948ee15d53b5c777ddbd9d0b9f99f8abc79f74d5c8604cb3398681f7edac5411e00544d22d77ba1a929ec1ae201c5ea7f59ceeefb02ffdf585d62beafb84112a334f1de686413b645e661e39f4a8a10935cf3fb596c68c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h3412c75207ab22170db925f7bd920e83c345b27ef6f6e5c593c767c4556f32be50f9e33c75cb31be4cb9a3dd849de58fef1f2d2a01675be54a6cc7a0088273b69e9bfc1aa3be026a44cff672968dee78e688b59b8a757c2ffda744735ead10cbcc834afa4f517e53808bc4512fc6f34b68508bbd9ba9db76c3a812f07a5cb1ab8fdbc257a19d80460e529596a945119b9808b3cb48d96a2eabff5fbaa0fc6a15cfc3010223b5af46129c6d23cbc0ce93dc9c45687f031f8570d7f74cc596d83eae636018c30df2a26350b7f7130c23be7b8a5fc77b8ea506c2733742f473fe0bad1d81f897eec49526802d59b4e117719bd57d477c122bcf17df346f040e00978663a119f2431f18cf0630eed5f7b3a77ef0e6fefd90d3273e780799901b41ec5aadd1d5f03cba32548634714370f83e0483902b0bf3b15a7e60e6668cecc26d8153653b2aef568528ece680a76467177102a3a0c141a07d5cbfa0e61fa7e299114aef5930e212decf4edf919f3af66a73c8a8f3c34378dba2869b776ba2342b2305553dcb15d4d64fe97b8b0a28716479a8359fcd2470f63a6acdb11d8398fe686652a3808ed5f244a09632c23bf896;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h7064088f2fc1d15c1c473e98aaaac3f131103a24e1bc51734a6d45cf122849c44b2fbadcadd8754c6e136bcc2f073220b5ab08cd4ef7f05a4a3ba38d8a094f286ae71145bd63af3605e58bdf122ef372a1e0e1a0b2bda1463a7a75129aeb92f86d40e8bc5e113153de336c6ed39b9b524d5ab57ce459f1fcf580fffd96569e77225525ae0b3eb46ec9551c2e153bf59e3c2df48a29607811579dcfc2a753109bdb56bff660b62477a8ba0eac14ca5c9d34fba0b47ab3414c418f7a45cc41c9ef91086d8df01e261ab4de38cf64c2775529d245a2a679f8d0c3c4ceec1990d324b29584481d4202cd832281564f1a02542e5d0181e8765782a4f039c7b563fe5c4e10051224f5aaf2b3b6a4a531aa8921a3b1b4ad2cf2bc48687df10ca0ed3448b8146b3a6a34942fb0652ef71c5a5a1df9db067eb5bb55d0905d1a52981384ef97f5bd1fe2b4eeda8832bc9ef8317031141741d6c0b169ad56b1471a85429ac5c92d8935d532a540e989e95c8ebb6ae4e12fd1fc7bf0ac532114723e63ffb5d3a14e44c7eebd9942bcfd7d14d0ffb258fedb078ccfe3a11705686997110fde7eba2851a92798b32fe890561728df7157;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h29ac97e5f1c9dbef209cc98cd7f32f99cd9392656d3fdeea948753fb6c8661fda100e90c1f178da34737fbc807d860617240dfb28b5ceb0dc50461e4ce60942a597ba85efabe7ddc1769df1c54a008208ad754163cdb36aa6771d2525debecd6fc936f0df3f80a48b401575d26c2945f2f1b16ff145b27ce93efea43a93ce566c12dd71c762b04e01827be3447cd0bd8b07152f74e9f698df5b82e9abbfc8410d2aa79ec4452a67120a07d1b5b04676f6f8d2a8187a279d63b217e28621b21c953def2b15d9771696488e4ff0f9341949c03d7b035246314eaaccfb1988c84fcebbd921216fea5289bec2cfc6af0b9c20bbc380ae9143f5951898d292f122376b4c1771870a98f0b3872e0b18bf7f27840eb6a2ac0e995b39caaef8087416e28091c133276e5807d324d4397621db8e1cabffd79f3192037c9b69e5cc38361675e1b2925065cda050eed72ceda32d24b626c6107af361053775cf83f0097fd882e38bea7db7d083c356353af501ee371efc34da2506264c1e2a6bd109b053c6fa929d35d455227e953eda42db4dfbc83671b727e7b6ceeae107f069b78be799112963a52d06123d9f2c12ad74af7e8e5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'hde5fc80bf2d6295af5e8f43a2d7a920c08af028113236c5a570e1dbfbdeab5a23337978ddf61afc6fc664d6ebf7cbaf2de913defdac14ac62d7bb07784870dc72795ef844740ab5afe00a8352863f987a5b992cb136a91d373c205169e9c0a4c60ef6226b4ff6e177d1fd73490b45d7871ddbdaaa2558c0b2cb2554e2ca7450324b38577af9d3303150276ea298bb889c7428b83314d718af7af7a5cb797c52c66192354886348e54e2fc712c0de9e8faeec06bbf5676c53bbd768d80cfb0957533c141c3a1dd3319d965a78ac667b373e16ffe49ffa71c87562d697a5758ee6ea122cb6074853695aa15dc61fe0b7dcf57c5457afcaa708e51ca1d7b969f38d9432dd1417ffe0c814861c7f56e522be48f5db266b2cd38e9b7b243f6acdbc4b4cdacc1c277480698f340b5b62d16d7f6513a73c3135dc00f95033b68830eccb17e5c57e1c307dd5778a3624b51d42c4db22a75cb467f426e8381ccf6d5d3c2dd1d6dea7e73c3184f1925e12dc51580bca40452172248ee4cbe9a0844c2e514f9c6900626029bcf169c6914162fc4e7d070b96b4d0b02294eb5dba0bd09339764476f4c7da4d54dcc39ae652401e9448;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 3456'h907700229f2fd1ec31bec19d915de921be232a881d56e7fcbcd7bd917d179da8b3ce945e4723737067a48e474555162967acd9a8c5f2f5588fea592c344db18841322cfb9ba4e1b825c6feb2da0d1d64c0802fa93a8ef6ea5794e0105804352af38cd92ddefc53920b78a91a4ce8897ca6f60cb453f843ad75caa5ec00c8d17eae178e730ffe7b6902885dbc57b4c672227e74268164cfb387b10213c01da52352830d10989327acd98938ff197942e8b21fef3a1d9e5ec434dd3884210e45c403449842cf212e94db13974b281bdeffdbea6c749787e042079c54ac22aca24c056eda5617a25c9063d383b95ffb36196f738cabec26801b84e17d573aaf1ef436d310a356b420e9433d9bb3022815770807215f8455058334869684403c4b399a920bed661522dab86c5459120d1df80506b99c2087f87444091ec2d5f388a27baca521a0b16bac113f3782d94a92c3c23a739c9800a278d036cb94b901d2b0f90e7d4698c558adf193da94a7ac182b20e39b8d7437fa5a02beece08aea6a7340766d1291045265220c9c8c46b7f255cb135f4bc6d6b556cfb17774f5e410b76530cf09a97c61f01ff5b06efea4c5b8;
        #1
        $finish();
    end
endmodule
