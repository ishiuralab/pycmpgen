module testbench();
    reg [12:0] src0;
    reg [12:0] src1;
    reg [12:0] src2;
    reg [12:0] src3;
    reg [12:0] src4;
    reg [12:0] src5;
    reg [12:0] src6;
    reg [12:0] src7;
    reg [12:0] src8;
    reg [12:0] src9;
    reg [12:0] src10;
    reg [12:0] src11;
    reg [12:0] src12;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [16:0] srcsum;
    wire [16:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1799fcb64e1f9574f1bb63e78b4980d522632b958e8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7d011618beb5978d1465ae3fa3ef0d9f81ec0ce6f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15b91f85bbd2c9d1e17dd5a948c7fd10d2168c85cb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a4220cd304295b0282adac2864811b4c3e07c6299c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h168897cf94e724ce250a1e31fc733d5f5b0276d40cb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e78007a24dbe773259924f9f6438b8b989bed3a4e1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h173e3df985de32516a4d88ebdeddc1eae6a17433742;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hda8b7bcafc6d4a365d680264afefd816d848fbbd87;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3a0fa8d6bef65fe476ab420e448d66878f3a37217f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13ed20a48bd047856b77db5e6cbc19d7b76803d66d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc874f878b62ac7e4d1ad6ffbf51753dd0b765afda6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7511d8cf7f0d563e7c7cbcda53881c223e71fe51d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8fb2ce558d18a809c9cf9b8f92c764fed210f4ad5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b412f348091c07c41efa25365196b2a03c23dcc2a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16704c5765f408493d63f28386f4aad55207114f992;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3bc1fe5902a3057d3b5d52fd157864452faa7372a0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2c123e1449a56613f7359bb68e030a4fef50f6be4d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e053d5bee8e6fe6a2048e74f3083ac03e6258085b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he99bc7eb154dc1594c2e8037c96a5095d1609aa478;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1487a135688316e7e67eb6ae52d9c86b3d3c1ecac96;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b1fc0b9062fcabab71f71c23ec1840768695cfb04a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd26b0402fea1a07fe0dc93678f905fe4435ffd7af0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbc1582a099cc17a058b6a751999686627191dd9e2b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18d1d64758958e53c4981500beb0a5ffcc6ffdc1e68;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18aa8431e3d395e4b9a5cbec5c96aa0c56fb717ad4b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c57f23247cfa52549007d3462257bcd6f1ae980843;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1af38b43493f165c2f5db8b9bad2e9f6124662f0e39;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h52c6c1453fbcaa3b5ac8234881cff876ef8eff032e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f74ecb33640e22b80cef848ebc28fc2cc0129b6392;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f256b585805daca15a9fecb424f2ee720bb3b4e890;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h101b6166f05bfb9fc126af0c548749978625a8d6cf5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1658eb488b0a63cf5a63531ca92b51189fe850237e5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcd5ec9b7795bc6c09c5904e91d29e29d94b720e394;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1555b7e01d0d39febbbb1089047f795b64ae0b6bc63;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h694ef82826f7e7be266ce3cec1f3d9bea79119fdc6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5979abafdf8e6a469583e434981e7fa29a9777afe5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h164d6d303f245a64f24cc6f78f93e810e30c2ca1b92;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ecda38ef3217e519b2941ce443c2253e3a5f76329a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hab5dfcd9a3146dc531646dcdcb44b788aea3bc5831;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ac87e5cc34965edc8f2df9beb898d15522010708f0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc7739de1540ae6b2d91bbdb6556258bc8f4c058c39;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6dff40caface9190fe223d415869b619183387136b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1360f36b5fcf540d8174b9c6eb5f286ac5eeafdf8a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h64e45c4befa628f607a15dd7f762fc800babe792a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6d0ba948ff97da80fc2ea0ba3c6019649715aaa12a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h69760165384ce2f157fadf2cec1696be1a52c709bf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11279a228d2bf96ea61f043fb6d9288d5906493fa72;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h174054edba0c755aa2e7997218a0d2292fd5680f5c0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h172b6ef59c186b112ca6e8b50294a0035a409de2e34;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h141c3eb5fa7d9584a3bafbf44715d83816e6b0cfd7f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1519eda726f012ef84b876dab52e2aa3bea6620b419;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e8ccb83664c68a1a7475b2e8e06d7904a78fe07502;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eb21358acc1e718ec4f62e6ee4c6c5e3f9cb13fd55;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h192210ce5015e43c5b0f2bcea8f1246b3f40c96cb08;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f3b4c39f767ac2106c2ab87e3f508ff7eb3d98d31f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbcf8bf00a8d71ccc4ca0553285d6db69f0bd4d3e7e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15ea1ae7a7e47267056e6bdafd57137df8eb6e8c406;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h191f2b031e8c3c84820777c42a46e79a035e0620436;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc9ae0425dadfd8d8fe7120d7ca245e76effc4993e2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15765f6b98756b234af7b480fb739e2fbcfb95001c5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc25ad533f992098ccc7b36deab6a41d384bdf2f29e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19e58b74a40ac9a656fb94fd626f8c8ff37500bd532;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15b820743f9d86d8a4037599bb979396c2a4be9e355;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h152cc80b284ba233512c8ef7faf678c2a4ed58db32a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a4020774c1e0b6706053f6d7a9bd082f2002e4bb2a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c3e50d72d31f26572e03bc8cdf99baf5ee58cd79eb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5f1a3c5eb7615dd264a7ce5d6de3b1e09dce1d12cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbdf1856b26f5e02ec5c08b4ce04925ceb903d8544b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6a81e8aba78d405462b9428ea29ab66b26d751f9ae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h888dd3d3b48cb1b36425a23a8d6acd03287fae6df5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15d0ee05b9fa1ea2c4f2804d83062e16108e108bcd6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha13de7a518fab829c344f879eacc58e38b2e8378b5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16aa8b8e5e657e8b6a413161310199ff59d3dc0fd5b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h108dc1de230cf868f1b8aeb45c151e207b84eff72d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h22f932da9f72e97986c791a39340c925c835d31c92;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h714148a75d2bcabfc55b7c530cb718bc3bd40aed81;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fce7530d787f8b16f781aefda6279ed8ae2dd0d25;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13d76c2791648d55113cf61a3d62c9f4b98f826368;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4115928ed47c476656df4773c7b7acd58101127dae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h479fb676675af0f87a1c79503309935671d02a31bc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7c48acbd857cdb5e7766952c0de07ed354ed8e3761;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbf03ba83027a5ddfe0b849a8ee10433e0f990adee3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9a7dcaaa5936b0182e923dca95b074af5d1302e640;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c38241363692a1bf92d7d9ba2c4ab396569cc6afaa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a49473729594b453b9bd27c164d07b5d96c0597084;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h110d8a3a1e072a886b6d836b3fdaed6d4dc53246d0e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h135dd94b37e027248377b390eaf3fa176948daf8053;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h182bec7a296650de49f909fbddc127096fd2b713ee3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he5d197a95ad6d1f9092c850628122780ba623f04f1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8da12ab58fd1c6a8dacd69f0031e8139b7d650c013;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13d32a5af100eecac9135e1835645e82aa7392e2651;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd30588fd5d89f6b5b86d6a269c1ebc32cccc33c154;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e4586e609734fca680548f69e2b1cf750507bb8fa3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h119ee77c0b88403867c4911757b7f11b4d557c4eeea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16548eb1a0d2fe63e367b8565dda99c22d1c088e352;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19e331a3ee4c180640b82d01bb94dc79b934f0fa0e8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d40396c78939a3d6cd120afe0bf5dedf9c541d9e3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fb10948ccb20bb7bc1269f434ec6f5ced8726c9a23;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18d51a03cc9e1dc882c3e4440c0b5f1c79c854f98e7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ee9b570dd2282d75e15f1669b39ab5dabea99181a5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bef15db0d958fdc5e2405dda2d33a013f1d254ca85;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h418e06fce3e0cd7af1d55d640928d214a2bd7c4416;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha3d68501706297c6a5340d553234e5cef23f5d4d93;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d8424025a77305f4f3dfde881e9795755a9c8cb08f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfc436b92ec234688bea2906087e20e6f3c03f63513;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cff5427b29808e53b064df9eaddd529425057ec1a4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1999d408f9f37d3d2f6b3bfb158bf5878a288ea63e7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eb6d6faef1278889371b982d7c77ed2efa667fc901;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h141812450d1bd9d6fe2a1cafaae8de090210a647a59;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5974a2144e99f901ae02987c4b6803b508dffbce92;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b0a468bff82ae761783bf3c4765a0be3b7a5f8402;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h48f541e4f7cfd507327718351db722f3c4c65205fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14efeda5aa0bcad4423b9d0ec830433fc1dd4212b81;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7358b3f4bb5df8272a1df0153b1e0eab580b29b220;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h95e7dd4f6aa14c37cb6c747f9684087fd858b0e88b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fd8187be74e04fca6968dd2ebb0f4f8ef400166d94;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9c4cb00a2167ce3f5d752ddbf03c8424f8656c1ef3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc1334c5ba340848980ee32763c190d31bfd7b1f1cb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6200af6134bcba54a67cb97acb73d3dfa4a8c9e96e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h131ebd3a6f43a7e2ae074fc616fa8781ed622d37833;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11a4b98c59bb5696facf76bb13c3b7a34b2f77b92d0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4ab2ca867ebaeccb16b16deb33626f3763e75c6cf9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5c8632af89abc9b6d03efe66edfa25bf87714b164a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1866da4ea801a5b849bfd31c9f56b0fa42050fc1949;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ff8e797e688893c59c939dc6cfbd29cbadf1a47688;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3c7431b6f2eaf0430e2208e86b7bb830c2dfcf381d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19a75d4be8e212b77569dd0e03ff81aacacc84439d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd762534c47b5de101d5952619682eebfe2a0554955;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he595e09e070213cff38cb3bbf857cf68230d3cbd8d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h81dad0083ba437508f97bc85e56f66fa1831438799;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12f0611eae740af9d464a305686bd54b2d7a7ce5402;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ca0922f71264ce85b2e0afe0e14d312c80e6dc9dab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4b4c11fe3e1a6809b20fb3aec34ec1ff89f46ffc46;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1acc63577036684cdefb4e566f5d15936f9821255ea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h624a2cbcbce5e64ed9a22a9363de3d1a8574dae452;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c384ebeacccac044e4a6c191c49b8f2fefc1a95c0f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h186932d39e2610424e18fb651ea5a567a1d66c98ad9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h97e58462ef704a94e53fe30798c94c89a280c6c89c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hba32f093badbd727e6aa3278d7d5a4e759454b6900;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h134888442298f93e1a403c590678fe1a0d905abf9aa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h43bf57f93ceace70528b7d7f3cfff07d8dbfa95d28;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b593a7a1c1562b0261e9c89aa608aae02161604c86;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h352039133b6536df7704046d2b224645a5f66f187c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2633f0c648e335f753486d0087dda4552d2a9b3a60;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h132195ff636bbb0449d3009983cdc4fb5093cd5ac54;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6daaf757e6a091a55fd5de29140573d232edbeac57;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h93ec809ae376ac466d2515e89c5230d358708311c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14aff288e0cf92b6c6564c80afa1afcea4709dc917b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19eb136255a0768e92f839208c08b1c814d79647f4a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13ac2ec7a2a7fcea8e928bc40917825787b7006f1b6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h169ed4c502165f2227978792c52eebd7cfa51de9454;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dd1f057f2dcd6766fa092e0396d0e3a06a4da4594c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10aedecc12cb7410e72635e80d858be3c94a399735;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3d260d8c2123ed7c9dcdc3a166352aa3ada44f4c4d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h87cca04a4ec11f3eb497c84508c255693b6ae7accf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e2bda1030273919df27f1ee8598be903ae79e1080c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19682f0b421e9577faf39de9a7397dfabb1f9860ba4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h472d2af9a019e3eb6eceaf3c0d9d38cca47a482338;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1004545da9f81e169271d4dce31a0ed983ee3f3774b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hebd17274fe0003a558abf6306d905e30bc0437160;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he07ed5d52751c155d25e9eeb9bb3e8b987175593f4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e574059172bcaf7bdcc2bc827606a96c59982bf596;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h137bc90d1d678a2137afee3cfbbd02866a1ea969a63;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11cca6e186f9af920bc9e5332b9d269fee44c7dac0b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9f720a2b78a1fe9944fb9af1e775042b922131352b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16d1e480390853fe9dd1934625bb30dd40c8d40a709;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd6e40ead29b9b7644e647cb5e6447075c8e54b910f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14b8199824252a04d3929e55b5d0cd83ff58a1db557;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h610b9a72c4bf6a3ea6e35e5a7cfd8492f0a46513ed;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f7298ec67ca468970079a07111fc154d581c73f68a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h852002525e484101bb8468ca3c59fbf06f5881999f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a73edcd48fbfecdbc36b6c7fc7286c113e29759f3c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he8feece3a50685da362bc8d5d805772b7f44797b07;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h137d6b5158026ee8c9e12d22c23af2aa5b2f721fe46;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf810d43db0d77c05918f244bb454f8947cd6876b5e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h54d5056ab8652a73f1744e0c1a6920965f88e8d44e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hecdf950a80484351d5461b124f80b64176f526e816;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd124ece36630f774268980588431468426a01a6102;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b19c8d8d027bddcb950496e802da7b2445d681c35c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h143fec40f4314255a834820a85ade99195a14332ed5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hac68e0dc3ef1a1d5143b1882451a47a17ecba3146;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h55401391a1bb60e89d91152c1e3026dd4fa8596c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5e810169b083ca78191de3375394b1ddaad5578044;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17a397ced19fd19cadb0b9b50aacc8b46159e15d96c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12b49cc78f05b93f691845bf0057f55bf532894ad67;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1950ebe599bf77da45758407d26ed35454c6657f9b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a8136498278688de26261723f6063368164c154da1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h190ea3fa916ae22a2fb4cd364502d7c4dccb56a2e9d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9ac93e9ff16f2a64cfe2e887d704175d55ed5a476c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2bd16d28497aff40b0cd8f6c1f1ec3b9fea927693e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a1cf4fd8f0dcc8a08c9440374139147f8d6ebf8b81;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9a078a033479e613a9e57a5152dda6dde00aa1b967;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h80aab2efd822899c0f3d14c81d7e8193ced212ffc1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h172f94336039fcc43b1e7220df63d51c53d0810c399;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha5c2bd18a98d17f904864873f6bcdb846315d277ae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1df028b9cc35b667aa423b453ef6ebe243e4de4c072;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17e0f8f518344b3ed1d64d5c47985d1106d90b391d0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcb7b77251b8f97432ca402822e397111d2506c18e0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f59d52ddb5fccadf797ed88d658fea570c483b75f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h156b7736319286ee1cc544aadf0332ac6d6ee1bee72;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1178e7f538dc48e0d62fc2f45ff332730ad2c2ea6d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e79c73d076a012d2ef7070010482cd6b1fbedf91d3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h154fdfa1f993c31c9e4df39ff4aa2404277e4b0ae0c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15d88309ee08e931e36fb97a8ca809dad8321984ccf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b2026d0dc79a107b2f1e36be7e8e6925753dc77aef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fe205f0f730c982864770ad595f3653d1588274d11;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3b4c2a3be2cb9580d23b536ea85f935922e6e0cb4e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h130dd5fdd936187414b2643814b0eafa0a156c8efd8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1015279d03d257bb43fe3d37b2855b8b7ef7f713b4d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hff00e4847a9e6e16ea9c184046cc17e6cf1969340c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4f81096365c1706194818f07c52eb022a7505f950c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf2f9cc2d88ca179355022f33323c2709dc8461fced;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he5cd8ba5c85fad4600e9d9a85a82da93dca26475fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5d2c398c436d9c68c791a18c34c6198d992ebf8363;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hec69b0d38e0f569dee67673986e58b225236ad4dd6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b54f856141e5cfd17c73644dcaa4e8c8a96a153890;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c48301cd4f2a954d16993afc756eae3458ddad11d5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h396d686d052893774290b9a26925b5d5b59ce24cff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f7d7ba2428ce5ce4ed8c253f3a230251e94412eb40;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf0b2cd775bab34621854c1c126f0b7a93e600c635c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ce207d5a68112d12424b3dbd63a8cc12a72f2d2fd7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc70afce43de2012caa076c21b557ea2faf8d7ecae2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1045aaa9ddcd3095a3d180cf9bae3a677f72a58a94f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10c1157af7b5b127b0694508060e65008bfacff4644;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14e7931e681847c27bb9389768012ad7c6215fc01cd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aa0b18ac4641563089bde4444895a9702d59fb3f11;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15c154dccc41aaad99ca61a2452c413c5cb7a7cb60a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2f192696e8c5d578867e1cf07eb4fda1e90618ffc4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h28bd0bb83ac70bb71c241a5fbbd0af51f7c546a8c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha5e0fe450ede5769eb23982aaf1d04398859f94d3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11f240be12bd3f6700aed53a2b1b9d55f827c3fdfbc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he19c28ef8d689beef163c59ba4e6ad3ed08e9907ba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a28e5073377fcfbd459c92fa8112a70b2dbff899ff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18cc15b5c7c4ad8b663277f7dfcdd2ac14862b0a083;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1edbcc90955f0873d0946336eaa4fda4d5e74872d46;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcbefb1932532ecc9d9e0fb8deb86f8779b8bbcc066;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3af585428c76e20723243e81bfd8a5ea126691fd62;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h143d7d72d72aea71ede75826e660a13686aabb5d8dd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb125c0f82aec37d5cb728678f7e7f0314cd73b33b2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ca222fe4df204579e582596c865e4a77e360baf4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h198ba2f3e9bcb8b7bdee496bbee33cc3fac2d819409;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h34ddbd22d49f92895f8b071399d5be9962582f1c58;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17e029b480e1c07f3c0fb62361318e0006d8533c995;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12e8f0b6443743dfa480e47f2918c8a50ff68336e79;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1405c21200b6e93e36615ae2384d7b9a94a94330415;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fc027f4982dbc783fa90573353d548f88f6866af19;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e108879c0a832fea98beb3e483ecb13cdfffcd8cb3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6a2c801f334fa95a403ea16769ab93cde5be9c54aa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf28fc6133b8b8d91fa71cc8cf4019b4b392095026a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d3b86433ccc47f48a8156c23d47e9423569951dde3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h113004368968f5df0c7c2b04fd8548af6cb8cd2132c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7e9fc439e8e3c6bb808680c5fc72ca24d8ee1db5c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h93a1d7ddabe6fb32e2fce447743e838ce71cd8bd84;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbaa1821b8dbfdb1f1eb2410119a8d9fa6be29cefcd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfeb9a6e2e1e9b324875604f0c8b79b298bf14ddf31;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e7204c52945775a55639d60a403ac729f1f07efdb7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4924ac77b4a8a16f9c03a041802a7a21dc44cdf08f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f0f0c925dfd6eff2be682c6ff22e8a8ddc745a0f2b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdc24a6071712cd4ed66c898f29133a72df23495007;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c8c51cd07edb0016378e823eaecde2f5e6b8d7f23a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eea98a2646e018dcabf97e75c1d6e4c626e37beb84;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hebdd2f7e6ae5962040041fbd115cbcfb8426ffe52f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h128777c63abe8d0d3db743eacc07f537873e0144b60;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd90a7902ee5b8819c1f8c3b5783298d31083c1fd36;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c3fc85cacd6565df6b16ecb3f80d4576b1ec8f481c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18bddaada699185c8abb98480ca46afb9245ae55e66;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c5a7e002e4a6e67641ee23a9ca262176813f8931c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd2325a36d7bdc3e29407f996de23981c793c91702a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19a5edbe29fac2065d2efaf6f10413fc95b551aa07a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10bd6e881983f2fffd07a6299886fa797bd0ce01167;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'habb653adf1170f0f0bff6303d15acb281b6fac6672;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hca99d0e1ac7030f796d7b1648dcc584f97c4904a7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h942fc2ab82f41369a43f5845941eed1f86fdc20a76;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f44a659826f904cb2203c9efcd2c6e49949db3df2b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18b8e01638cc32c4d521c03b5d3647ed9ebb6f9542;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbb2ffef2f92106cd002e1056e82400bee560fcc0d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d608b362cac9a4882c4238ab059ea7fa36e1863963;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11d97499341d568ae0bb295acbc4eaeba8c229a91a7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16d91bf63d4969de452b6fdb4f0e647637d9582f79a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1355efe3bc56819fef870630e8a81f29edac8885569;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h505844a0b386ecf020bf3e212a14c93836d73e4419;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13ef9e49e651807a728c59ce9a92805e9fa215ce86b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h179ada6c86212bfb18dc41fc57b2feca051efe08db9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e84574b64d3fafdcb6a0513ec85e9ead33c90fc65b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10486fbf266c4d6ed11d519d097a7e137022798e622;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf7e9597c993fb8b498c2c515981aae628d92fd2e4a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h74f152aa6d7a5882630d2bfbfd36afceabe2c82b7f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c7231330faf06524c221bf187ee8c166407b47509c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13eb7b7bc07a9d5ab9a7c2d88670a7eb38729f9a76a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16072c1e9d94302b1b8a623a03e08e4e45856ca601;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6befcd4c734396f4a166b1b80e87c02fe88442fa56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h61e595b6875b531b3299161ebfff7b7bd499299414;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h65dedccaf42496d43c35dbf52c47e53b44949c6bfe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h97cef02275f071a168e0ae4404142cee5b05b48dfc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he51e801fffbc91332c9fbaa90afc800f802d7f21b5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h101f4e77093dda5e71de8f8517019c16dae904cd32e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h244237ef214852def07ab40774a5b5d01c98afa280;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17a464b1e888820cf90e693bd119cdf28563a87c28d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d59e5f0675c70b7e41ffdd73064f5185751355fb0b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfceaf8e09aee512e2ff97160f6690287c342f52e86;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcc4f588a1ac3a9400172708a25ecbdf4a898af63ab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h442fddeb440a1603b9763c6801f3e0954f74f618ac;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f254b72249be4ac8f21340490f0ded3a2ad4537c4a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heb3900c35fd5b16ecaf84b2fab49a17d886fba79c7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h140a82e5391a51f4def9a9147e20e621aa24fb15b06;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a2ab943685a50a9c8970252e08653ed4b7a971b879;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1692f0706f78eb60acb197852c8d60ecde1d2004ef3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1780d2a7ba7e48c20d201f93ac411ae399254654a56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1685a7fceed804658a5ae604b824d67b4bb671c6c03;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdd2573e313052955a41b84f14abff9766b811e82e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9cc06128bd6e74f1eee874d36b3a56ea18f2b53c31;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10eb416f794b29c1d63d13292f4c70447ce2b036ae7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h123d45debcf5b879a119ad4742d4357b04392d8aa9e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h97639232e47d6a0ddfea74fd178f13a32a611277d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18fd39753b5bf743bfdd41995498595266108a827d1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h994d3f2e843783ca69476344ebd61984eed106cee0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h367db44f35ba81284d5e2359838ef1592c3ebdffd0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h42d9c8b3d3124e90f9aa7046195a143198a952fcc2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1de01af27340f0fae630790126d4ea14ebf6515c89e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6876d6e9bc30ed1acfbc015f69cb0e62ab34913b7b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cbb92f9f8a15a8b49e5e7f6dae4761441688de062f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b2cbf9d82c5d76f846294519d7ea4dadc2f158dd9a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2035b615bcab84e5928af868856c76e6455b3f1bb8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h114ea8671b17e723d3f71dd9d5b3c69f5066e254fde;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he3168707c38d7c2e1f9827d216fbc83bbcab51b55d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdf10d5a767541eab6e2954d752f184fc7980380521;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h85d7aec5db19bce226faffc1cfff665b01a39fea90;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18bcf3c6d53f7896733bc1239c26738e378437fe7cf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hed62b8654a9fe706f9d073f9ccf1d43762eea80b5c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha2306f6e97ae7909322be793a34e1da6d88671e23f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h97f243b76c90fe0eeb85202e15201f0c55a5171035;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h327d99289536d2affb25e2a84f1097f705b7358313;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1648e93531700902057b6f2848d752eca0f3741d532;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10f55eb5616c853af8d3a1a191a6b40aaee7d73c206;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15714b7fea86c72997eb966cecbf91da493974cfb03;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h983059538798e506f99677dbb9cf9dc56840b7ad90;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcc08781549e485c36b6a9a3bc829995cb4679d2d51;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4c516559699799ed3b273b62adc71d3652b3239577;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb2fc1cfd04c10d6aa6735f008ce6e6da7bf94ce759;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc2305ab8804ff885ccdde8ec77e641c3ff8b8795aa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6cb608907b44a35686bc2e74af9e3abb3691ff0ad5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3c18249ce4983853f56d89f62591bf5035918fe1f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h116128fca8e9a2655890a45fac2436ad485f6b9102a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h161f2a24241f7084afcbbaea6e2e7dd8cd90d54f2b0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h124a62a234016c21ecd657f0a553485075ff7bd9fbe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h144da2850555813c769797435c9f837cd6eefb56656;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1962997564e69301b55cbab00553af781cfcd1390b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbab48c4f271ab067f78e69f69b2345cee5af458839;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hed9630362b9f8f8485e1c6a431bc4d16bab5b10c9f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1857048821370e2b080b5902614dbb1830f54e7fa5d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14b9842b81d7e8611bd5007ed0377acc2aec8702425;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc3f60d43eebcd78c093a31c5034b90d0cec8ef8d16;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4a5ad3d5ba78db3dd84683220b6736638278dbdd7e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11b35aead6df8128933e1ecd84d9da3d3fb24401b0a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9e150784bd3e3f7cca4a5efb897cd76cc7d04db989;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h99d262ab101d1168a7a90812d1773b3c5ca7a00042;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a3ebbc566ef4aac7e14814bcbba4ce285e05ec9375;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16454350721a0de373f7a267fca6b354909ac959991;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h678705d14cca4875b2783556f088ceac4c00b39d39;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10d61c3d71514aaf6b96b4cd1062ddd50bd19625504;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfad70e5627091c9d48af35b6e8a22ed73531d741ec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc12cd519f119fe371537be9351e2cfbb19c684761;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha28b9d07b4b1786f9c417f74b08ce6081cd53b6807;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19cd11e46f05cc068ef617360cc93443d28712df25f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h122a97a447635a8880bc0df9daf917a1b05bb887113;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he581dc3b54418910ec3d3e533c70de07ad27e744b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h195413f894cd4cb77733abe37a585e26d326f5995fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha62b7d2887af42c2efc3edb2714f68a8b209785c35;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c10b87f2892380b4c997313de0484dbe33d2970c2c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h31b1307fd607d57e2a954a15996defcc4fa02b7f1e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd748b6455b24195467e59b305656ed4eb761b89739;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h616f39d89be4c4e2896f74dee2bbc992d107c04236;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b0e4ab5b8ad0f6598f171f64d50dcc41535454d21b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ab6c6067ac9c4fac3be2db91511ad3d66479298030;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfc095869ed9a879bd6c9e98c9c0890b6d8f015ef9f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4eb8505bb86a32e43bd7f3e7c7e625c2047dcd9eb6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2c14580530a97f8cb22b90d934087e3f83bb368507;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d87ae6f9ac658f7e0ee190c80d9ebc2ba31d322908;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h166108a79ef8ab0aadd359c27da4d84cdc29f24c5a5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3d4891455db57489bd5dc3b3ed5495a85566a398a7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8340792a8a645a8175a0d4e76d7580c53e45260306;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h161536919943a9afea8116e5c256ac1e84ae2705816;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h139b1b005bedc88b89c6bad360e285139142ae957f6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h84c93fc5bf6087d6fab83acdac46ff83422371d97e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h50a2dc642aab7f2603c76776eab5ff1cd8f37b6f87;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f852047847ea63dcb6c10fb0be0f9e8de2f3ea4a9c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hda5b876bda4d78e2e5fcc51bd81f6196dae275e58d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h53b3c72b28d6ce383884e9020066504f3a83516dff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b4cde7eb8cb98d73f0624d637cb3ad77ee82bc8a79;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5e41549d33f9123889307e18e60dae96838d5ca1c8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c0b43fbf54fc4793e7a67d3dad6cc46783659c0ca8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h127ab58d695cd02ad56e6d3472b6ebf0927f25c0626;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12c7930042007ba1d941ab0836b797b4440be59c75c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haa30df145fdacfd0ed7d92f864153d30d27959b6df;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h300df35b32018a6a8c32ef1e129d28d2183e5c3d38;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he4cacd8e78a7225d472197e846e85e8521e2c90c50;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6b39114aabd8ad9361a6b9c533718e766d9840b5b2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h52b40632575d40617b3dff9549f14faec0498c5a07;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfc1b68c71136c2fe32d39622b5e5fb1a33fe77154d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1389fbef81991d8f67c832188aa6cc874da7d9b6689;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h148bb660027b99f7f434827335bd7691a27191a8a7d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d9b3d117ae91a02b830a3825d2344472339e07b52c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17948d1d809aa404a7f46b9813bea3356586ed566cd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd176ecce3767308f87f90ee215747a5023b660829d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14833e515a9b7f61fbde61127c7db55ff7f2460e984;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19bb3862895a7c3003f8259abece297a1d3f103b467;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13783e7d4b93811a97b1567e4116361eaeb3b173166;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h197e3f301ea33c0016d0216af8e0bef3102eda29d5b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf52f91adb75ced46ece33b19bd5701a0adec686928;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc4e363aa02896e0e60a75d9fdb78670aab46d2c606;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h58ec3ebe40fc4a200f0f8ce1149ac856776736b0e8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbb199dfdc8006685cafb3af6d78e3b635c6ded3cb9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5adc2eac90ab685e5b24eff2ff115cbb37fa7f3936;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h112f22815cfbf2608b01bbd889f301a8add51455170;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16b4e6e015caa16007a1898fa5cf0158c1b6b4ff17f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a05f53893c1bec99aeab37403d3af108bafcf48087;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c070e9267a5c4e9f047f20845ba5cb9f4e0a00d7a5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h95b2e9fbb44747ef0e3eb1139760f869eb65078428;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf2a1b9e1d786e7c1ce1068fa5e2163a872566d9270;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h50ab3a597370b2bf72273dec0b3fe2f54859911a95;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfac512c1efec4e49d8d3004af0f132677edfa4857;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12edd203e6ca56c3cc49cb53cf22da85a0f659f8832;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18f32ff9c4e01cb491392cb923032b08ceba418c6a5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19f72530a70bae09ed6b01079f9df668b71ed64a297;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17ca6e4677dc7d95fdac4c25cc3fca49f91bff4b765;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4727be6a11bda55c76405c42ec25fc5b14b7243b7d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fb12cfc76d653b16d48b270f363d668427a99f3182;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1afcad4255d3282e650f83e1f8ce6851eb1be5ba1d4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19a07eb7f2dc691aebbeeef19d0db8874ae07a8785d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hae83d949ac3e69f04f04e8e6bc45747675ee9412bc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h118ceb81dfd7138e3fecbe3f7ed377f9648e810d453;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17172311200adaa0231eaff14bd46510a2baef904e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1635db440796cb354fe03845b41f81b8d436c8d5cb3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2f1b820fcc8520be4ecf99ebdc2a452013d09b695b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h171b92dcb9764ae47e465a8dc48712fcd3590d3d9e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h38296d76a9b86dc23016d37240b2eebc72cfd89a9f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h174f55b36989d0d1adf07c0a13aa68723dea321ab38;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9e6bd88a1ca0d7e46cdeee8e0ae17d9eb72b9c0d96;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb53261b4ae22c525d8f1c87a601dfc9386016b21b9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haefea2c6465b80c60d8318f1c744bbd02b218c1ff4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hca5005803332469ba197561067b292679aeb621921;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bc8a70bee9dc779f0b24dc08b200181a241fb0fac3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h197dbcb9d691d07c46cffbfff2fe8531ab36c87582d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h171f386eaddf1fb50f0959a941ec93914fff9322341;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h773d2af95312bb80bb39dd4b2ea4a75c528600daf8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1506b92508b6efb0d725773822e8f152b418dbe8952;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17800bd5f874865a36a14bf5bb9997bdf9363bb1459;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16111f42a4b84396429d57865e68fc9158ec8c2e1a1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c450e468e4f0fb4bdfab01742e741470566f74083b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5790856b638a69c51c794c6e9c0f3270bb7b80d1c2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'habeb2bcc129fb3f87b57e5585a69acef1000f2cc22;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha79aa5c92211e7dc0f8b537ed3099c995cf9e795fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12d6ecaa0ec788ad604c14175703e378a27ffc3785a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h171d57afc18d6d3ec2a9ffee59d27876763b85ff8e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13ff86e624c4e1df9ccf6c719c3e97dad0ed0633363;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f2b6838477ac28cd7ac66947a96aaffddcfdb58ece;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha0bf7f7d517e15696dd1bf31363a4733915be6e34f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf4e05dae14a4b9bb76c77eea3f196f70e0125a5ca9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc80eb06586ad783584d4b7d28f1872021c00f6a7cc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc0826dd47e6d4af6614610b077d72fcbd9407ae5a1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18f805f926212720a084317a022adc025e9ad4654fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heacc567b6a134671d7a91947bc03efe2e474c1c06d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h140e70e0b09eb8df16c334ae50e09eb0910eb10dd55;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h173c6b169075a9ba60873359dd4a23e75123be82f1f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h389f79e73c20960896600c723ce8c2b47084f08fef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfdba08fd0f71770447ad30c536a7a8c99bd1f0ae5f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6053d8a2c546d9fd210c0ffc1ec33f690efd5b0450;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fa2c03a2f136959756c6d6f9d3af9219b1d3d6a5cd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h22c975cb77882e923d08235dfe846b46c57fc455ff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3bae57ea35a8450a257f46a8144e4d8846cb500f49;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14b3f4898120880a6d4170decb7a1839475116758e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb5a316dd896d77e2c4610d4fffae6ce6fae20342fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h147727d89868076c5505129baaf6a155932f29762;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6efe23ebbd3ad6dab76ab631268b6e3aca5f69fd71;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h183392b36d769ff36aacf06e3e6b5363a671b6b67ee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10481f8ee94a4f6107f3f996488945556328dbdd837;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h237f1f05ce293328df327b918ed63a05d78d41a14c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd661b3116cdb45010793525bc327c43148c9425d90;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d9723ae91a2e11bf6810471307dae1bdef8a8656f5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he6230351f18dc04ea33542e96580d56132cb91dd03;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf1a4aad34f71fd3a651411e8ddc9f49cec8e943503;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7a2063a563f9fec483f5f4d168e0787a691dc01749;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16269371c5100501c5cae6a2d6169b5576fa397c690;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18a37a8258b3ecb2f7dc8b5983458316e70deff1722;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17a49e7604e6d8ee0845c9deb780490ff163fae543;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h107d3dbb18829c1e2fd5518455a88aa8736a74fedce;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha3d621b35618bfe3150ac55e05cd2b345adfe9371c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10c6dd702bb67bcc1ebb99f659fca9b0db55ef7c89d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hce7ed6213ec658ba85e16db23b5cae2f6a36eba04;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2d6dcaf26e0710c37e8ad5d12309aa926705e70a7f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb77b5bbab131c5c8a68894732774757751a026e757;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h56d7a74bafd42664501c987103b752b2f9f28a3de1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6d181831e2c78e629c5dab3f786ed5d8c253bd0956;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6699e45af87b0c4706dee11449fcb10ae9fa9a3f94;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15c74c32e2e7174098e1b95bad7a828e87a65906737;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1432e6c717f67ec4d675e1b66eef9fce11db7b4a469;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha0a5c6b51d82859239da8828747fe419322b360ed3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h57c364979008a9ff6d5409bfd04e2aa1dcab54c3cf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc064e6b20baad8a4280736622c5419bb8d8e3ae3a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc443b1e012a8a741908231fb64aa7618814c987aa9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14a7740730581feb5278047d081ede63e042ee3fd0a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h171944c733256d053aec9bb585a5388e7e600af89b1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6071bfb107baf6dd52716eac2b1468a83febe6c188;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hadf314bf2d29584f80cf8b7b5a980d6845383263d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hceaf462749e4f5069b10c8c61da2ecdca60b7ec82e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d9652191fee7b95c4cd980976a78761536ab78a7a3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbb0dd4d8b37c72abad6a24d34c1908679236267776;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha133b4b7b81d6944b1136d9cd70234df02c1af4e07;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h974e9637d0fde2e7f324ca72b2ba0cdc4cfe8f1b13;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hac625d23aadfb7d9f7998fdcb79ac62ba6aa4a9222;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb59ad8bc095a844d44e0abb42307bc7f9af21553e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h38597dae63dac1ff3af64e38d63647fa00b13bb9bb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1be9a9a4ffea8e16a618580b0ed03066dd5da267107;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f1a4a1ba663b6ef00d898b7fb1651af8df22c6930f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb3036f0cb4bf684fb862b59a08e03c89b901dc83b6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6ee98ca4d48536a5221977a59dd0ed102c66f2b78d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hae891899ec0e48bb9701c64d51fe3965f4b0be5967;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h24af87fd85b1e196e8d7aacef4454d2500f26418fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8068267f0f064410a091ef2da833be0435cf726af1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b383864ad4afe0bfc68c5209d2e04c595d5c6f40b5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb664818021f079d9a22b7c14c8b3ad240e4272ee25;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd3aec54d4e7319fa80cf5cd676df60cda84b4fa63d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdf12f94b8b5c339c0ba63dfac776a83b30dbef5e96;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fe8462bd31f5181a0e90c2ec40b3005b6bdff7f48;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1902faa7825f19d6800cbdcf3075db469e7bb77f7ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h174ee106284c4652d9dee54c849a5a346953c5b5837;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h513e9e788023f951743cba1f71cad8e7c4ca0c7664;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h74f79e35358c9be2acb89a4882343c48d97c003deb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hce15e671aa5bd3ce9a25e577352f3d6a866193e098;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h320c9b198088e746667a91d5d9a65f61f397dda963;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hae0c3b6a2b223b00a00196bc2f47a90e7f65dce13e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17d6f8e5b8e8b570a670cd42b0a9441c5444cab03fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19f18fbe50dd76997495e47840322cad29c6bace732;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc846ea2b069fd7c513925e81fd17db4150fd8075d5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h582948b3e3984bb4fc02ddc5fef062b23e48e26cc4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ec03b580f14a3982cb924e5bce24908c22b392dcea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf61a6feef0b6c27d8aa95e8108a3e3b59ab1450815;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f6648e337f0c08fd48289308ff20cb2ad0cfd6fcef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14c246c812c81254cc66c66e066254010c4b92e3257;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h180ffb340ee0f576bb883392d78cd64b11cca3ff3a4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19f988b46d5e927114c999ef0c940345d1cbcc31457;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e1cb3b74c534860abf5d47445b9c86cbdbacebcbec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h81ffb1fc6617ccc50abe82a69af591c957d9bc0624;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13559ceafa50038e53b3718adb63245c32342398be7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h472f93af36d3772c2e6085709ea2a55255a54e9dbd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h656edfd396cbb30d0c6260042c353b5b8fd1aa87e6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9dcf093995fda5d7bb3278ee8435f91e476714d36;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc3c92f5e09e4c2f4df3f7b9e28f3ed1fde2d8760ff;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13bec5ef97bc7d961e58055e583df834e1bee11a682;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6b606f4d8e677417d4feb0339bab99461e81798346;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d85dfda007fb3777202ac838efd478057719028525;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haced74d0e4c5e225fe51fd96bec43a728a29a725be;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13f99969cbf8ea2c1e4cf7e544f1559516e3df26bc1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bd23f02a0348edf4f1d9d19e16a7e5d968755bdf22;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10e0eb6b550b58874eb0172a16e91f0728220f014e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fe410f8fe5d45ba6da6935e10c000510ed4a391e8c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h76b1a407344ae66d8b21b347f9e1638bf0fa13785e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f2b52e66afd8d894b8175cb6120afe5765f5b0432;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12b2766294285bca83f52c62ecbd710eb5946130590;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h145e0de3fb9f74b18d9f0999482c1c1a27695f7b9f2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5fef0b65144acf419749c433f964ccdc3cf65b178e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h161640c021c2aa558a4e36e446165e33e4904df045c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10d268b0714c1877384a813a3b42648216b6f1abcd3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13cd73ecc6300254f47ec3c8049da14f32a2c49afa6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h75eb0157220a6bdb3dffbe666ccebaabde326e897d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h87ee1aab99f625f75d8eff4dfb04cb09ffb0e19af;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he1ca64d009d3b9d4d93477ea4d892412394b28f826;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcb1d0a375d3843eff44f231a86ce5a7ab48cb8cfca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h121adbcbdba3e452ab94a59f4e4dc76caa013cc43b7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3614e01a2f6bddc6e58d5d223620829defa03e4411;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13110f77afd178f40a9104661fd417dcf44258297e0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h187b9c251deef5daaeca20a6b5279d3649ab0eeab1b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h165eb1d0d0aabf8ea44f220a962066066ad38cefa60;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c02e8c3a3dabda083ddcaae6c1a0b103f0a1e1d97a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f44d0d79b0588997f3b7799f30ca0f1e3f2b838f8b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he10eb4ae1cd331c87ce2a4e4e82c473d6f5d2b25f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h121be4964984669d0ba8dd3df3b72bc71acd63506db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h163aa13a5c7ab283c7dcfb9a30577da622878e8e443;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h49e8ebdb0fd583c9fcec065a1598ab0f8f70bd8f3b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18c3988059307884298d3fe0d77bb597dbb44d3bd59;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19fc8c60f7918146439d22f6b37ca8fce015b0945ea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h125460a82b411df5100231bc4e5825ac7446c5ec9bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b1b057cb2775a5193dfae7cff0dc1a2904dd4e91c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11caeb0e4d898dca38cfdd2d26e103d35b6e38c694c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd35e01862660843cd44c2f54256c52d097b380d18e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h104825969987fb1bb9143a3bd5e77177bf0d450197c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3bf73d25f01c09f4ed99f9ed323c3e4d61a4c1ea81;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13cfa76b4fbbd37ea4fc227e4c0f7b6ccc1e7291b3d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd2169e611acf5e4d60bd14a63ee2b624aadb3dc2d9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h132ba66e4a8d33f6183180479841195715c98bc4621;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c764cb0155e6fdde52111a6d9dba93ad91c3759c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d9dfe43900babfe79e88dd7c7fbad9efcb11062103;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcad6a838d12259ba2ee934c1ac621d7472e2233695;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5cb862d870c031d66607229d1f6339aff013276211;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc915aedc137422417bdb350c3b13616da3bf76e20;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf8393a90daf4f1db8d5e692278fd425481a4a806e1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e965634cdef74ba9e558d0bfc90840c265f2390d84;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14c73bacdb78cec9602baee7b526d3ea70f86900b91;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h270b7978bbd25757ffe739927b933699ca1be41c39;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h62dc7a1ccc70565d3a618ab9df156ec45806669c79;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eb1aeb3912de000b59c12c98773b48ceb79ff2d90b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7401f2625ffce39bd53ffb3aeb0448d47c8cd0f4e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bfac1584e6c1963cdb735915e8263b45eadcbf6eda;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h39163111de2acbb6bfa17f6b4f29422e4a9f7aeb5d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h120ac7d523974a14bf4a697f1812b83ea58d41a58a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc7181f0fe5d65cedd33f2577acb4062fdfb9173fb7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c2e8d35bc6adbc9b3904505eb345e044ff74a4bce8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h124c4afa11c98a138beb7a2b93e5b7c32cf676ff597;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he13202c04cddc1d6ce9e1434c47dde6d31f947aa2f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15d23d922c0b93c3d2b9932bae4b61353b0e4341737;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15340924e1826b15bdf9ff7d9e815557293eec88ebb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h171c4e097d0b726dd76c777a272cbbb539ee06ae241;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfcd010dba42ad34c5ebfd54fa11a4637f52e152958;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h169e897150df7fd0a3e733e7abdfd876bce4456ccaa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8f14ead8558864d1bb23016abbdf1b5bfbc2fe499d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fd24e354e65bab938209020b8fb4d25d7a98e25c52;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc0edfad7b289af059ba67026e2f77292948753ba3d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e9df5297fcefbb367bd23e54c9b189c6f6dcbd9edf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19c708e95e83434714538c2a7e223e7c7585907a4e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h30d5f4ae1be7d4ad284ebebd86688ab01ab7e301da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4347afcc1e727a7f8878854a1bc4795083728bf25e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9a92b5bfe18fb00e9a517573641862ffc8eaf4654f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc7de6da2c3a569c5bdafcf8e6e01b862a5b712795b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h192e0c91a4e385429435d580f5b4b3656aee8e1810e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hed4836f5c81a0bd7eee589358608a1cb6ed062fe6c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h147089f64753d09b8ae1b72cef690a4cd0b7d7269b3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdf492ee4c99de7f5b4de2918c421255fd127f8aece;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12ba4132ef199a4ad265ae5dbe8fc86c876067fbdd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f5f3fa2eaa4708b3311604224543184db87e52798d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e6c095552f58dc114af82bf47286f27859e3e6ee1b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hae20ad0c4ec4e831693e6e9225ebc268a92e74ee65;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d93549119d5e017849d2af375933c9cdf260416072;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1366bbe3aee2e53e57a699aa876d2e482634b9d440;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he53abf94269ea7c99a8f722f68a6114aba0eafb8f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb9f07d3539c51d250e3c8e21ed7a1a4d512b998f21;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15d1e96f9129db9046ba56c24b421ac393d7c6bd7c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hea89001cdec87b41eccd289229fc8ba80d82ab99c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c38c5f32804bd6739c8c0eb59ebddaaf516c0689c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h198537f9ab7cf521234e9d3bd69ac601665fe327d26;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h184dba5dbdaeb4334cfebee1f3a2f507bab8264bc53;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11a5b764ee5df92cfe7fde3699e29a6b625c96b4b16;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5473025c33dafc115e79b195541fad27aaf2d3b1f5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a1d17df0d9fa7f8e7fb0e6b0ab405e5ff138d1501d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1197a0ae33c1e0f6653aadc7730935149e763df7aaf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h63b823b8d33985e5bad3a95f4b0e73bbbbddd9d2dd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1301ad14dc1f77cd84ff19401a0baa0f7241046ef54;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h144f7b5b7b9156ffa49fd9af9d0e28b7f4e8ca7204a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dc053bb8a2884fb3ed5cba105660e4ff72fdc26c08;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6842645c43b07983e9834ba1e246227e5f1c0e7548;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h964108cf614a2f332553c67c278fb73149c757faa6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfdaba788577cb52b1cadb0106d4e279422a5924fc2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f17a2ed04f7eebf65a7f5e710b5e7f52055ff257f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2a33cfaeb779e01b31c8e09e568bfac9d75efdeb76;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a2989c77f1ba1cc3cb35fe75961a4d1e1030e96a08;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb948ccda33dc3009cf3d2f312bdb4716ef3cfd8ce1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15f3c726d6befb6ffbbe699bc21044dffbe917b5241;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h68de7f9ec45f31c3defe06642e79014d73d66f3875;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h821e4c1e59145260069ce958eca8106c602d17dbdb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h249ebae6e1a7f03f11a8e8a1f2532783c293ed3be9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h33b5456bb1f387b06b4b47789b4eeafe91f1bba265;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eca2a7dd6f4848e606a75833fd097d346f8e73af3b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'heafd8896dd0d63e2cf7fdff172d4b8745d7955fda8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf87c6dab32be54442e908188ee4ae1c60d9ee8b94c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he8f28e8a36d2fa5585becd9dc33fccc5fbd34d3155;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7c0d1001027e9a98622227ff7e6429e1c915d518f2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h244b17d52534dfe7dd4ea2f14f5c1bd3663380d637;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1063d1ad8b7223f9ba02883ab34e45128a440240b77;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h57a2ccb213f67fd0272127058599a492f62ae6c6e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13582ec5e45575f1d21d938d66368c6d4cb0cce2eb7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1568accc5b64628b8b3cdce3adf0b132ef400b2621c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h159fb099bc89196708d276e67ce104d9b3b51f15f19;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1777131916818fdc8336e3a922e8443deacb817e1db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h896e886c313aea1f38260b27151bed07667bdb8688;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13b57dae334465c9937bbf0a6632c5e5f0314074fab;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ac90315bf3f50856d7260de213d46db034a1454987;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h58e869ad252500c861dc1543920e480f89ce6d095;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1dd7ca355a3bb59826799b84118e770dbf84db1eae4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdbd42571b2cac89b0dd4d4cb825f520a2d8942ae38;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b916da6856084daae753e1e1ff227c620a464165f1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h126438e641224a262cd3566d6002861c404a3dfe4f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d03bfc271254ddc962d063c8035c85f4b66c7004ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h743d03a2580deed8750addc5a986660752924045e9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16e62f06ccaa8e37a8b1c5286cd9be84ac5bafdbacc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc7868f007b24d41884db3ab3e22078e17481b4bc8c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d6afd3e2ab848611bebea8da77bfc6ee2b76c8f39c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h140280f19e75ce3232338807970168fa123eff6f1a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcbf1315e2f21fd5ecd7d85bdc904be759042e9d932;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcc56feeff2ca8e0a1da561526fbe9729fc3a861a79;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15cdcc3295c27e8792e9e3c45ad32a05c553dd51809;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h195353d5cb5e91d2bc66564da4f96267c093f88b979;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12c85212748587458454aa8657a898df1047a4c9a0c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1018b2a6305e491572b629c9e6f29e47497f4146b59;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9de69b6e7fb8235dd9e2447a20d8e572eb36474d09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h93a408aa078104147a3bcc4b71ac140b2b7b207e56;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12bd9d46c5e12f397803e76e1c9eaf814bbb17c35db;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c08d0d5632411dd465971dda714096c5ceca416c4c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1063769340e3ba62ce13aba66419f3c34654d76d224;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf15a6d3d8b83265f8d1ea1a16cc2d6736518ab7ae1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1eccfba26ec6f0b18cae1d479715c2c280fedcde7a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9184b6fb561e8a2ce32664a24e95821041abc79e7f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he3db4a7434dbd02cb781297e195272f727de424341;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hafb1fbbcf80b7ad3f23ecac9a0c5038d480b891b9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdb30827d56937c45e2229fd6dc8510ffd68b9fefa2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1bbda005c723d57a76b23ca9d278a472496d09a610e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h122a3d970b0fefc2e5de271a6e44c9931c037ccaf0a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdd85bbbefaa996eb7bd78a9cbfa85ea531c64eb946;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d34281b2a2c45138c7fa9a112ad2916664443130da;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha5bc2b96876e913a2555c5ca7d140ae6fed2f9fae1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cb0a2901f370f707c5b6f63450fed5e7ee3d89d27a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3bb688edcb2a0e53e636c1ff482f1abc4d77e26856;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7c5c6583f068ccb85ef0e5c0ffe8b3c6f450d19e3b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4d10412c44b09e33561ed60209db6c30eccd2657b9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h70bfdb4cb50db2191fc7174e7941af2c2a1cf76e16;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e6966e20e3e2b54b427b8f7030271abb2dd754586b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f5f4537aaaa35ae483ebdd45c957455dc33a7e6d86;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b39914e87abb583d871c23d26e6ef1b90d1746ec8e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14fa4c7fd39ebffa297ddacf09b1ee4bb6661ee766b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he73b47b4158d8ba37c87add61662ffb21f67f7fed1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h89af880df7cafd59b7fa563e223a9b2f5f84dec549;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd6a3296be928f03d772274a213ecf7b6c4cc94e531;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h269aa6dc9fc3c4a1024cd33dbc0c9ecbe08b286e95;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8821214569cc31d6cba75d0c03a116748fefddbfdb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hee1690a92fd2b4b1513024b3318366c0b57afb5af6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h117acc81d5510e90d523e53a46017199b7a8ccf2961;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcb307a46c4fdd7bcd11e80486f022bf04323a86aba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h116acfcd6370a698fdbc38fb7fca65801a689221b1a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he1d78c8e61f27e796f349e31bf5c1ca490cb2edb6c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h188eb3ee76896983e037535ff779dcc0eef042779fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hed440f8a2218b2d6f5b882474d543d56976d1c8d02;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c9450e8549beb944e41fc93c450fb8b0634e921be4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he6f2de658d0346d48c39eb631546e4ac1e2e0be081;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c124cdd59641718329d6dbd92c34da219c3311b722;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h122ac71f35c65de00542b1d2693fffd86a5f64e3ae4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he65ca769ebc27a78b64e14ae95dda479ab179886bd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h52c42e499e619244d53f34c805fad3f12dfc79eb3f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h519979eb05721b3ce005b46b8aa91961b7fa311917;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8a64609ada9d8f898dd997aa83ce358fb535cb5a30;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h157258ffaef39bc900d021b931873ca829507f5bc3b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ebe2eae755607b04ae5ace91ea2903a54b2794a4c7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbee868659824fd9512b4a0692740ae0ed7360907d8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13a4afdcc79371afd0cc72d9deec7949067f0bfc268;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9865b1f893f216a1388872960cfad97948b1e693b8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h83da998dc415553a45a36fd168da7ede6aa94765fd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16374133b4d18e2ca3b9e8eb1512e058e4cf5cf9a2e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha0937d8f06d6de270027730e2d364aad9d74dfef49;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16c5700f8f1addeb8757eb4705c8175a4a90e633c6d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d51423cf6a38bb95fcf1a15ada4aea3cdbea8c903d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd678efc776ed13a91159181ccf3f0d01897c2c2ef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4563ca05b1b0e419ffafa868872ee82c174ffa7839;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hec9502f703bd18f1ff95cd3d5db837c1689fd2dfaa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cb90712857542a696aa7043d1231d87dc04962cd8f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11b5690b765ec61a9c01ffe0eb93d75acd304c7e06a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b98e35feefb0c649d2b5d044260403fe68f757f935;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14fb3bfe69663655bddda93c54a31887fb2ccdf8ff4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7490982c093564df0647ac6855b44ecb351e17c60f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha943d995a6798692e992d7c4a4e8b7dc2ba724eaa1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h142cc25bde8e559c47103158b68c58dfdcf6226b924;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c60b33c4d1a113001b071083b479d4da239634121c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1361628e38b50b2e9c118744d5782926a91c233629;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd8a915f897b8b2b544b5a152bcf5628e6570a715a2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13fb54b8c37f025987edb35d3fdc2828617d7a71ff6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6656de8bebadf42dabdab661d47ed27482ad8a2d33;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h60b069eba2e5f2325eb75932d3444686562367c3e8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d9dea970d5ece7ef0f483315c74d420533a896f71f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h175072ffd39d5a3b057181e63d33d5387ee38385e09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcc96c7c788aea0545e49393ea7e66a062e3c90b342;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16f721101988b046989086aea30da7f3ff3b4012dba;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b41f626fcc33fb91154b4dabb1c66d46058426a83;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19ee4d593cd523a3ae3a6ec3ca5f7133a009fdabb58;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18ad6de3c828ee9c8de5c7ec80e80e0f8e6aad7cb3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ff39b71bec8744ba99ebf0dc433046804d18a8c852;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'haa78a2cb646fc991afd7b9f61817afaad391f6d0b4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6e1342d60f66916de57fd9dd414def528f45feed5c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcadf3352ce5ab063eea289dcceffd49c721657a48e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16ccaadd47579ef70757a9195e99230bb11ff7e0ace;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h77161667c2fda39295015d1378d3e02f4b024d465f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1244660cb62e2942b2e86cd3178ed601632b7b74f01;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h54080312dece79c270190d657f198e01a0e31792e9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11dfab6d5ce45c3b7c6f5e6664d550c4012eea7dcbb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h78a1ea4003e4da4e64a13dd75f1f0f35b6dfc6bb88;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17c30829b94e026541adf79e85697f51444a0bde1fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hec67702dc1fa09b0cd1aa274cdaba26a46149a7412;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf3d2220cda92740a876db5568d1f83c70d1b40df2a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1965391acf31ed5aabcf4a56cb3e3b3ef3238f26c01;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d2ca91a936a99a8abe296d6f24211b2c39b2f05f92;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d4e8870a7a4ce66a6ef10d4d1f67a3c247b22cdc7e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13fbcdb14d3ab972f3bab2ac20f8a5b3645320453a5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f034acb5da90bbe59d1730de0b1de758e1a810beb5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c409ac2c823f141fa62c58e53b6fdfca83ff24a4fa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h399b88fd9e279975e2d4a68c9b7237030062b3d353;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7e79b7eade879859229531135ce04a3ec06cc84b9b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha9d372a217a0a065c2c8bfa8b8ebd8286c1b1bea9e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11233d34118f06708aa164c223d8ed1a0262096b585;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc9e37d74dcc1750ec1af79a8ceb6d429af8210c2fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd0ddbc4b3a2ee037dfa70dfc27b3512c1e798f8c8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h39e6748186f52ac5d3649f0a9bf734d7184f870508;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15e9926aaf50694e1b410fb0db5fdc41b1714afa720;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb5214ed8ecab688ed03eeb60c4bbb409f4d308c17f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcf3ef9c8af11b46d801971360deef0d7c1f3edc240;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h90efa91036c1f4767e14509843d9cd9299e645e015;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18343c4500e7cb25f8a38d52453306cdf3ea6264770;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h80d2eab0d23fb092a2f6c7088f9deadefeba0fe874;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h82797c349dfa8888386683acce56e1e66244c61fdf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc01c867c4ad8322014b03b91cfdef3e2c5172945b4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcd53d71b6775d633b0e7996be1fb59f242e60d8657;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h738776f2a81d25c7d1fc17a9724ab7f8e47fbe7588;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfe02a2a862b344564557a4413293e24a7ff3d77110;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9b9209cf9485cba527c6b86085ce0868956fa0d8ea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11cf7c80e8dc1e59625c2a5e7a888e2f54ef23a363f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9c08de61417d8d8607b8345c79fe6a900ca8c204c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h99f75865411e5233cdf0be4bc98e9d7df7f35fedbd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h638218227d2c96f525c98077c0fffd5db8d04b2189;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1df2f6dad13afcf604c92301c5c6839b18b0874181a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4de57aa5687df47d8103c06f80377e1d63accca6d1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc88ca9c6402b6a6b0e57aa7799a1c0fa3fdf9d9c27;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h28e7795d1d3b036fb5a7f9c3c6bcb9df930164242f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha2a5b0e3fa6efc353bdd6a355e78225fe3cdbeb485;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18a651de9f8c9d9361ca6d78b5036496a2846546c6c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9a14355c78e4fb8b5c567aaf1dec81714390f101bf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hab7ca7f8d9f7c06b36368f888fc912052922556e54;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a1a19be788bec37f7cd518934d3c878422b7e24fca;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd4de984837fb125c0c244315c0399220a9d7cdcc2b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h271fe28a0ce5257b4d48c663b41fea4af06442ce10;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f137b5866e97ff5aac1349185d8e9fc19d14cc85f1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1521fb94314a9bb007de5e2cb085c4b3200588edfc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11bfb5d17fb860e20d632161c2e82135dde45195e8e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc6a91c0b607704071025357f00159dadb4a6d2828a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h187b8d8fe7657fa340ab191a82c7b7a78956898da0d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e3035006b9bdf9f65ed89576ca70606a3ba1bc66b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc3b465c8b328770dcbb519e93fd30d4aab722f70e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e00d5e706a8a68280b5a55e9567524599956dc7dbd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h132753e2cea5beac1d9ac458132991ced2a73a76055;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1203deb5ef1d8b3cfd37d6da4a3949759f24f6e9783;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19781299bfa8f3e7b1fa8c1967307323a8aa08cc960;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha02c2ba6e3ddb3c61d858d4a13679057d0d7cfb659;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h172f76761bd39b8315d0097d8e9ad185fd7b0f5fc78;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he2f0f7361861b214906c319c865893400cca4ea5a4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hda665cec78fb43dff7caf8f55e90f05c7da9e23c91;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hff222d10f170e4f039545d885879f81ba5db8e7b0e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h23f8fe8e50d38f9f9afc666a04abb73fe4eb5a60a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1aef2f804688cd5d8bd9590b1c97fb28d7bfa6281fa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h860df17ea220da2ba1c7127a35ba1ab8e7cf941c7a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h50c78c12a822f47cb64af35fd39346cbd8b6b30423;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h61b9994595dee0db4a54b4aa1cbba44cca06d459b4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he0cf58f0be5f8443e54ac75e080a1ed89e879ce025;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17387b99afb08d0a045e9664b1cfcbbfd0ebdcaf889;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9f3c155615fc32adb0723833850c1dcae4885153de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h151ea28b2e6bcf6344a98db8053d7d3e5e403a1baef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb1d4e04d71a5063576ffc6d9b3f4d9854f15a383f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h70259d0e603d02872e4cc2b8c453c6adc37852cc71;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hec8be7ac32df79b387c1f9a7e8701021f58f725c37;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf02c3aabdd811e34b5c25b33449d0013634e2c3e20;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha2d818c1033e598a328c8724d2dcc957f949fd6146;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h150693937b5c92a0e570b60ea15b08ff5c9ca2c3386;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h175fbfd43eb6dd8a43fa5d8a020644aaef36f84fd41;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19536d9610fd4c65d58c2054907a122c8574975a7b5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10ff66199da24f10f4caabe53e25a116886872835a4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha24a419c79e140c6314ea98ddcd88a0d939421b8f8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h55f467c81215c57eb7d06a9f311df54221a2d5cbd2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hfd16e3b43f7d9bc065184247c0d344509649fbe6a7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13299fbdb6d205f2b8704204a84012b67367e20c82e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc41a5d4f8b1c0be33c4fe206d059832917d70b7872;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16c21bb891bff58a1679db2474a646f1afe07cca748;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13fdf0e36fbc55a5edf54a0bd6331378d40b98643d2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b4992cf4bd44b77342f98ab65d470f8288a89d3634;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17700ad814e072cf8f65e92dd2659ad5abafca5c41;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbbb109032c525ea55492df57592eafdd1ed2d32b12;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12000bc50509c88aae1f576cbdf94aede8aa4634c2b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1198c382f1d941c5d19483a784ea61fca420f095a4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h180e34c3be3423e8c194aff18cdd7b2b03ba72a3cbe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7d847ac5b595a9554dc6f9d8445b43c170ebd347a6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16effd38a1bc156dae1133193f26914d35a600bc681;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h52d14fc0aa66ec6a420fed030f3e2b0df141307be6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1490967d13aa4dd7fd4d18ff913a9694c273dc781fa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1967f236ae932eae2ca1abe88dda59bd1db31539728;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3705ef3c1e1533e2958a2e2885ca482067851b7a1a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h126cebb683efd651b850458ba9d892f648d430b7394;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12c2a0882846b441a14eff8afefdd7bb0cf42daabfa;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb88f2fd3e83ee41cc0188b2d9f1e835194cd82b537;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h5f5b54fe7f27280146676475b52a5d5c606563a179;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16a135b5dfb361a7e82fe268cd04dd9ef4eb95605b9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h138c921292984481611c847faf48a321fd542a7609c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h50e2a0779b01a4be6e3949bc1dbf49cf881270c453;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h107397677b963c964c5860197c25c8af03c71f25c58;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h169926a21b6e947f2c0e8a96f8d76c7dab6f6db0d0b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha6bd7c11dc9741c6be27aa468ee2c357f73e8a29c0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10517f60ed713922c2142d3e132489384e8a226ec7c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d185678c6d857edac531c3f8cc5e12acfd737eb9d6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7c8635d6a47734ad9185249526d7794c7f41c395ee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf15b10fa0a332340ed9385541edb525d9337bac7a1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c3a221e909516c117454aca6f676baa11c2f17b1b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1866dc1518ec96e65b5c62cac155187b1329c9b61d0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d529cd17d94cb02618d5112b1e8d91e0a164e07690;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h8637a84d32d6095ee34162b2127223b34b3b951de0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7ed01c0c7a8ebef3c9a40af2d1d008bf8808377fef;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1732bb8f8c9b57195d417feb2a6c2053b9fc130c9f5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb99295742744c3926fe5aa4e4947ca847054763489;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6c8be8f0e42d94958bd737cc10991ccc1f7524cfc3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hcf7447505221d1871220674a12cdd4beda9f89d1bf;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h105bd19a19e140a30c8ec2b37b6a25f644d943f7e92;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf1520ed533472fffcefcfbad05ac2bac4677a1ede5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13d8acdbb52d23ec1937fe8844854bf35fb1467f402;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h138270d6c1d2bfad28221f0d95f06d7a63d4ff155b2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h45f626d106767c141639b465fddecb8565b1c6532f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2cfe853e7e80ac5eb6be2563d707f02adf8f211492;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h50cba19ecdcab2ed2653d4c0714a616362549df9f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11dd9985604c8b60be1f35777dccc322fbeb00d2cd3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h55798bcc58fe2cd9ab70f9d3a77a9211d567ab0cd6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h978319f6d27f6b77b8f7679c7b3da6502c5c753ee4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9c5edd8afea1c9234c5dfcd45025f14f42f4626661;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13cb47ff6c03313cdadc5c1b6cdb649f2b53c851b28;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb057009f1256622da97a61dedff5aa73dae6cba1cb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4488cec82986d7ac7037703b2db0c3110b36e8d513;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h108be4e704b794c1f8c39c6f6930a4d247d0f61faf8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d4c0647299baab03e0f982e0faef791663be3922ae;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7d0ee55bc8e0719a291abbb1294eec474083e155b5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b8a2e3c0d2896bd20fb45a9b8cb068f6e0ebff1d0d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h29f2987444fc7ad18d201220bd911bbc92dbd5be31;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11872a6ea04e0a351759bb3a3600cc73aae6f75209c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h197d00ea26d56b8beea07aab7d3276b0d5e34b393c2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16f728ca57f2379f1df5d7c46c3cbe76a4fc7976f67;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1be78f708c33a8fdb3858b2350005feea5c32d43fc7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17b77928b09ca1e1b30e57690506dfef34dbef85415;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b8e5c96e60177b72b71a4077b6d9de5ca3cb6cbf87;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18672ee8095e59b11d991bd15bc11c5e92931a482be;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h115d3b04a17b225210a63ddd7a23c3ca268d55f21a8;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha4fcb9658666221a532e024311bc220dccbb718e87;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c96a790963fc006d4332b4e8823560a5d3c0858cf4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7c1818e737088b9c5752261c86176aa2140e9eb064;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha04adea482c8d093778876d11bbea5f1bfd08c38fc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11df1d3fed5550163bb170906aff5a992b6c97d56e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10321825ba168afb71a3135712a5ff751706e39c0f1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h171ce78d4b65cc2860c9c9610b171179852a4dd6b3d;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7aa3b810518deb04b3a899b54375b9978617e31d65;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1557a514b19ae0d6f6de105b07bd887cb0f3df1cbc4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18686af305e22beb3b47efd24954ffabd3df96f74e4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h109d431ba2456941ebf6c3abca092b78ade30efdbdb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6e4c4eff95187959a6895aacf553b8cd1120556cd9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1486a058c31a7142e9d55a7829db1b3848c4166fda7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13bef638c8191ee13fbe2219ca01bfec9b31fa8c98c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'ha62d36e37ec2b023db242b09b0583d90eed12cc93f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1136bcdd0b9857658f7eea63b5cd0cca788ed174f80;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a151c668e89320ec48d892bba7fa47c87877402fe7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h108b8fe75822982432dc15967b97549eb6f4dbfa570;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h10338163cd4971849d9ce84f720b8b17de816ba426b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h131f244d6b7d363795440e5cf0799d880697e14bf53;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h59ea6a89f049bf46553cf8e6648ab3d24f987743de;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h844a39bbd6fb5813ed90d9efae5589bb5accdec15a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16e9a52a33a4cad90121b16d35c81838d2c0196b007;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7b0025dd615b661bc240de18fe3fb207eea683f3cb;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h145e4106896b4d76720de4407d886a98dbbe910a16;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6506906e436e711c9fde9a7617d0e0bcc5e73d05f9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h13d28d946fa01c5ea57dd921c885eafe5f119c10cdc;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e742d9810381da7efaa18df306f6d7e0db8701a19;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12b67a3c397474cd5761c1517c0a9b51a81902c0c43;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h167a7f168088304d5cf8588c160e80e0dc69eec1068;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ca9ed3de9ce3c24ada402d137f04cb8fb1dd5d32c9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h72bd486b5d22e3ede5b89802ab902ec384f34c7512;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h172ae52f3f7781f1b595b00c1f5261f6c46a5a01a86;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'he312c615413700dfc8e1aad69fa6fd8023c7ea1b7b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3d19cfcb0c0cec9ff51db6038c2d63c36c15ce0323;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11d908e19e991d75267bb2bf0a8928f7bf1cf24b0ec;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h14908f093ef8306812623d5b940603110ae3dfee712;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbd22b63e300b774da59f1a5df906f4aa3e1c9697e5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9332d1f6319916c5d7f13c38bf7c2313303391a9c3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1120865f3eb2b67f7cf6d324469140acde29f949a4f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h29b73355ed2889d079b49ceb4fa649b0cb2b089d73;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cbd3006f7d00d30cd0a41bd535562475ea0027ad5c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9ffacbf54dcb703e150da3523825eb070ec2c8c4f3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h3553cf752b07fe316fab5a9e98f626df5f15d69cee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a258c6b1aaf3430a79a72756889f1516fc1c1958f7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf3e88c844b8f2e64b06441de2145cb1203fc9e4477;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1e7fbcad31cbeb85ab5192322d5db15742f49b0d074;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb32b2d06034d739c744d691153dd9d18abd60f537f;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1617abbe2a893af7a865e104424dfc0bd89f724ffe6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h9911689edf0117130631ec289ef17e7e48b90abac5;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d9aa2a2772edc45d1e0724268af247a8e56f6df243;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1c442cca6432d06a8ba47822a743bba9a0830f1fb04;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h12e78eafddf723bd96ed91bb1c88d31ac1c4c46085;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h15b16eaed87b805bd4e0ae6b4385758f733f69a01be;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd85bf41ff4e1c8a4063a50f7999b6b9c26c49f2c46;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd27914ca1fbe6f9743ea6fd41d23d131ade535aa24;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cbd95c7a3cd765a4196621b2823d8aa946c95fc78c;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h6408dcf5b3d18f93fbac30b5f6cf1a558ec1c3fd19;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h11df1a33eb52349c52c90bc4b66b44a7667f1a0165;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h194d99cb83848531f4b6c3a51e1c36d4334df942da2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb1a62d9d7a9057df6707c92ec8c898b8482ed9530b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h18cd188782e75379b010df164d52ccb5a7f05f97e1b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1ec649d1e7d51f6e05c56fb805eff0e18430309d503;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h179a551c9d9a28853aa7a0461118f227f2d37425247;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1a8800deb4e24a8a43c59298918897041db841eaa75;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h7a6a743f149001672f6450656fd9ac02f101482c05;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hb34725227dd15bf3d4c8cfb7cb7e73f7dd8ee375cd;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h36fc45f4093f21597348d56d7f47fa787592eed1d9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h16373161b7348ee3b03217a6ba826549bfab9d391ea;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf6454b57e33962a6c562aab2cb4a657d1197064f68;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1d4a689de7f0816a4dea534e3642f4bb76c566d741b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hbd7019479db14d6b98ecf1a646334636920c1ca83e;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h115d535dfa4e851b566eb494a28064b6940095b7254;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17c960e96ab2c10ca6207d9952a90e8008503baa20b;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf0bfb5bba9258b30b0d66cce0593a97e86ea9734f6;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b11b06496dfc2170d398025072216f81d1b81ea6a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1b2441cf09827b7dbdc3097db2ae9fa5fb7047cd587;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1df79949c68925b20b7320b8339180a9d0fd78d82b4;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4eadf7ae890e4dab5a59eabc2da96266c172485304;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h2cf0ecaf4d062241475e740807a201dec956919dd2;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hd1af13cc8e4660a9735cfbb4dac330defb686f2e50;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1fa59a74fc23055505ad52aed12917ff919e894ec94;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdfbee14df681f32bb664a4d11ad21cd2ad5ef6effe;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1853c3a039ab906128ce035f351ae9d1f7e6bc7c760;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hdcc40bbf60bb4a26d58a32e741485d743ad7c3732;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h19b5368e84678354779b1f59cc32d44a819091b11d7;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1cde23a2b1fde2a7469ecbaf58819324651d1397c09;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hc5dd6a54d1d4457064db673e6b0e89fab486adeb86;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'hf4b7feb735834ad5a4d821cb7cb17bc907a3d06851;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1713868fdb962b62616fb2a22cd80b1b432fdb5a07a;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h4521980ad472d2cf6232e42a8e55160ba381b33880;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h155b4408ddfa1a0e0b749f5c328b025910ce53462c1;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1434ef9732267942bacf5dafcef6b770fcfca9b39a9;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1f5822d1fe5b6c60615276f35d17dbb947ad2a80dee;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h17767d8f580dac36954eed3eb0d4098a803e401bb3;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h451a70b7bf6543dad3d3a72c83cbbf41393f81ab0;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1380ac15c5f27b6bdd02d7d343fe568ae03321f5578;
        #1
        {src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 169'h1df56d3d87fa1ea08adbc8e75cb3faf5fa61e7cb3b2;
        #1
        $finish();
    end
endmodule
