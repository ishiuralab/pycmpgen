module testbench();
    reg [16:0] src0;
    reg [16:0] src1;
    reg [16:0] src2;
    reg [16:0] src3;
    reg [16:0] src4;
    reg [16:0] src5;
    reg [16:0] src6;
    reg [16:0] src7;
    reg [16:0] src8;
    reg [16:0] src9;
    reg [16:0] src10;
    reg [16:0] src11;
    reg [16:0] src12;
    reg [16:0] src13;
    reg [16:0] src14;
    reg [16:0] src15;
    reg [16:0] src16;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [21:0] srcsum;
    wire [21:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb9ebbf3d510fbecb0137568bf1fef2bf48045c3856e14ea885238872b78a0722a64bfa68;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fd948ea7913406c175e53b00d2cc17c1c0d33b99ae5776151eb89d6503e459f539d524d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb1e04d8f64798044128a136e35811ce08b9755803751ae76fe86c58ae64031edf0b7d098;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12c9bfe88f9860a110716a5f7f83032033b6504918978172f638f5ad1908b20e100f8d1a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc0193d7e0e28b5c0590ab5e724bc80feba8a73bb967bb5437357376ef69a4dd043928f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h38331b3e40fb3db5810d7ed786613f744da4008ae09d6c569af96b34217ec626a4982013;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h52a5347aa25c3317036505791bc1ad32da2dd6ce60a153fb07cbfbe867ff69ac6e07c13c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1af81e7c5f24100d246364b2aeec1be65bffb057941426b5743d9f4a34453408ddbbce193;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19558bb1d03f6bc68b4f19388eadd54f1b48b0d2538a26a67aeba090810c26dca768ea5e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ff13fa1758ffd23568a64c11bcf483c17b37505603e79d81b5d9d18bbbce97e0d988d2d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f8603e86ec006ee7a25fa057fb3b84bdf646ec565a7f9fe7d805b09ac623cc3a8a9e4ae2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ff67585150c5ffadd95313919879496c912774071d63561a722372eb6b33e6454837ce7d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc5677db5e4737ef1b9742f6e7e15f58addb5ec31a83561b4596dbee7308d15aa7dd1196b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h925660f5676644c36fcd996429b4a9ec87938e88808c484be342c86402d67f5625279b52;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he9c0037e16b1026188935f662d036bceab0713bfd306b6facc3b3763052374417662b698;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cd68b573d4865cdd57c93dbca20ebe61773f8551085b4c4dfe2f8ecc84fd4f4cc5f92dc1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15b258cd5e113d62eef64633b8c2590704beacc9d726afc62b87983f44658ceda19fef3b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15d015f1cf4adcdea316be019fed2004fce7a5c22ed37f95f7fcd691274c0080819ab45bf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5432aa4f208461aeaf4fcde897a1cef2e922bf5fd1cbb72765be7192ae0c75bcf64e10d8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d664bbda3f52969e47814fed96e1982841d464858f2cd15808c706f1b6186f768b7a4c2e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfb3f0a161dd5e4de721c42c54f306163d5b93f6efd93733e6f78944d794d4827cafb6eb9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc2edf4f35d85c6e3693832b08145b28389fc5a536813a9efe22c4be5989f380d4f57d5a8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h158ec145d97858cd2665c58be1ea53ad12752fbf7a611e68c7d80bcc618e306eba9765820;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18bdaf49e817c7903f2dab974e87bede7226a632977f774121670014af4d411cdaf7073c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8ca8680921822418eee3dce80125adc94e96410cf6d3b2b72d953a73f629477f44d5337d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha663317847a5df46c5d1bccc48cef664bb722a820fef66bc7d600df4c08707bb507c8738;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c53cad84940ffd6cc5875555cede0c744fda4cd634f7a3c3868af644163ed614ed25ec26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hadb06eaa8411b303662aad8ddd589b9ba175cf5034485f13e8725762bec206cf0766f98c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h133d3f6c3ed185e8211dada0d3b9ff5476dcf7622ea4d397ace2a780d52a5720447d22cb1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h51058f41b2df726a4b14080dbaa768afdff41e1cd2b4fb0e6e8d671e3c058531ecfaecca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4a05cead24c84a56d60fd5647fbcbd0eef030b8262f229f54a56ce048758f2fcdfa3c16e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1832cc2226c5120308586d6452a2252c60288c0c5be3848f0a60324f9cbeafb992b1d410b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h136eed1ad434236c763c5ffa842d59b4278c49902ccc0ad1ca97add5314452fe94ed03fe3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9316f893d322f09cfef87658083106a3e0c740c479e5b2a1888092324dd502d8b2151ce4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16e2c787c2818b6274c5f9addf1787d1bf603bfdfb83e8065b5c9366a81de3f0c1a84ae2e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d2057d0d74659cb5f95e98b0ddc8032d3d60a16371d663677b4ff46853ced87187764b63;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha80e4e5a9b1bf6ecbf5b9e30e0f651ec0b2841e95a0032335c9ef0f363aad0889820b3f0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c887a8fb4749d5392b12806149294a65c404934c1fb08966890d31d9d946721a0c9c59df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d82892cbbe8ad8c2a8b60ecd05edb59b8dd7197beea1da99bc6cb109920ab2f4e7a97566;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h861884c2ab74e2ff6340f1fce2f42e76ec26a48fc3a48fb77f392b7fad2c8948c42fbc43;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f36931327e02226be5df8a6bd46da9f45a78947a2695acadc6afff6f66e8300272ebafdb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1229d9237fa99b8585a90a12703e419ae6c201773b1cbac21ef3da632b83d81fda7bd45ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a3d3179ba4e337c8e39697ec8fad54654cc50f3a583c3e9847721afbffdf6b00a13af3e5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ae838155c60712fe471c16c6c7b6328cf0d64dfc22003a1758157606b79f5e0910b38e6d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h75af052eee0c3cda0d1794ff7d414c3ed25c541136890d2fef2ca1506ecc04115a987a0f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8094c5d44d2afd979c198e247d29039cc1f4d6e0d5aeab08be1b31fe7ee7fbbd46c1415d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hca52807efa29ef2e0b9caa3ca0dc22d0c9a5d5f8288e1aab5747be2ab97248e14e7eb992;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h48e76ee8652aa6ad2924dfcea4072d898a0bea73226fa1b33556faad340927a42a6dd7ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6abb0550a2605b6a3a7a4ceb4c6a8d0efcdd8acfd778660586fc5aa13780c4f9505cd363;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17376f248b9e16a18c2367fba9d42a0944feb93cc9673f7419fc17c02c4a4e63fbab328ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fb6eeb19440e9ff12bb881c49fc23676d4a5e5133e151c636754bb45640b0547200a7848;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcc73cdb6077d999ef5fe7217fb9ab718f7e1ad2b5979c8c5d5d6058edc891f5ab69e6a2c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14632e4648a27c89f7b12e3fb4bd5d6196df0f73d03069c142f8eeb1db4a5ac2c733922fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fc224bfad4e818346402c816f67dd515e3812f252af11fa56931e008e10b0c1d6bab62d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdf8d6a1528ac8f4dfc9ab817a094777d55f159508c905253bbcf216ae7feabd89619614d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12878bec382d2c8c9b2c007815d3cdd95c2dab76ebf58251e44360c41fb7e82ecc1b4baa3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h86ed673cfcefec6bc78afaec961465c7eea7a58f9db83021eb567280f2e297743f764ecb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17f0a7458d98cbda7413d7c2aa9e0aedc046fae7de128d5d61afcfc54a6a69f223cccd790;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16e7285ba8bf2ac1d6618f3e39f065237fc23b8a6e5fd7480295ead8f08eaef0b91a8cd9f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16c743394b741035bd79308a959a87a8316c36fd55841f885b1d8eab3414da23ad6914a82;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha305cbcce1e9717a59fc0a25982ae129c2c3c461aae6c31cfd9393fb61b14b4b5939b5f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h33b6695025c850e8208a1f91412651711eb3c3cce5d31ecabb5b046c4dc54e56f94559ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbf221e9740d7c7748ea626250136967156fd467b5f81536dca83c8411ff9a8f2e127e7f1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hca945e7996f2dce8ea91ee0f0d10f3dff3eb02c0a4f74171fc8bd2e9ac4d26fac2b3e1a8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h64f484e67d9f16808414e539c4bda24244287da305b6c39794e8aef8e6a6b2180ed4bb05;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15b209996f48e26d68e0cb25a69ce15d7bfb6efde033c6b4793bd7e4ea168468c6ccc69a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h632b60adb80cd8e3ff4a53a84e19cbd6f2f11193de932cd6f694cd1990b8773154e78a3f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13238596db3a67c49ce2e4eca4df9cf55e46551da0940e01158365fc6f3fa01ddcd86d1d4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1329f86d5d360faa3e45660d645a4db7acc7628985c3f0e6dab25a626e27a573cb515c86b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3934d3d466b90bd556065a708f5dd8401929497d221fa84714c3cc78c622d2aa53ec62c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d0d2f08b1a13460b577e45d6a60abdba0614a0887be2839eb76309f820c86388d6fb5c7d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha2a8056b83a1bea7fd9c460d28145c11ca3cc67a7347fc7e2b71d30bd40a3ba784def0fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1866fbc97296b8871967fe9d451643722531080e126bbb74bbde57c333fc9d5a03fed1f8a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h145a880761523095133516ed39a16d0c47b1dc6bab8708d7fb81690228d326f402f12aa4f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hafac1eb98f1e48e1a771a47323539c2c3377930a3b8eb3b43eab2ce2a8927e87fd2d8634;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h807168d2098bec4294583e3781babef10a0247d92a03aab75495d7b3858426182ab66e43;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5df426d4bc5774f4ca05567b2b08165f32053cca6970a8f07b70f08496fe579c7940cc7d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hded0ea355404c2bca4f440aa100830ba4a3728c1e25b92bb25cff5b365d0989623668d8c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1478d69ddac353575b162f94bfcf637e363b4a673ed4cadc46a8d48c121c6defdd49321d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f95fdaa7a43a3a807bc300ec3df03954943d0bc456c5af07939bdcf8ab7d27832b9339c3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14cc8a01e5d9b79f8c5b83a7417cdcf58761aa53d63eea23dde5d7f1cb89b799cebc39792;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc2e3554f360a527c1aa0da7a0af6a3b797803eea5f4a234aa50874bd1049c7725cfa5202;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h179637dde5f21fafc27e4beeaa8aac9bc822d853e4efe44d9e9f8273dea285f5f02d2a33e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h111836f85fb5fa0098af6db794268495c732865f6a5ba7e969b28130f2f89a56e66804d4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1abdd32bcb999286bd38f201f1789f81c3a0675972c33d1c9b23127a77f64251ef01e0134;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h65a229fd5b5593b6dfdeb651e48b8aae3d3638632c3469d8a606c83061e1d930805091cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h666f177190bff07ac34494faf403d1225875241300e5cb469b7245557c3065560079dab0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18f4de1e69f5bdf489a6415137f548ed132a20a6ad8159fcd8f401313dd7fc37bc699a293;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19250c8b51b63322ac2ecf45ac824a6a05b76d2f1d6c83765649ecc1b0f013726ea7e8853;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1700976e3765a266686621142175ffaf36c3b7c01e176ed24f48aa2220b727d01df9108d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h152e4fab86146777363434446cf162f2c60e6e30dd22322c4c6e719174bd9bf13af4fa3e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc508213ffc2c40186c66a4cc681788bbfac8c773e0f15c45f7acf69e9a054b2785e8e4d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d50975324fc9e821e5d83f364f9be793d210b0163061ca9cce932bf974c3f9a951dd7535;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb0585ca5e58934ea02c00589507937f1419902d44fd61bae4fa56817a163b70fbd29918b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3180b17004c8f1789b006b99b651f4ab0e3ef6cc5c8885ffedc47e8f2c36d1e72056b935;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3fcc886ee8925d0cec4b8e7db41ea395a07a3ebf239d2a6a8647e483004c0b1e43569234;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1508ed6cf82ee4236c2a10af97cdc1aeb494cc24d093a63fb39f30797d17e8fd491a3c6c7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc31c3d2a3e9704e32211b5ecc49ebc289d064fd6c23ec6392771c4e694db5e18fc1b0d0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec3e2183bb4c60780c03d165c0b1ba7c669ab46b84cdccacd803f34e67d64dd54df7aa9e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aa6c78184fc22a5d2ccb1df582293ee9335b0a779cfce0acb4dc68a8a91ad79155f21bbd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d860ec36669aeda9e2a701ff5e50c2b78b5edd04aee6ff2531dcba6636868cdeefccb22f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h181dbb246b274d4483ac0455dfd54bdcc82ec792c26cc6f49cf7527aaae4bbeb917be52c0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19afa62d111736c921b5263d8d247e9edc4553bb77292407c78ae73ba6a7a4be9d1960e9f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haf33baa1d132b766fb3c87a46bf82c50daf62d167f877d27eb4ed6e550a1abd799f6eaae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13454add893b2d306f956c4e9415efb68beb078e67b5687aa4d8b2e43b1b28b7fd42fcba3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb5c318a43766e8fdc13c84fd85c372ca4f1fa38379c955fd3879aefd96d9bc4b0d2379c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1110a00ef459bddea80c155aacbd6216aa13e3416fb417bbf10ce1ebd15432656ac720e04;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h93b8700bac1014f3d835b4d78b68c9d7528d18606db515a20a33c7df4923a889c92cfb5a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f3bb0c0965f6eacffc693bf3c593072e13fd99fa0f8cf49c1ff94091dc67230e5a4c782b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h37ae1da988aea93ece5280a1c82ec71567d92ec1c6b363b2e2eb578495bca54e1026033f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b5826953bcd13ea451f11943731f8c973f30261a02e2612e9218258f5305ea367db0b7b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h850a732915b20fd4e1a6a6d8e5b172520d08c2feba0a9dedfa179340fed0d7faec1cf282;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f5b73590d27bb45b20358304aa8cd7d181af0840e79d71002917778f3fe4ea3975d4872c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10b4c9e4d0de45b38604854ff1a53e0e1d4b77146ec1a321a588737cae819baad53a7c29c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h56636d08e4502cc06b4bc2c0a66fd633f33cfd69cc081600c5840e3fa2c12c9e89f3ce53;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h137b56bfc6a347bbfc54ca882dc0a0d47441bf586d38dbccdbdfe35752d17abf62379861a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5a87cd045e4b59157f78e0cac8166a82e0a1d2a746628897940bde8738ccdb588c93f72a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h945c912b857b69bc0a456bafec40407035304e3fc7ceaa77fd2d8750989af738bc38c120;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf67e6846e1feafc8794a6dd4fe6363b32ef1d27e42b1d6c8ac4575a7520ed41a424812db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h165aedb5e85bb98079b13c0e331491b2b4c90962c0dc76ffe246134d2a3dacc0bb4747f96;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h157bb2864237c909ff434448b2127a14e3fd4c14a309979392fc5dc529d821ed7d92288fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6c90a3068cd1d334f5856a131e5ef417c9b870c29c83264681698e62a0ff83e0189318a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16e3b9e321a9fb07ec3305e8c4f37badb6dbf85dd25ba1f1522069f5e75d3d5f8bc621eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h121546a833743938f3011fc3e26c01f7848b6a3f85b1fc134632d885b85fa5076e6a667b4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c92aa83ddd41b06ca5afcea77708bbac7de51169b04dafab0fd516a9708b449a473730ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d2438647503a2c792be76c9240cfb8d657e1eaf0efc4489c724790c4abd00fbabbe90a19;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18fabe07e3c9c2c696c1c82076b3a179719b44cd88a96c010d322966c34449da5c817d215;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12941143560077d6edde83a5a8c614fb1670a5930d6e0893753a982ffb5cf22702367899e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h97b63964af82a42660d68687b2964d9394085b835e9591ec913d025cd40e0ced42f3194c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f4780fa6e355f26dd108722e605e267552f74a4e5c7ef8039e889ca047104b8755cc89cf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h31d8b5e94894d6122dbcdec61e5afb0ab021bab28d1ddb4f42988de0240edb16b2af65a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b37b96b2afae7bb0ce94171bc7dd254ad36f9b1be350847e9b5a3e2371e501b7c719667a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17f53729cbef39c7f8aa5dee28d4000ee81a93e7d25ed1f55bccebbf448248cf6ef0a07e3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h524bee0be82958ea98795352aee0852eb3c75feebe605fe989365ad99bc93350d3ae2d5a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h632b1bfcfec992c3f3584f713c0c7496c59bc60a3a80d31b5b99b37ec9272fc18058635;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbc9c1f3b0223dd4baefd35196bfbf374938af50e59990528be9710d9d667741dc4d5726e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a484bc0242b6805038c6b1249b8a9b001f1792c80590f7971cbca1e6424bf1766d1e66d7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a7ca246dd4c0371afa030200abf2f29f2aafe01939daf16f1f5b5c1bc166e92210ff079e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2b2bbe096c26aa6bdc2c36047e297c7355b6971b768d79aa30ebcd5a52a8a18a3db464f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haf976e7d4ef3abf45959ec4f080b4cea875f1e7795a93656aea7963994923950802cb164;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd210af48dc77e849a4edc48796dc7a1ea60ebe2c306e9261dae7535275bbcab5049f436d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he461379aee7b37f63d10044616c5ed7e58bb735d5d979f1cb41d4d4b951a4887c38e488d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c9f838d1d38a719e25d79a7336dc024b47342e9740e94f2b246c508d9851c500494ab844;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h107c6c017ebfe0c28cce26fe1539e2af3c1cb6fc30a55a7227f246499738e0904785edd18;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h897b936f62653308a279a2c6a71adccd60f1a01595a6959512d9fc327f57dadd9046623;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1743e8072a55f6c2f1882ed662b58e553c5826a9bd5a06fb95239755de84d83996913a720;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hef5460c3cafe391453b37595916c49b53d0eb2b1c03e24c4603032d12850eec23d4e5f23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h61c5da666ec7037128edbf56d8e991ef83bf0b01bc129881413f7bbce0844a8ef7aaa32e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e4dbf09c018aca2bfdd9daf8dafaa599f5e20acfc517f1c0676d847f8dd178c95edeb1ef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcb51a42f6b2976e66a862b717c227bf381726c0ce1f2ffb167f5f2430e83944bcf9a28c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc8b60f11ac92dfc9ecadb4784f21ae44585d5f0195e43e596787cbb83d700d0fc3677d9e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8798893df3d88602c771ea439e1065776d7358de0740eb5d76b7e1b513baaab4eb9d68a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hea1b9dfe06321dd7c78b971ee3288ff16114cdd846c556cb5ea53a8f77ecec8c04dfdb5b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17c9b2ad51295e750b8e414eb43d463b320ffbc8c0e7310347b66644faeeefce32a1f18f8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11883507510e7bd285fbc67001911691db3c388fe37717a749a721bf1531a8ede3fcb51;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a85588545e8452984e296767e2dec7271aeb944afe0a1b998be8f94239101c46b675497b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a0f695c5e70f158b24a328996bedcbf4645d09c8db5a44a0ab436d7ec710bfd14006aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he90a39d132db3d0bb9052791b357786bae32ec3f3a6db49385043ff8ace0003874ba1c28;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2290a15631dace5b61b8605e1bbd291f7540669677ab22b8c377bf0afac635a3644e3de2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h62eed1bd055caf454bdf2a3cfee44c89b9ff1568fc30a2af3972180633a0076ef1c40876;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6024480df2d5035bdbd225be0f538415863f678d56b037ebfdf0ee878b653a4cb8fc6d13;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3497bebffc2fe10fffae9219f4fe6244c97976589706973b06cddced4fc1e08f652320b1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf93054f6ff7c465602f6a3a3f14fc688e3d1f548ef5426a2b38de1d2f87cca50ed4842c6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h198e95544b27c3e3b3edc7f50eb3c3894c01aef9c75ac51359fbcb13ccd4ba6b2ae6f9dc7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h115d153fb51431d64b403179c36255a3c1a81db31d0c506fbb52418debcef2420173f5e4e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h397dcfd27c182d26d106af7700eeb7eaeeb2e79b838dacd7b0fcb8569a09c49064f1b31a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b46908572ccca73be105f856840aa9f98a8fbb38bad517a4e889565ca96e67746769271;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16f0cccb67427e686f64695bf9a3ecbd25df30b6665459a582bde4b961c5e8fb4448396e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdd8f063f9dd0c96be5516bc4398815f748cf5e8e44db5552c5c8f8fd623566e81fc8dd8a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd84bb8a4cad9d995e778c5431f4b59356f469bdc1d616f6c540aab8f04791f97e56a25d9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ef50b0bacacbc643aa96522c0c5b1acc3676fea1234489dc1908f6a97ccb7100ef666f21;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha0ffc68a84401ed17722eb430f2810c90773d9d0e3df32786c8a6bdaea5bd1d8aa33c3bf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e49733c82fa92c21af92c7631567374c39f393ac79f379056fdd7155dc6daedae3c4e89b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h109431b8031af10e7af2e8a8676e37fa2d0c76fcfda7a226468af69c977337fe5ab2466a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10402a4b6a479a271ea60b72874bad56837fbe68a2618c15c29651f6316228ddd82a4b66c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h465d40deb7792d5fb36c7cdf7291eda35a930222dedb8c7236ed942f6ecab2c10eb896f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b69aa8796672eb07607a83c2f68ccddbeadf54d814540d25078a54b20f00eda74d094b26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3f64a7879d04ec1cfc5d4110863075b2df976a9920ea9eaeaa46a8bb0e06779025d8c76a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb69760cf114ef4a78ab9da15a171257061ebc6f2c31f1c35b90e25b7fcc468563094c326;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18e2057465ef2e87250a3d47b379d0f33e0e043ee224567119f9529b9cc163f69e272694;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hecc45b6aed8b538f8206f9c2d5bc490242830c843299559a70bdd18ead7764d36e7f0f31;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h32c19451c1efd0e4efea2ac627334833bdb89443c2459cc6603c0f1303357526f094de1e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16c8325a2392c8319fe6c65470b8475aae680a819bb28e8a18d06bcb7da9c273d603d407d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h127f59dc6b78466eba8b6c4932763ef37bc04c8d0ab01bd2d389dcb6e239e4fb5aeedca0c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc5568a9053828a3980042c9fb9c32027e3c4b5bf49bc69ec7f03ddeea914ae36bd657254;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5f11b3bc6195094eb5f35f4130baf4aa8431922d3041077282d4b224d73cf6c12c1fc64b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f6847091e86cc8c3e834be71db19367131322efca6463120320c58bb54e61d0dff9fedad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16761d95c5cc69b62a845f9b421cb9d58bdd1e9f298b853d78b43cedb1b89f3043b0a2e93;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4e69abfacc49ce4db1b9c50f1237c15fa465f188c2a7b713f3f22f15199ffd09cb4d89;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dff03e0a1371ae099e9b6050340175ef873ea0e4ec55874e905c8772ab621cb5e031f67;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1663dfd3a400e4d634511f8babb8d683a1a44e1a1a9189ce0495caccfa7908754940e520d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8dc8323f70de3b784604f594ecf45174dc27a39e635c7871bc45c84c80e541650ab38dad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcf22b0e99e2407efa97421977851a8a6531be151bd562ea85eda94d8bf4968be64e3fdd5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a32f28f7bcd65e2e06a0fe5df80f8510adbda8f8c188b59b985643d9c804262e49e795c1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc38edfbcb2c0151cbce031654ff5068067802a90f33ba54473399510fa5dd31b8d2f6357;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h183967cfef6ca2b72239808e47fe6aab236bcac702aeb9d81ec482453ad58be584ec29b25;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hccef9dc4d19d8b474f959625076bb5804173d6e9cd70e503363f94dd35ea2101baf309c0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1262f5a4e7cf142ab9dc6c4c43b4e385e5a463fd8d9a67902fbb4903c51a772d4951cefc4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10bdf41a2dc187611116787e113ade856cd47dc70e567c7e6a879831c0ae1db6b3ef67216;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a6c2b0b1a35e208b682a20c9be7c7e8c1a0c87447a6b19b2e3540ade8b4c339ee29066b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hebdbb529d81389ba61b3267752fe2d031bb5b399d6c0ee4538b762b372c520f79cac147b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10d88e5c7f0d3cf3f0298a1840f6cc451c6f9f22de2e7382c35d128b216cc53b7f6afa8c5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he20af4d7edd92c6356682a60df046de445cbe2d8850006abeca7076268e1fdb2b6c6512f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf71f329ad8d9ff1aa007d4434fd144f84e269bb57efd24389d639deec69abed65d8a03ea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfbd0724b17e827b0b679a5b5aab6628e284450cc178eef9e35fba9c6a4a58f8d0d9ca00d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13cb5a1491c767a2a6d67d57d08e89881533cb0695c6fa9384c706b556fbfeaa0414781c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb83f520d2d7c89897e5a224c065f1e7214dadc8d1a93b099de4c3e0bfbf22d1443638c3f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hda81b645e8408662b4037e74a8e5732e40d25f893091c8feed62bacb981e83d249af008b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17b5dd679832c292d9c5b394d9b7be9c75ce981accf1db27c91ef0b9c21e52d3e005771a6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h185bcda64bc168f3312d498cce7851ccf8e11f170467ea2a0c94ef9da9749e18ffc4584d4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2cf0bb99781121af6e314d01f76783347d5fec6bf7518f105055b9bb4ac76f42d1ec72f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h36f72c47f951dff08dadb72d2e7c6c9334c492a3e1280bf7727247757a0b3dfaf8dd4f44;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h85945abb4f5d8417a4a097b2e6ae95e671fc9594d7acb7b174fbe3ceac88603d1eed9834;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16b194bb468f2dd097df53ccaf44c71ec7461ea52b94084a369f99c1748f1118ee94f51a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bc80b329d0d3102cd5fdce27e10fea87e17d0244f48670c2d977d3adafc4a2dd2b547e85;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbb694d048c8a537ac4be65ab97c1a2129e9f5519b40187522ebd46bff46d3f1b401fe76a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he5f440db728264a23230183469c35adc99bf30a42ae01022639552e8ee934d4d8af11d35;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1786dae95a49c1a07a397c84abaf3a54405c2614c80d4779d4487a67d687056778f67c352;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10cb04e4b9ba67d41a3a9cd661b67e113bfb04d706729ff073a3ab47f4fa07d092ef28077;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9825aec1af5b03eee3b1be5ecb98e2c756b5c6c42ba7e786dc268503a0f844402df054b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha651428e71422574ae36dd91ad55a83cf952d41c578db7b6d06c8d94f0ffe9b25f384a46;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd39fcae49d5fea12f7913a8136ed26aab1387b45ae685a52ccc0b10a4402eeef3ae9afb5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h107ec3af23f6b06ad9c6dcc7d6e727d3789f250c26a8d7efff5abb8d269e43b4d690de06a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3e79fdc8fd7e24dbe2e3a0958e7d418327951edfcdca08e885552862cb7251d7ad7b1150;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcbb7b547538405c00cd588f5da6ec1227e0cf37c9a52b8680ae36e62f0b4f4127be8fb11;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb87c4c783602f09dc49f475a9162bdd421caaaeafb3875545647fc8f1949c7e0fa07279d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c4a1df397602e6eeaba746b08774fa56c525632e67354c71cf37a4ae072929fb8a73b58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haa7e504fa53ae3e22ac82792695c93b69d312ef83f51c6b95584898880763063e16ae5b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb9d5a410c0f8e60ad68135d8bc829242d89bda6d8064a7427e4745bb3006d68670d36842;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dd6f27a224b290fa81968fa48e74467af3aa22f145ccc84e1365712f38cd13725dd05cb2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h188a1d9f2edae2c7a70671a8a65d61dea61d2d08a41bdf44f38c0b1df8b8cbe1419d52ba0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17cb5a345c0a2dc3351ee5b9e6b66b1d1249d8040af29669f66dc441037f0eb8c760c0a63;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c454ffdcc3533fd02d009e1a7975c6374b8be4de8dd35b25576aa0c18f748370afe72c87;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14a5528325abae9547748406594c8991fb6ef36ff931a8ad83ee9e2a0f23b11dd5b46d6dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5a4de075e343f1c7630f984867b235f09a45168f3c99cff52ab32108693fe5eb510d2d11;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17de8b8c66c2e3101088c64da02d2bdef57d71d0b18a5bc6889e36e5f0a1ae3290bd8b631;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2d5eb10087860a52f677a2dae8ddf1b540b18b48031da5176ffd01472fa65b26809d4ba5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15f53ede3f0a928f8cf8c4ba64147a2377cf8e46544ed7db00601a925e2318778e937be85;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha9f2ecb05bd9eb06c463dab9e8c5b55587295b8886c8b8c498b8f86184c32faceffb76c5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d47444cbd3fa722b71219fd1d0e0d89dbc2f1d9727f89398efa9f617804d6a30771b9a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hafa24903381d3390397e63363bde203bce9fd8aece722207d130eb504d4ceee1a584ab51;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aa25b19bcc304a1e1212505e91716340c4a6306b2d705808127e7c7bc330f1c4e59fcfd2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eeaec924c47a64c8b30096bc576aa1853a7bfcf29961808eb4af524f4d7a4a15f02dc831;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h49eb20bd8ba051b91b96c12a1d2124b2dad7bf8b63d6a188e774c4af3f06c350c974a430;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15f61443a12f4f5e0ef4b53f0c4a1a6308627598eff438fcaf237ef90fbc7cffe6641fac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hba70b03794de98f6ad1dea9a33205ba56160d02f64f78bda6914838175a31833d9aa8c0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h162bd2bd829d7db3073b7a493e089851dc182265ba0efab977acfc6cf3bf07b90eafdaa13;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbefce684df730fedbde1e58c0d0aeaa3dd73f30baa22bcfad67be41faef9bb3560486623;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h105363fc310c28184824b03dcbe17b4151f3de1552a205abb2f69b7bee0ef3ff7b9e098f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h90ae356c2c564c062a7b61c6bfc92a5c825502f8704ed5fa971e6a9589f4f43afe5e1e01;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1de5b4b9c8562e39858dbe3d8a7c8770b346c61c93300fd2e7dc0485767afc5bb361d3269;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h117892df296894870643057ac6d36184181f1e1daff0681d58a6e000847fae6b690dd7c65;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16246a30fb2eb66765f3ac0637eabcedb3b2fb72d6f97035953eefbe2fd2f112446a029e2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d68a93776c9aedfcbe89ece72a7a491ebe9af629911382ff3f82cb0b57e79989ef2c2884;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h171921a8f268b482393b5c8ea3d9b06cdfe437718f394f480ebea1480df6dd922b944850e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d83637732e10d3e2cac44efe90b5a83c80a6da2a06ef288f0f8eb7ad31841b7ae7aede10;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18e888fca9ccbc7e227ea2317963f348cd347868c51ffef484832c6807a91db7075e12e5e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1130f9ce1af28860a31c06e25bdd2043c4388f2e843ff8824367ee6e97aa61c9fb56dce53;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c263a4a3dc1dd904c36f7a63e006e74d3e309de87ffacd57f6b10ea05f2ad6f76d1e8ef4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16772c4828105d6f8eb52b76ce9de7eccf2828b7b6c2c074258872f98c77f5d6631bdfe8b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cff791a9d7053e9c875d32d9914624aa9457bb3ff285382c3b5dde1ec7d4de6495a93f12;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h27347d955daaea5e24a652592e955ee88bf4f04ec1236d013169ddfb7e892b17279c8388;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h264889c58e1d3359844b74347416b38baa9d7e87681dfe6f5610e47d445d753a14a12fc3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h144fc873a8df3d0206a35bd6d11dc29cd334fa196c51800e2ab14e612640935c153ad0630;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b987f1a7c9fe07b3d787d574b2d09caeb9a8424063479f431c29c5fbd5b2e8b2420ce672;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc84d60e9de0505eb88ea9c7d6feac0e205a7606aa6da86157eb98732ea2dc988cc48df2d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eeb37af9bfa5761c706e8353a3f213077a6d69be062d6df1f54c50951bc7f06699f4036;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d35cedc699c6d99a1720cf6a31674bfa2d427f4884c48cdcc8e72ef0fea83b334f1dcf9b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a0fe4207a8c6920cc371bc7039630f154d14f75cef1449b56f8216f382fa1e5c4b1ec90f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11fca7dca94e0c6bbbca16e5d952aba104a3a0e5135a2f6df66342c04afa1f8039ed88383;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11a984f57e84bb38232e24d5166408acea7c085eacceae6d12b44ce836e0e4d4be7b163ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1035c7f54f4d6c786b40bfcb139ca9db40942bc4f2e6c60e7aefeebf1772736229a6557b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1804997c7abfc31972a03d7cb5f10da5c4db623384bf31d85425be3e9e352d5a4361ba890;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9dedc188b53f4b6f9c25250fc3cc360d43d8c39b032d0a67714d248e62ebd249b6ba5053;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4eddc0051e3207cf7f9195922343e14cfd72b6bdc61f37969bf6ba8cf4057d21499ef30a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3f366ead3ce7a5529021d2542bf38be34e8e255d515bb6bcdb71d8df0f0d407346c91e4f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b8920fecc8ac3b9cc3c2c6f622b50a213f5859f79c55c097baedf7190d1c74fa20110fad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6a59f21047f5c0e004a607ef0745a2756a9b3f75f6705a106d68025f0b299bd4bd8dc3a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19e6b561180487c0a52fa4033a3b2b17a1e2e1c8723e65fd7780dcfc4ef421358c16038f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h29860c293ddfff4c7d3c2ddf5bc3093320ffa7d14f2f853dbbf9f25a4cc225fb4d1443ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e7772f3e277394982e7eaad66ee8fa69db75bd70cf5967bec4db164e914b09104e05b0f1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h141f5a50d0fe6df38add75e72cd7a48b9135833c34528b96ca18dc6a9f84c1f9e2b752344;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb92fdc87d648012cef66e7f3f3f521c1331d25bf662b33df32a10552eeb99f5a81e72b51;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1613e3434d9ac74f766b0115b22083b41102c38160ca65c22355c32e497883df9cd6abd9a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h71d596315d08df2ac9bfcbc031fcf2a003ce333883dceef47297c800e2348a434c89e22f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha3da882882238b2a505bab12e7cddeaf94aa2205d2949b74b4faedad28d646b15c4a43d3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f6e76afe92debbffc86459531bda7aa3bfec0358e9395f6246c2c43661c5926ecd1c821;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h489a4c69c7369b73df066186e64df5a929d2403fe20366bac129144e340b5aed0e31605a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hda1f988f2ceb8be0fc64a08d204b8637660624006025e0fd2cba7641557f7bb884021e88;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb25a45e0b689347f5997e27e32339bca5628b78317a4990a8d642b14cd954f692de3b1d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6ffdce603b7eb6058a4a7edd3c63efb8acab69e3e09a528363b226ea3de27276ce8ae3cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he9b4b01b250ed4fc5f8a7f01c63d818e788ad08ed9c40a9573f0a9c69a01bcb5db6fe56c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc2cb012588e6a9f19332d773906c3f99e0a9409c39ba5cd20b7fad9fc51d865ca665682a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h537433b73da14989f7bf79283a1f1f49d060d9a03c37badc766f5f93a65955ccaa00d25c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ebfba237a7e78eda145740356aab59c18e729a158b6474322b1fb23c029fe2ef5bf3b5b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h147c4690cd667f303fc2859c746dd439f0363600376cfda6bc9b125f9be2d0c6cd5e817cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h168586f0b754660f8a2cf48c773c5de66ba337796585eb4f7373f644865c41a71472f839e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb8f8a0fb2dbc369c68f48fb04495ff30580c9e49820f22636fbe5327db2b627bf04e6b66;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4a79fe2a811374b9b8e3be0f9b27ec5da81d35dee29b3ada81180cb93c8df0f506245393;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h105e826fa4a69217b0559562075a742d04cf799c310bc287b4cb92990b8318f8eace8330f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9acd544aba06ed31dc4f48b901a58e6f31e38645d8c5bf9d5f00805310372d6b5912cda;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6a0a783c83ba654ca640a4c273ff72e81beed72cde6f7862f2029573f732557d7c975810;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd9fc941b9a0a1971f9f54bab438ca731f9450941fdd5534016c9715db3cfe1e81114caab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5aacf0ff160940b41beae62d1c798fbcedf5b66d17ebf126caf552599689e75556550190;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf0aa8048613f4bd6904b4994d197134c32cf72ce5381dc875376333c3db0ac3e9c1feaba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc1e853d12d22a37d3316593da97f656535fd227065528a00b6b97f68c7e45e6e42eb6639;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb9a0078e629ed8eded348262cd9ffe949d1ec829fba056ac6cb5e73ff04d5af8ff12caf7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8febf16e1fae1040ea2ba22a7afcdec90f03991c60a4b8054ee83e343c8bd024363bca48;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12fc9031dcfd277410bb404b556faf4b3d8559df8b0c58d0d058dc423726968ccde64bf75;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12253db89b667761c78abdd282aa2b088d261783127d265ba260f62bbba66b354e13b631f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd9e6d5efda91f9d36c79aad8669dd7ac10bd178c7a2bb981d9eae42fd7e168eb9c92c11f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h184a685a5dc8995c0d1f64654ae9e16d23106f981c777eb13eb7c955a10b49df7c6b7c924;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1794b51e6844cb31968ebd198eb4056f1e6a083905ac92f2f1d11e3b6f3a8d365ac332b1a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fffe82f7b586312a3602de507e1f6605dd680d4b67dada7ef45161bc7e65ba791c129442;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbe4bc8101a029e76eeb92cdad726aec0824df70925655a403d748e6182d98477e64ef5e9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haf938855e6387de215669e62545c810596b3e3facc4640978ef708964f9a79d983cbb4d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5a497e34ae35f28ba5ab6299a91026f6ca3bf7cde67d7faa01f710093dc8e62cc72b0e09;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h154aad47883568de68e4802c57e1f7881c0501d87521b7be88fcb0d2ed21410b20ff06978;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd614a23f94fed7172b6f66d8e57678cbae52ce0875c194f23b2c39644801a9f5d1c09a0e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14283d43b17423ee3a73f5bf191a3522217fd004166f915128676ae3347ee9da8315a4489;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd00d75891b524f7954ed2edffebf8ac617f919f2da33a336808e7bdc4fad614a5a8863dd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19d988d2b4949c67e3eafaac1e66399089f6166f14b57e10a13a7e8da49dac1ff4732967c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c34c915746eefb258456abee08eb389283e356b76adbf036597178ef0460b4d88ba0ac1a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3bc65bd3e0da9635e0ec08d38544c1556a3fb5d47a4e751936765be75325707d990a973c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10954797a51d815c1f41e496af23c39fca26c44d1fcaa1171978d64d013ef694204dba352;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h547248cc77ee6ef79d74f25f3b436a624cee25379037ef85d27d7a8ce423cb0209cd954;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b6d404a19694148332798c5fd24da76c3f324ecd0a30a9160a6b69a8cc63e51ff174621f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8be44b13b0de1a4fc5d1cdbfe6682d576e6a50d86deb90ad823d0d8a97e9f52d49fa59;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1193cd402b739ca0bb115c4d8b535de31b6172fe0ab024184e592e563496c3d302e774d73;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h151d3843bbbc3f82435d75ae597f521bed897799bafc1e86b0b08cd19d5c92aa3280dbd3f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eafdbf5f7d75a381d83631603450873f515e3499a47ae382d1bc17e49f9ac2bcf4db9e6b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h221d615c5fdb97182ce7cd175e8974ca1b123726e60d97fd29fa3fc14e08ee4fc220dea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bf28b15ea2339333e3a9e1d1e1c6ef0b0470bc86c39fe4ebc6e32bd5063d468333d48a8d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6b8e678e58300ba04d873b897dd8faa06d6c1fc5a719237cd96608b61e070de145f3d03c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1266baeb243e2900d1bab3cf725035ebbad63df4e20241502d21bd76e506274126ec44bbc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc7da6257bcf9873f3da18621bc17e978144967851e48eb17ccd86156ac0abdb52b7f5b58;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19db7d8d5b78a065c854b43c955f41f6095b78ca1022d92cb4c27aa07d5a65169df7e41df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eda9ad0f84d4b58ef3840d838b21ba38bfe41d69f5f145508dade8701add10710b5a7361;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eabb363b167f358523099b61d084415f62b5368bdb433c85196744588bb6ef22a3b06ff4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18930221210133d1c92f687abaa19bf3d5b55ea83b7ae1ade279bd50644587ad6084245e0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3146f9f78dd661a7adad3618744686b375f7a6d841782607a5123c5611fd2e9ceb9d3ee6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h198c6a41a5cb1b8c624f623cfed52047713cf184fbd9862badee7874ce207ac19c4468c9c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd3b3fc72c7b91dfe3054e32105db49ee0630c03189060f6cb8796963ac4cd37769f2853d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h977cb43ce161dfc6e526778ed368d498a693ae7c05556897b672f489e6007718208acfff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1da4e9ccad95fdbcbb5f3aa0603549c5a22c9444db8eec5f331f2c5eeef09942e9c2ddbca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h110504acdfa1c0fafec24f87466330a5e466a98b4514987735abf96245f5fb384d9b8b297;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h124f35687e43e0bc3c0285d03247a8181a942eb7c250faad3ca4016a15f67f68fd9d3dc7e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2cdb64fee1dbdc9830cbd491432d62cef4eac01863918267d7c7f5e92fc0bacf95c9358c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a098241d2f2d41962c3f8e5a281b1a66b4544d9b609059dd32d170a4457860c4eab6f12a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11d704761080055ddabb358f990906eabfb1c5a56a931dc0a7e938b1a850e8feaba627557;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e750b392590eb1e7e1025e582a95471fd2b0483bdacefa26ea7daec023758e2d3aeb0fd9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dbaa563a6cf66e648bc80efc677aab04ba22be9d406dcf85f2373025baa484d9fd131be8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c65b3dad0ef76d6e12f5a25dec7bcc62d4a77a981bc74eb72b91da61db304e16249272a7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc47d45601b588731652efacc82ed938f6aee157dd59dc7bacb7179c2e3289b207cac8903;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h85ca7000cd30369b386acca4c41709826c5df47122cee9a6adf38e7129b62d3d2bf0a295;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12cbb6dfdf98fde129b92b32109a8c808b33aca6571ca50d85610985fecb9f36f12c5b01;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e4abdc0f4c3e027f88d827d0f0a56f697d8f383c471ba91d2f46d25e8f3b8fd718c385db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3b31b9704f9686ead2f70fc6719fb5817b764b1493e87fc2c0c445bd670fc1673342cee2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8022d80d631075fa7027d370201ed85bd269c6dd8b833075c5659bb0fa4098b064673b07;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h90a228360c0d6709ba94b7dafb7758c2140f8e77068b53fab83b5dae5c863442b41b3168;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3a841746c556239819e35047554a30b503b08a2a6239d0be456fefd8d7e0f8d7d4d7800;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15bef51338bd3b0442b9a3279edc96e91c488c0bff06ff436a882f6f477f05a362dfe87bf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf27419850cc883bb3bde8af5faf19aefd1b36fbe0d7361ab18cc9a6190f01a2260a23147;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11e585bc1e16719c167423f47b76c7cf1e3d94bb67830e063401e147cca89c0144f9f8232;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h26b11dfbdfd3cef2146905e77cce5a93a24499e9388f15603af0abafef137c77802b9b90;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1644d49ef63ea42f8d1e15949b672fda3492fad7f3fad6d07ec4876c1f9a15615dc20dfc5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e1fea2e336c5802a3ef152da6861e56b7db2b5ffafb77c571bcc07d54d41ba0129ad2975;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3d18b0dd36cc845b7bbdfe2e29986e03daa9c5b4ea1458efaebfe47f765584655f4e17ea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h185df8f728a4d3a539bd59800a77e4813a40f2ca5ae7a4f1d338f3b02e11b3bcc78840cdd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hea3898afd1b98a71293d25de2acf4925efb68ca7256f87f09c1eda7b98179f84c0946e5e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb7e2e44be26c823fa17e3f0b02cf5556f5c4d5d238970c405d0b17008f3616db5f79643e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16dda4082610f54ede6675e5015f8236abe89fa65dfe814361dce95fef2e3599acd021c89;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h23eca5b3b004cf0b13cbb471aff6e6dd66c0f19e4be929fe04d578091a8aa52429831931;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cd74e328bdaf100a6e223fc942e6fa56235aa6d8c5eff95a5396dde829e77ef36a0d7aef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfbe7316e354e492c9cb5524f986668f462f6213d15925418456c7123f738edae5052a8c7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f90041dbc501e1ea65e1a3c15e819fd22a64fa37d156c4a3e36709302acd72dea99edc4e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he2de8e83a81faff7d3bea793ff3acbf13a98d730afa0336b3bffdf50dae9025ffb926086;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hed034765bf3fa063f78532601de1d38cb23c209a8c7435fba60ed82628648f4e3c84685f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h94bc5c48dfacbf2ccbd4492473a397e939b2f1b803f556f97d2b7a29835eb08ae0093b42;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15b0b8e96a38a27c972e6270517c5cc69cebab284161bdfc74f67a9939abea0b87d2f2fa0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fdb6d2ab5420a0a9559be4b47a48c57755c682ad84c8dcd2e36765bf48bbcbede08dca27;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfb12c18f45c18c52e68661c1c8a06237d8ff2922424460709d7e03f2f9a4af9bee0c8137;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbaa706c316bfc2901fb265ef5dead57dc67159eaac70815f059c26ef1dbb2f2ba6c00570;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b659bc224828fb863f151c846df6fdc23ba94dafca3ca467961705f30171dacee9625dd7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h24a7a3b9b4ebec795aa432a09f2f0639b867eca0e940ec27512533ce990774e52ebbe67d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1313448a5b50b181cab5ab122ed0be1f5f65cd89a010f54ba91433f251cf48acf02ea3f71;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h125a7a74c29709bcc42ddcf8f33b9836324a29374d6111db0791dbb4651835e04267f3b57;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18967a0aadcfdb2214bf2fdb8deb629e4ce3baf513a382cbfb30a2750ce9578d922a7acf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17833ff31b1d1f5af5fa5433522413f8a19eb72c81970f6053958bfba2a3e7269f35d737f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2a0a12ddea10a7c1a7c485f05b19a2cbe03a21bc21fdf5004c4170e59837ff29e15a575;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c8d72f69d0b786dfc5622c30f4f72abd73cac47e0c5cbefee273a1395aef6c5963247dd5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h107c0bac1e6c7e1d6090aa2c5549fae1a55544c92e0726a7f7802d1d2dd7cd9996d60e584;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a65a700244abe5405f71d382fb877d64ff30a434e792253c68309ce94a8a8401a927a167;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6acda43978ff7f0c8a9a7374931607f6dfcd0fbe97a737b098b0c1c76b6f23563a694a43;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1acc3d4afd555785adbbe30031020d2efeceff29b2352777b01b216954799a2e74841b20;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ab0c5f1fa7e2f9a587da57062f97c13b4ab0a845ddef87132b72a3b145ca90c1d89a6810;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a487e905a203dd70df351560c2454f2645490b80cf7ef433a00344e5ac0587251d32324f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f6e20081c1fa3805d567f51693cc2af54510686b44238b934d7faf002d71c833d3b90fce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h380d92b655ceeb226949b93190f7cb2273aa2d034edfc588ad688e9bfe3e50c82b83b634;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbd0182990b268b1c940b9ba5c6f94454bb1d3bd9d6b4e5f9820b239a830d2b87bff8dad6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h97b27383ff11f43980351d3c289a87dbbae9c34318fedaa7cc8661941d3ea172cc51478f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19c7942311175d4b3c2b728e515f63c503b80d269047c667a30243579f2e518e90558e439;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b89fc00128d47718945a3dd8ff8e26f0e8fadd663c9e06d75f6e4f4344816a7dfa3b95;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b3a99c54b2b986b825b5c3a97fac90a836a0bc9d1eb5b705c806f9a5308b1ea03d2420a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12d24c6abd11ababe9c827e99be75898cc3dabeb482965c3b8254989605860400ccb08c9a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bce728829f3fca9f33829938786fbefaa50fad19729e9250202825613355fe8acf4f87c9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h89250a915b3c2141deea6498044788766057602d9d8cfbaa2c557bb2c4d1cb7207cd0c55;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h22647014da2af0c487823341af6933f812496a17e477b8711e1fee2ad4a75bf76b6204be;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb3d7bf3ed03e0e6b1ab53424fabd3f2db620abaed956a25d22ee107a451d5a3f161efb9d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h148b4dda03213b2862f94f564de4e640ac85c2b42932ee9695fe7cf783689553d99220487;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f8f84560c0332645e4e6be2676b9dbc09656b14652519476d8fd9fa4470cc29ee887e483;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2b029c2a950c1676d2193d283377df1f3d863353ea91102d5768a37b9214bbe67bd3f7ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h241a145691f4ee02a9d51ca67e77aeaf75bf9fd89caa270fe143a0915da56225b53cd881;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15651a59cdada56b4169f0df2616573df66d68e8cc43e6a6e62ccddd5b46bbd5a62bbeea7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha79e646918020adece12dd58471c572fd2eec7280c07eae205de6a948fbffe1a2d9a025c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12b47a16e9267155c08769fc4a5b6723712a7f302ffe39f9e41089893f25ee332ba95f2e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h760bbd8bd5ce8379342b5a692bb378d4c83759104435229cff3951af1cb51b4ab2ab25e3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a6efdae1354ace30c9ca60f347d928d508667346f05193251d8ea1cc7f9d771c2a61726b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd05adbc63acb9dc844865dae7cdf00d666afc248d09e1afe88662abffce314a04c897a7a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1be90e8291a40a14cca41ca8e2aa4a6bb11ddffcfe3ff2ade7ac27df9248524b021ad7ca4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h195918ceda3aca82aff2a7643d1ce544156fa9195200534bd5fca1e638d22682fcbd6732d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h107c83a97f5edcea79705402c5d7e3650263241de3694bc7007f04e31fc3fb965ad28db4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f498d5854ec6e873078c1e4f76dd20376bca933d31c38049fd5e139be1a4c7706d9fa1e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e47a6bc5893b96582a0d491e0862b02543ca2f65a8ae023f708f5a5027a098190c1d5b67;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h66c882d0804988cb445fdfdd519b6f5d53be836b1958fb823e1bd8b8647fc6960c6bfa48;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6f5115b42809d7f2050a604fb5b8769506ac569e2328bcafb300603ea853730dd9b206f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc84f5f38f94b4a4be7be29d34196b3045cb0e4848eb7b4dfa88bd3b6bb271bbb93445c99;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10469ead7f1cd1f4bb35efeacd5b393c284ca6e92cb3eedc9fe0b25bb90a7332b4918fb1f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb1f1eec3f3c00e06c08d0b6b3b4663caee2885fa9c28755f60c80515ce371806fcf77d2b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1b9c8efdf231d4536f3589676a235b43f46b46e5a51cbff3e5f72723761ea89d1e458b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h160efe34c0744f8f4ce91b27308aa54222f44689c9362aad352857a54b598da4cc47909b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fde913fe705ba176a4e824c7c167f6a7fad50568a55e40c63dbd156e2b9b4ba24aca6105;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1676a6dab7a6d823a773bd403f8b4eddf011a8adc25fceffe8a9e342acffbe462fb0a6aeb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1067ca2bda88549337d5913be659916a0130b0a709ce4a79a06a69a6227c8a8b27f8efd87;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dd40a7f85a74d174495a835408e230e2b8c5aacf5bf4d4a111e517d817f508cc31cf369f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbc05b873d6d63882324ea0ec749eb10bad35c8864c31de2f876c40ad1ff085936353bfcf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f666563942732105a22267a4e5c39fbe006b9f020d9ac4d472bccaa88363a0050789793a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6b9d19aaedbded77083808b642414e7e1153ad66ce041a96567e04cee70d396d481e72a6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fc0ea8edf6d0a79d1e1e56f76190a2f29870e0cac5c345c8a72645e3d72ea67ab46f829e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7dec5ba2b0a402071a27418aafdab067bce0a1a922cf62c9ec196e2eae23bb038a28fb18;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h776f0dc22fe3309544e7ede6d03e5f38640c844cdd823e7351adbacb54368beb328c5b34;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1950acfa56bfb1d773c7ccc6a30819eb02ae2fee27a0898d53ed4613c5aa86fa7f17e7bdc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc8230c9dc57f461b5f3a99e909980174b18feb9a410d479a9b10274c9da43ae8b026127;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha3e447d08022291bdb2f7ced25bb46030eec8def8cf91cdc6a7fd8faea57ff8ac25af0fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h356e7ee0126e8a324c49abd0b2ad0b6115d67a180c8cfd5b1d1c3a61dbaa21e360c177d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bbf4e98499fb432db6fdf5b28480e1a493f7e55bf990333e131eccc873616b69755da5bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12dde265cc37aef17350e9e0d2950f8f243e98d16a1d1334be9dff43af64ceae4ac4ed41f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1723cd21ca02aa0eb2bf9a4cc0073068dd3a46383ecbee9579a5a84b70af490e890b00656;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h34662854db03d12a0d372ff0a76414bc3084d07efe11a204bd5cf796217fe62a58f20cc4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13029bd683f2ecd739e289ecd612792bf926f2fc4204c89a2ead7ea3e532859959834f394;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5e494719c42136f06b2e1805177ace77b6a5b47429e0b99f9342397ecaac2c6692c0db61;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14c16e7e205674953b0c14470607f5aff4bd9b8b03608d3bddc8b96afcba4babd2e8b6794;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h910abf44c280bcfcf4485714d7aa550236bcb508f2c83b900697fb83c6357535fd4fb772;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ff0bc10f3a090d94be25c559b7fd260d8775550ab14a6362267e7bd82053720128fc767f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd076ac153187255326459fa8df419dbf12a95f5063338f5588c160cc90b3f2f0903d84b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc0804bd11bdb788b70c67b1aba2ccaf304314dd0de3f42296f4bc0384841ece400aa30e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d1623cb6fe5a693d889f8e2aa285897c2fd7e8e44fb8ebb1fd8188e6b6cc7e834df5f864;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6ce518d63b5fec3648805566863e1f737a6f33073d38fea47af5ad775abf2aba8d3189c8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8b97f2c58c45417aacb0219bfcd15d54bd33bc9c5a46fe7186e27206e1e534ca7af2b96f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cc1e396a74c1d41b41d1618a09ad93aae8ec4dae0c09769b60bb8491126a4b07ff07a7b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4037125cba5ce1e628bfa1d6563ec95fde932eaf6c650adf1c3a00af7cbb724013d60c83;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h484bc370ca3b54bbe123fb4f0a990b3a78f2ae8cbfd15bfa1da778f331a00625f0cbe2eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h133106228697ffcb85dd3e720cae72aa43c01963d9c9ac106f7dc88ab9b432097c7798a20;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11bd2ccaf109147cc18450ae0c9cea5243f6de87d8a067ffec4363956c4a349d1466c84ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1822ddaca9c31a8fec33d9cc8f09a7d92207458cc40ef6ca7693f0f8801cbeb5ce13f0574;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eda84e72a57e6f078ebccae2dea125caba779fbe3a3fd232c0dbf198ffb8b8546023a610;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha3f0a07ea4a9b5e8ea3bdaa04d9f1299d8dda331a96ff9983f5d206176e3535d3a0ab9db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3b0ab75b66f8fd4c8ff4d77d5b6bddc4f5852728d90fe89f77b0a8f9b5791bc92a90aff0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc2593e330b1b8c22132322cc997ed5b240c3ece8c4e9c14df582d3aebbc70357d3416ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h134d1827d11d34fd80d8c4ace8566785b92c5a030601abf67051474990c2d15d7fecdf633;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16ac47733fe9df3377d7020c0c598a36821f7af8176df5c930f89d192e17a8f78fd113238;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h208f0e6595ed4cf5ef4eafd003af0e7e7f64b6c096a8fa2c419b26cb098867d81b79fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18d640d01287b0ad04e0ef0fbdc147847d5e820f523eece2d2cd4c663027a7ab4e1581d0c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13f6f210be299a8c925500a1dd8bd40aaa9a99fdfec6e72f50d8a298617eafaf6ba0b52de;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17ab53bf8a32bead0b6ebecd95bf1edeb6b90034aa469d1e070fece424e879c4a2ca7097b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5cb02b729b597bcffce86f76bf7660ceea8e1320b3cb61e8b6363aff579cedec73ff757;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f785573300ac9a069c138f2baf1e1ecca2511d8fe67e5b65a9ed28ceee526ac7ae81a6dd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d49a73c89ed86be66204a484c47dfc5a8d66f16d72ed06f49586f45cbd328a5f57fd1568;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19cb5b73ee153dd27516ec9921536a827b6b8ecb99cb7621f96239f434d96e3f2833e9581;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1299bed938c614cdb7a91ebf07102902683987d31f6184aad0181ce80a713b2b948237300;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h216cdcc34ef863d1624fa0b139da3d4fff180f4c990da1c08e7f4c39f45531f5eff0457c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4cdf0df2f40985f278aecb762e4e30f4facbea687809674fe1a166a40a4a358089c54cdd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hebe097b5ef89348b5345468db0c7f81bd1db5be2f7679672a7882cbe5f3de0e86ee6f7e0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h166e597a6c9aa974f020a80bf7ddb4d86ce16bcd93d00e83c840413db6a7e19eadb66f64e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h62c36fa026d82ec201e9835aca71079c5dad13a48c90d601252ff1be61b2deb0fbf598a2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h69d67c3db3e8fb3c64f05f96da3a13aad11db39501aadc7611799b2655ec8ce447e57116;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10d6e67a4dd2a129026e435b05d892fbc556208295993fd7e2a7501aac9a71e9b3a3b4127;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h347848e19e47f0cb477af95b5b58b2a65fd8bc56608679088c92330f76b43160bccfc4ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15fc45f2518f0ab1f3af9f0720e6780730bdd819dd48c9f4fae133c891dbf044bd2fa42a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b62da4a87bad649ee3346450646cce3eb7b573c65ecd8fa5d94bcfb975564bedcf851c2c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a715a1f45c2239a4e51c154f0a07668468ed6c365ccad27d94bec86ce88c3518a590cad9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h108a83cbf7898877d610e1b1a667929033659219525fec7f4314b1f51db5a703606f654b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cdc5414ec1009618230ba15d6fc226289b7677662f470d2df1e29e1caf2eb08a50f9239b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a354ae7f6aa6d2339be720cf7b61dc9673720e3dedbd86bd63f39446eb6bea409967282f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e5f1f7aad23fa9c5335c4c2eb7d4b3cdb9f19fbecb55a9404f3bf214334a5ca03b5705db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15dcde81c91436c982b04e08d8b207daf6b57eddc060812a3bb130252c5786cc13b28d02d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f63b4ce8e322198c131ee7f2b7d9b239977d5e2d31262e8a3cb808332b040d35b9c3978;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc8ab1646d65b1f189b315bab097f36842e3cf80430001bec102c488a46a22abb4e5eb803;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h554e9e73d2d97931d7d12f3575c6eab21bad221c9eaff22c99bbc8da865a95a5710e6a6f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1347baec45837dc36c495792e1ccaea9a6b35c503e0cc0a7fc5c2333589ba951e4120c1ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1941121ff5f57a242ceb6a7706b30296de9d02b7872c6499d058808119959e495ed6f143d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h949b4c4eb6110f4be9ceb8215132c8e9f7a2179afe5063c3d5ea3066973c3c3027585070;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dadfd850671ccee3d8b13966282795a0727ba87c610bab88bd1f11589611099017d7f75e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1562dfffb178699759323621ab02a86d249e8e4662aea72eb0636887353390c12cf9d2f03;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hab75f77203759d29594108912681f2bed8fec4bfceb470d9e5e244500ca5a772235e0010;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13434fe325e1f390cadf64ae94c63e06f294078d02295f7ed88ddbc797b65f409269fb9bd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4abf0b107cc9e05625b61753d73f8ef97329ab7ae5e37a54d8fb66b0c158310dc3e2f4ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h604aa4ad6b0fe9b0d571893343285d7e9522c336e9024f1bc821566a9b9663a997d79c26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9b6dde9ad2e82984134b08e777e52ba06657bf026b385f8818c77da88ee8fac197b52c55;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf4ab920aa4effedf2ee4723c274453fb046778ea3f3111a40a08732f733a0c7eb1d34080;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1014d5109ef0b6f7f13e5baf97ae730b9251fba8ea6798852287e3c16114ec72171427826;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3f1f9e703cf8506e27ba17d1d2ede820a248178f929e7b2b85091a6164403b308b73af0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h152f68c524324d39f36ab177a460d6a21100f47de8f059aec4ce34f054664d94e202e698c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f41630b1c8ee9d4d82d74de8b49b20231d536bd7d204b8adbb1691fed57bec1a6aa3587c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11e0f81bcc5c8a25aa23561029f8dd9fcf265f13b023325e94b422318d189534ae901e56c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he9e4189e50e3d5fc19ab23f57d1f43cf1564a6948dfcf78d5eed939b031c65ceadd6fd7d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14c668225695470653cddf858883f77f19e0acf81ca4d31b08ee57ff8f6585db8b4670f0b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5efab8ab340bd0a2035bf33f4faa76d0a9c50aafaf81200ef42a587c87bb483a390a7369;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c670d08cfaf55b536ad241b5ad5701a2357b694653ff9429fff901fbacc8c61e98957f61;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfb4e7f0351e38da17aaf654f3df55cca194a7eb598624c00f6bd8210934438b0f0a462ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5d82970e4fe2dfefa1d5f5ecf3d4d3be73cf9664ad34000cbdaf0c3596f3b66ad762b2ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ceb6a9ef6354e381629a6823073be35fbfc010427bbd03159d727d4cf23788e6d813dca4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6be7a925c04e6998b3417a0b76e7235d7c1fd90efe922784e04ece6ad5703b06577310a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbbf6220ac4a8a9ffe9ef59c715dd075ea55104721dc5b32afeee3d67be18721adae81bf8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h114aaae04dbecfe1dc693979e2e9aa3a79f80e63c8fdd5c5c5e9500a13c9653863f36c303;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c9802784329a26242a6c67e05adec49f9d4510a0bc28ee6d1b966a21371c651a65caf263;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bfbfc7fc88d0ff7267f239acc80b82229c85629387fb947bfe93327ddfb1e6036b636bc9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h111ce9e0dbafbcadcb119c721aa0d29435e26e8474ecad4d9da593f61a7be2f5f0ef2220d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8aa27f47ebf02e57128930f4363626a28ac6a229666ab2c339997d9b4381f0f9f7ff34c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16f6b5f1f066de483cd1c71fe639571d1ce2ccf8e0cef11393bd3fd596fcd754d9e2baace;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h168e6362e6a03d5d0404572c81adc10f8db1b6cbeee70e571feb67dbe10d28994f045d054;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h156d3d941f78f261546c2fd9fe59d4304be1184f532a37ab7ede30cd4a8b8bac3bb1d3068;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3b31100275e780eed45e11c87fc89ab8da9d86af3dfb953163b20647b3f5d8fc3c9fd0d8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7a36e097d6e6a06a731c2104251022713c73fd083ca2fe36f546ad1b763ed652558c088a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha5074b81973128e2287a9e33ab3270dd46376911c24b18194d74ff7e32f3b320b2daffc1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f8287fbeade455bf8c2d5fbd9d1fcf8c8f05c118c271035553850d47757a1374378e6af3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ba9c101710545216231ac1811cbe72eb8a01fd7269fa751890a6473ce10fa12a094aa27f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15e1b1e720fe917791d255e1f18277a67180e3cb91e72b09cc6034c2fe19213003d0ddb53;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3cc843ba7fbbae502252f66d60c7a59e4c4c3c1f2410d6d0cdd4fdb49dc7eaedb297cd0f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1402b9a866883339c9f8fec5cd539c3030e0e212eaa567fc5a39124474e4f31edd6be5803;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1156e7274e846923f15c6daca9e9b38ec2d0579b3052e22b1d57eceaa2da81d7447b214e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h195192e1d8d470c0d643477de3fd22f5affe3a373f8a2d488805292942c9f951d11d3a850;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3a6e54dc6f3f3699c1ae225b2664d796e9c207ef58890c75769c4f557d56cebc2b96698;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5ff0b8d2056006e717b6167bb07c650297bf1c2e10cf103d9dcb2cf52141946039a0fcf6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c6c9f4b1d6d83d9551e86c5c734f62665266d7304c8b5d1032defc4e7798eefbbbe93c9c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8eeb8dae6a81d38dd6387dd415c4954270936471e566e961d78c3436a16feffbc68651db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ee378e4dc71b89c0ec5fcb791d3107bb5c01386f2f3668c98f7dc05b1c64bc04f0873e4e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he6abb00e3ba4649a6e512dcac23ab5154a40d03d5f60541705893018cb0684f0060eaae6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hee0657e0c34b36efe2c864f9f2ceeea9e9fcee8939585a02c205799b11f9ba6d33136397;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h124c5516eab3de8d2e2ab237ece174a49e0aa7d844bb0d05e0c23c5c5192f51517c6758d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b9a8f25f76ab7a1728d6cbc9f79bdf34452470b7c931f963cc364996c968a40e8fa7f8ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3de028c979f535f9fe0777f48b0a5a248698dbd67c6ca7c3be23ed1e912eb15b0d2a9f97;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f99c9db2ac612abfd107419a961b95cda373b9d0f67cac29e8e7244fe3d2ac250157bd40;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b01ad33940d5cac4a52820cc5e33d3664937f2026ddf463093cab1673b9dd7b3d87369ff;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11ed6b7c1687e2a24fe75bfa612fed673d656419c855961af915abb8165a822122c46c484;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha2495dee33659e364efa8e3695ed2d75d4939d31716d4db9546e70768cf2be5ef73fa5ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6631d27825618f7fa3bc6da2ba9fed45a57033faba583a63c87e44bb3bf14ff61dffacc7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4d591cdc1c164bc8d520a4a14f1317e8ee42d1b37d60171bb7c6dc6767e525427d00d391;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14fca0442973f5ea59677f17bf9b9fc88d0598d024cd5b7dbf98af1691e787893210472d3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcb2f2748bcda0ccc2e790a14bef19a887a7432e766aa0e1b563a8f7de678ead3ea6b376f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4cc58c85f857321d07bc11933619d7e572336c3481726025b1bb8990916d1e48e92b9905;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4019bff1c2a6c8018c0360062ba0065de7c7a5d5ee48e845761f8b9f92bf233a1cacafc1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc35e21f7ff692b37a6ddfa5ee6a8eccdb6a0571ace752836979306f092ab38584844cc28;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c4c9e734cd9d9c484b83a0ce2304985fabbe549980034adb9bb4607d1855e57314c6d9e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h98ce965b93053efb220031f304319129aa625961ada17972f8e12d0f0b46665257eb02a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf5260ecba360a1ea63f402dc78ec7ea98146549353c4d238b148ecd5b7b9a57735fba5e0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h363f00ffebf1fc89aa493461a08f8856c7b7cf39250e55d281c1f5da3a1dba0253eff86a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h85d4b61be2b56e95c9a696f83c6dcacae9812289f4dcaeb107c58afa92e8cf09a9b962b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd8b654ecd1ccc98585cd1c08b18e51b60880116a21f862b745dc3bcb5c1adfe36133fe4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cec542ff6b30a1586d2584e92daeb261aebf60772647366489f9f3058f48306a68dbe58a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc7a737fd513d0d6408f439c78e55821097e619fccc7f581b3e0181f41301945f8f6dcca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15e6f61de8bb0c13014d5b16e1f1683d79367079360a89db8fa401810b43069eb4548d271;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h840485b9876511efbf98c9960666959927e79ef77765650572aef30409f6970ee0920eb0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a22cb7a7acf8bf4c850b884a9e1e39670521444d0de45e7750f047a417d2450de7e2ab4a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7d12971b9748b058f3b0ac5fc79a3cd1a8a9106b667c0d9f6fa23462e37fe7e9a7878120;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfba97b8d69514935b7df7a3d2c92077cab1d96611c3ba4059bc81d1c93f4d739b3ebf2b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h700c8f3191adfa6dba9814209b031815a763d5a0d3c485430da7730256d63d50a5bd6f53;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dd2af7230f0c37b8819b3e32941b1439d5b8d65b9301bb283cbede44c8b8b0ba1c859795;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8469543b0064f2796830fcaee2cea775a72db49a2afe4772ef72cdb0b769f90d8da7ad17;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ce2b958c9e722a132eaf8358d737f709838afd0aba31a6a01c9ca6a0ec8da18bb07d4601;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h199597a9fc36db1af051e281ffb8f0943177d306fd2a86d2bd64f542f33dbed73b0b71f71;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d3cda041b4a521a992dccc79b67acc1266a24fbbe128ca54692446879589ee5fc3aec20a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h30ab6605902b034b764fe0b063eef2fe4ae9b823fce373a9e1d5d4bf736a00b3dc3ef975;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h137cfc2cc9b79caa5381fcc798539a1f05e5dcda5a378907b7c6d5c95d47e314f08e90678;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb7e3a3fe2533dcea40d638384b84447ff926e172790a2ad4ed9f72e5866eb8e5455dc7d5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h964c75cadb823c64028d2c347b24ff2319dbe034d8e41bc53ad8c8397430c4593122e33b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5a8304a9417bc836f7f252b2c16fbef5c7cbab08a78e0e8cc186781908da0469590cb5d3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1171de75dbf00dbceea9d5e8a69a0678988c5a6bd33d7b0daee81b34cf1d3a16589eb7860;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ef7ef36a88d588734067b56a82084f135d9a9d14bd335cf25a7f5f8f2c4aa696e0ca7047;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8dbadf16390ec4a1faecbc3a552bf6bffe654cbcfa302e91954d0ba164fd81d05781d5fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h175d283896bfaaf08fedcff1dd76ebcc23de845895e2c0f87c33ae7759920e5345642ed4a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha809d78394c8e192c788959ce67b19af0955dc089c1293c6ebb8bc98c7b67db8bb19de2b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c83e0dd131411ab032e4c35753949f7a709f3e6d8e383da10a1e3075ea9c4ff3b5a88121;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha287bfb36776ea498451747bfddf619b55252ac39b47f44bb5bc61cc6bc6270f6a4ca3f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7913060a711ef56ed1d2903a151ddd7edd78aecc1b84f403a60fb80859154f98d65ff030;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h151e70ab50f84b01568dedbe401eacac4d53b9e8a18050622616085525d8d92576b859ff0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12cc3b72ffc6b18685aabac8e298df000110fc32bf9e9c5ca3e5f51699840079088895638;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d6979230a1e6944632998b767a4f2eccb53dd1f7dd89adb7b91ca601df4720ec82f4362a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h155e5a61f00ab690afefcfe0e9b42483eb102b59cbe95ff67bfc520646475084879dde427;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13a3e52eb42fff111ace4fc3045cc21b174abf348b8b72dd9b285d758199ff4b5ee60fbd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hda10a5c36caae9f21c469f886de329b0f7f1a779fee72ad455259c391ffd42ee4ec8e6f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1922ccca032fc2455e95f0c2f17c3be296a715bc53a079519bf8253aab9fca3f27962a148;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hea7bf1299ea0d2c64c74cc81ff472f470dc96fa9916f87af328dca3d54b234ad64526608;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb9c3599e9928c0b489dd9dec1a7f488ae079233e5d09b83a5ff74f942c0f67a715ee16ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a3a1539fe9a897609b3c70b2d81b86407eec4f5a99206964e77ad94b1a4d7c1e99eb24b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7389069fb400f75fcea904fd9700d6d04a11cdd487b16ea104ec7fb328ed20eff5e53881;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he1123404317c3f042cd351393197fdb614a1cb2f6f8ec41ea02eb20877eb9585c392c0cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16c776ad7761ff91e5cf2d1572d20b546c9f98ec9a65ac84cb1d1907967f742597c4a3fb6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h42e0221f7e837fe3b2c05df93ce6011549a9a735400a8207bf22e1fbf8bdd35d66fb82ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6d004d60c9abf41f51f0ec76c4e92495c96df7d98fef6bb24e5748cf0f8f3138af46544d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbcd6810e3360437763de7393db3c60768b59da2e6b655c5f781bab364b1893a734bbdb1b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he179b0f896258c6d59c98f9e3592bcfae56b65a9aa6086eba87971202eccea841654a07a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6c521c0c46d8987227eba79247a6241c6b1756e49581dfb6023d1580478d823911d5d8ea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h196448ace55e742f7a397955cb52c9b6ff9f3631c584cdd458c0462b5dd5fe5a8316be75d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ee82e0f7b1186fea747705ade3ace6d74ad0d9d4394ff2c55cc883aae58fbd28ecf7684e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9d2ab350f4f2ce50a373520d0f49d1fd79a29ca077bda095df31762bf76cd1c908f8bfed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2510085dc1c88416fd5520cb5f4f3f43709e0fe52d4d16d673083cba6845b6895bee9a11;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dc1b988b4bb70ec1d36ccdc021a898e59f6f90620a8340fbe3a05d1c37e10e50b39a08e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha91690668c01f0f5f5f0fcd7df63b5ef6c23e713e3d4d45c42ed058b234c4178395a5acb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10cfe6a7f1d2dd5fa6b70f1c54285798a597f328dbeae6a47020b198a71cb75d8b9ac2c1a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf078f21ae930e9be56350a1b369c51796eec12f36ce2b13f51d9c43e06835d333f358717;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4f34f72d36a054cbec06ccc884d528c13c150abf1c28fa6182d55ead1ba22ba7542c4036;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h36b785dc80e607cf1deb0c7bbbf7d55d6fee6307d01a65c24da7538415ccd689645ea9ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7f5e0939f693f6d49d6de4a35496b47f180cde174ffeddc7377c870a712e09c5dd69e0d8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h65bc984ed205eab9d83871038f26004842ac0f8faf2d0f40a727ca9ee4e4b2bf125ed451;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c961333034ab016332a5233c82f07b01ac268e7b0ef7c0cf0e5194b0860491e32a76f05f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h450bcdc40378c35f504593150b20992bb75bfd824ac645624a75c1c2979e71df13c6f23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1844887e9476c803a07944822515ea1f153527cb57c8d30cfea9397422348be8419aa2c3c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h190848b46ac5c98bc9fe71a2984e3bd04e05f7075e814dea81b4b3809f693b6638c4c1760;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ec85416d53128469a0d53d7c9ba3c09a74b919e57de5ce8e8e5635994fb28612776e879c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10bb6ecd47e38d76bff492e115e8b530122bdedcad08c8702bffd0342d51df28ae9665c84;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h110e1293f083c8cf74e3fb05405cb8872977608ca4e448a4a3e5fe04603f2f40ddd99411e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c69a19a03bc8b79170481daea73cf161a8c849168fc01acf50b682f13ca205ec47b43183;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18b3fb8f9ef01ddff8abe7ff50c8568f372e2c3e0c5f49bf45aaac26929d7621fc991a4b3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h117d4c7a4d6a8f788fed8f5d3a45d05d260be5d85b760e6e45be79cd9b9433a2701674955;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12d148ed5eb6090386b3b4a60b04ac18ab3486b4f5ce2472856b8d574f254130edd28949d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17d86b95df98846e1f58add6f2f4973dec326635c0cabcba0c482abcb9122feb67a3b6fad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h617f29f4e5fb9d3e106e75477add5e9a3b8ef272e3eaa78da2e09b0d5627011a67b99cc4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h81838d362b2e8ff07081610e45da86317006f487df81d044ac159675604e1d496888e516;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb20857d8ae57066a6ef4f9ee9661328a2394eb749d025e770336dd7b84f3308b7e639a2b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15cc7ddbd9dc4a243276c90aada229c761bf8dd3ae0853b13fd61510a25b381d29a0b9560;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4aa3f7c1389577a8bc1042ede936023822feabc16ef8a2b6c59a6543e3bdc1c925990260;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19af3d7d638e0d20ca08fe86ac28cb0c88b55ad2e4516ae9f0cb5d2bae2738eb487636051;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h137a9d2d747c3ba977015a3706bea5cb0bd68b195a9f7feb872d4feffac622289b9a3884f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3beb4803c2bdbda4f4e7b34b3ef60e337d18fbb3c884a531f400fa29fc44f82286ce16a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19330c7af753879275a5632b6830e8ac3fc2b608cef30707da27a978aca5f2f8fa9f41708;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf46f23aea0f483adfeac2f56fe34234bd9dbedf690aaa59b52c6975fdf6bafebac605177;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbee24e683ec7c07afb4e1da4da759ebf82d39c301d0efd2217b357dd02a888227525a90b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18c8d7be0eb439dab11ddc0dee93e45ccc05fed93800e2d1b9a0cdbeb638fc28052286349;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h400ea37a3a6eb179fadf8a544ac5bc78adbc5842685f91d906b363b091e1e8128ceca817;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b97fe4cf9152288a834ebd9090b7fb4b88d9b16fedb2e9eee57590492aa6e39a58ed79f8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb69b640ef20f46bdfb4e0df93a71474c0ae92cdfd5aaeb84aa10398fffc47736b7e1a553;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16a6568d4d9cde5da639f3b5624a25d42cbfcecdc3660f35c03fbf691dc37de05dc4b1666;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc49d0b926d3a80e73fb0930912cd6af103d75adc87b4c768f6642d9f8e50cf4a801d4f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc561b487c6dfa6ced50bce5fd1d174150b153b53feb16ea3730398531b8ffaea3aba052f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfaa20b72f314d9a32f239ce611d7baeadc541ae8e295b278892f6700b7a538bf37cf4aae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13a2e94481bb9aecee4b2c66d10d7853b81278ad1c2866785cd9a340ceab4bad5e45dd6f8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d9d52863645dd72ff631156acc815ffa40ecd7807964895fd74a1df9407fdab7bc231d82;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h192bf4ada418eb6fd692656bec180d1a25f3ba708e7b6eeadccacd8409814708c2e7a501f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h107c2b0d15f2086bf5f0f7bca0ff4cf239ecac368617749e4964514924049d21427ee28d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h136b7bd1bdbcf2b6548e3fc4c472362df02863dc4637053eb67cb43d619f7951054dd3174;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2e78ce9907ace8012fd8e956551208fff939a9a52a3bd7c7d5f5156dc75b32dfdb3c7748;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h342094567c930f94f5db9197a9767c8abed250026bcfe01491739073bc2fcbc6589900ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fd46e0bc57ece4bda65695b336b6b09693ae1694faaca376e45864b75d232bbae38c696e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bda341034690bfa57f3e7c53e5b80661e2cc7e36a1176fba2ae5d6b1e28cc965005610a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c3a7d555733fec8754e84bfe5e666a79773d781ff5b192a9e95ce9535731ca2899c1124e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18e059656b2feea32e0b8d3a48ec865c0b63a4660cdf25667703ebb006a10f2b2cd8804ad;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4cb4f4e1c551877a200d01fb3d3df98816645eaf641634ede8023d1282670153eb085819;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1eeeca74b5d86e4a3b31c5a7bf3644a9a3ada2a636e64ab97fd94046db1b0723f217e12c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc67d041e99a4263f992795046534dd977bd35a628bbb255da3633914e5c52c6f9b876011;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h136f474fe4a81aacbe3469532e963da14947c2bcee2f774cab2f9f971a3efcb18847c3684;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf453d241834ebf1e5c03b5bb76983444499dccfe2ec12c0d35e6a14640c80166b5a13754;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e89a280f8c1af2a3eb3b2d04a408c832cc66c62ae2fd9e175aaac81b2cb86d694dc139d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fb0507e47ae660714a1c75cf770fa1adb7a588a4d4a6484d36e01d8f4525cb9f6e7975a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17b8aa745d49eaece019b433f8eb236227682b5fd80683e150eeef5f3f62d6906a725cd83;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h892ec834cfd03fca4df19b2e9222a6cb1c9e782a5f9cdcb2b3800f8106d62a5849e1a547;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h153c97541272df4f4c1b983240d1fe6b399e6703ca0a1d74e1e0649aaa5080f3cc26d4be0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10fb8d9abf73972cb19f452cdb1dabdbeaf286abb6a6213c14812a370f24e7ce22cb54115;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f8d5fa39ae19216b1e0e27544aa03793e86fedf8c23a2185b00082324e6cd23bf6d9e509;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aad3e0ebb0794da2e6ff2fee2234a01440fd436a94360151bb7f343ba9d3dd5c8d0fb33d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8941b9b1c9631aae5307b454276240c6121c616ba7cc040828e183f83b777181e5bd5a77;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12ec750d6a0e2389b99c9f2929db198a69ae44096332e31e1e72ffa98cc8a1c3ec6248abd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h39df10b795ea1bf40d07980731e65ca15dc855c4b297bcce99a66b39d3d30adb88ba7d11;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e716bdbbb12af90c95fb76c7a5d409a4070f03290d5a06eae03ed73a80509264472498a6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8009205b657c3cdee07d7d01685a0f133a85002fd859f73249cd4e88238aa7bfbb3d118d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fa8d8bc986794f33677116c2f777c09c246abd677f578a53cb89ec4a81973e0c1a5550c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h405354e8a8ede135270ae60193698d1005c75950078f5188589078268e843a7613e5c910;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17aa8c695415678b31c5b9263c62b80c072a64cab4e8c35c6d0e99c20cb2c6059329736dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13e1a192a02652d864cc2bb4dff70b24bd6280f173e1a2c0e80db12057a6c812ce2ecdfd4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h122493bd3a4d4bc5b47a59cec30acbbaa9a43e08d4938b527f9c76440951717971660ab54;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c56c31858f283b7ecaf2129da21bea7280fef21fac7e177ed9391e6772ead96a488318a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc51964d2d667dcb7d8b1c48173e0b9c8aa247444d90c40377268eb6edfa1e6e1296b8fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d6742cd6de92d0a7d76c4c0a70e528704a67d2d82c39ed55d22088c7f4f0f63768e7b0e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd0baf7f7eab7bf40a7841d2ba289bd116814944a7ef59b2156377ffebf30fd06ac267dee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h146e2dd347b6a07e3c98107423193422fb5e0652cc23ded93d60563912b5d8610e945c71e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h726704d2fe5a7b5075a986cf062b3a4aea7321b8400cd60bd5a6b619271e2d2a7b90e4f8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14ea161c8cf58e2fb7d2c9a0125f89901f9b279c79c688619e826b6035dde759e2bd28ee1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ed491d4ca7f4f53b489da1d394dd2f876d5ce62b2b627978346ffbcf2ad66129cf23c863;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8f5abe3114a47666cacb71cbb1fbb55a9fda9e652ce65b17a4102f05e0f57e8086a12280;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h156b44cda5cb0503ea3205c22f6be622e85d7fe3f43e8eabfefed9323083e651623dda13c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd00b53924b2d2869e0229665a8c5715f2ce9b9bde4e6127f6a28478ca352aa1fcf475a3d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h80ebe972e29d10d5236e601c2f07f353aa61ff3908cfa8b8d54cd9030ddcd4a329f52d56;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b6a0ad402c1f47ee5b7504c11a0219c87cddfe7f569eaf9c407b0a81e13b0641223794d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h112c1ad584a7ecd8735a7a0a2748c696b851f544cb35d847fbcdb484b68045337bc413f36;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h165d444008d234df5f3593782b513984e3a886d9b0ad9d6af0a38ab53c2d65276a406a813;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h691c1524c2414a14b22756c02eb23193128f9b089d7c59a4853e6086daedece2925ef7bb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3ced0cb2b5ab4a7bf97db6502cdd7d1260ea20842b640b381a5bc52e7266a4e0c295da5e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a3fe5fe052b57a533e24bd3ec6a68070682e90d6cb1dbdeed75acd00b18dba91a5d463ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h97e02b60729da6f79388e66f61fb735db66bd27394b92b3b936aeb9af415967049da01dd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10a888bce3a8861de53b2bb62b175016f8a69cdc36708e935981b361a9ea337a0f44c82b6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha82d53698e57ae91b6d6a92a775478c4d3cfb3821b40db19f421795da5d56b8bcaf4f2a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf8cfe64b4c3d60811ff5fdbcedf3189d3c01a65e06b9495ded52069932b7c411c3518775;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hab66a5dd012cf43fe7382797824fec61d43e01059eb5333fa512385acea1ae1ac6a18457;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cf7a004ebb7e5363108c24b65d88374cd83056002cd9515ca3982bc7670a7363ca2a6638;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d08e35f4bdd9b99f89292e7263e45855f7856e39dfe152564633f1f25b91707be9c033b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h177f3300c1fe99f4ca629a88b5035ec06d73d1d2a60c267f85bd8faf738a4137c57740d3f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9073bd622e758b01f89667b8c0160a981fec0a90edf4e6b614315cf296dcd3460055fa5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h304abb0bb15b3326866276306f24cb37d9103b248ebed34734290ddb6d1990a1e51363b5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16561306446c5776fa2eee3c6fce5e420601be17822c9f60a4d9fd17cbef8825e3d326d05;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf63a356b3b42cf1a0456420d614f0228bae5c09ddef15bef0bf0736f47fde40ad078db59;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d4522a84dac4efea8ab3a5e6835a33eacc7c1c9268afa1bc53bf1eff4de8b3fd664348b1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f25996a0d11985dc5d4c79d05996c910e5203dca4e5b64a4a3605b16a3e7d44cfe9be2ea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h177c8cd1689073b12550f98fe86dbc0d4e349c5b61b0f2be04b83cc09ffb852acb601baa1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12e857da123e00af0d2ababa357dc384e4b80d9495b83c8f559756eaa9a936a4f7620277c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hde8ad215ace3df348ad28bbf8284785ba72197b6d15110783f0cd5501b762f99ad0b5ba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h375005c61165c558263e9cda000de0e0e5a11d10d48cebd5c8cfe5cb6b22902e95e22e23;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1020aec3af7531f81123f095949fba16184d987e46701e8f864f8711f31fc441f050b3aeb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1846d01a9c0e6a1aa3938173bf56ca1c3609bb239b9d254cf3aa3202e5df142dc6703d81c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h967d58788a20aec7150348b2fea3f14f7a6961f23a5a40737ef72fc25125518ea920d389;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hec7fbdb44e2f692147c1add915c3a98c50392b851eb5c6ce70fcb55a301375fa4058dd3f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h35407cf3ed640dc7df8152b7f29e3670d83a52d1eb6eb8b45e37c2cc1d1ac258144ec56c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9faa9c94379c69fdb14ca6dbc02a2039e3a21933e449ca51982044346ca06c49132a45da;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h42471ee4c53873b6ed83e5186588d6fcfc371453bbd986fbe7f843ea5080b73039f1c90a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h125954f63334a2b941040380040d187309fc288121a86bb00f84d0dd122b393852530ef2b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16b03f75ba38b5132e3936114e023dd4b55f1558356d1189a839f121bf6acb972d98e30cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h57cfe875d4877b5dd1f10493cdea679142b1be158fb61741770243c675ffb4bbfb77f175;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8477446227119a448775feedea25a695eb9c1497073ef9c63688a48e1f7bd5f3d61d0133;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h182730792dfa4dbb9e3593f293fdb618c29f8a82ae6a19c0f36cc1c7df847eb7f3d4e3ce3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6d7cf0f3c64d182c3d1f1599acd4db0e1a3a3ff44f8062e6499427c6a266f03e89377736;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15bf0ba93c39c68016bac01efaa8a30ab752a455074d364bb3460948f96f00efa8673e27e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1515b5300405597e4fba97a45e2643f8cd6ef9a271c7876b88f74521cd2a91e3c26a75ba3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3c062ea88579dfb67c249879ebc2097063ebb29b38df2f2c95f11df89a3c4acb0c4fddfd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h71f24f9505300dda66b4b9693c07c8f4101a1882694250175321470a7f790f7dd7c94133;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c7a11d6ad753d5b639e8ec50784ca3439febfbde133697a1ec19ec0b24706c38d974aa5f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha2c15f4da6fba153bbaa32188d1754fedf4c04bed6312a084f262dade491ee742fdea0e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he449d1c81a369666c75d4785d6713f4ae738352cad9929e0ccf1d8b1d8da7124e2ec0204;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h145da75be096ce2f9467b38dad33e7ec5feeac51cf0e5d35cd9a248bdab8b90c1217c23dd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h59a77447264214e34daedfac48fa6d141f366c30d72379289faefa1ebeda86d64b25c852;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc0a8136f4997fa8f9d154363fdb218cebb81c3e08b4dd8a95add66bfdfc2cf551bca3951;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7fdba7f430d5618553c2f2a4c63224a224b2a43880dedf132852fba02b8b6e41f743a165;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1680314e8573f79009269eba3cf9e4d68a0c21da6c8aee37c374fe1095ed387f584db3036;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h45c696b3088f244f244b3c52d70f9c28a5fcca02238dcac1663379b58b4c3312b702e15b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdc3acb679248632b64f9ae20f12e0ffc31fe062ffdcdabdb2d9e01d09494e5f17c3c91ac;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15e9af5a5bbacf1dc3de4a3f1dc83f35b2cc3d2f6c0c6476b4aa0bf0f7d169ac2720f803;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h21831cce333953a35dd9ff02d8670012a86e2f904e5739b22c6c431b17ebc0f3953ac4a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb27d4185522a03525f6c49109495e6f67f713bc5601ee97e175b10b3d1c7a95b536dc9a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a76e16a86e7d386ae908e74572e1e6116d446534977c5631b9bc55d6fb72ea1b05d5e5c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12ecfff40d069fe9e7fa732a007ff8ac22500a3f052a0ef0f7c8ca52bbe0a49a5317c9eeb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e20f558ac6cc1b4edbbdb185b5951976c4b952af8994b6044fc72358881d0ba6b709a3b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ab43ca6f1831d5530e0f12c25e8c5ec22312f3d3af7a7df63e43cf32c2dd6d2741ccea9c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h181bf971da19054c0d2ab34653e3055d0fc8d9e8282edd4b1506b09bcb2b06d0a8e821888;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbb846f30fcf96b99a3ce72a65f2e14aeada5ab787efaefa9690ce3c7c1ef027e7724ff09;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c0c274daddf2ef36e6bc4bcfdc4e9c2436a62cea4f16dfdf057f5b0d93d04f80beb1e38c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16f6f6cb16b1a8aba81c3e0a6cc9a4d9c6d4df53b7cde8d389d15f82288592889ba991109;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8fa326de91dc8d7bb06dc02a2be2c293b3ff2d9c6481719fd442b738575280215e807a4d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb88ebda519ff213329fccfbb0d37c33aea8feba319f0d5ea047a1b43edb99466c3029aa7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a5527f43806bc4b72fd046e08f23d910d52da6ca6bebeec45b755c21ef3f5d7197391606;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2bd9c8252deb03a3374c313f2ca0ca081375d9a78fe668b1e3b61a2b70314a8121c8a479;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9fc6ab316aacc91b6f2f3bd1e7d3e1e21247404d9d33ee7bad56ce271117c7b71ca87263;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h182351de37f09bbb24bf6950c33911176e582563081c99281626848bec592e33ace6ae741;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h157dc617723ec6baaa26575929763083967209adccc7da18311d89c6cf12c2bde678fae27;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3cb305944cde812e764567dc2a3d41d21329cfeb17d5f7653a76695417c3956c69d5f13c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3679848b29747205d5c9e9e39742b208e709cfa2bfaf7d2a947457de06d29de7dd11a984;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1504a989a3d70cd29f86eef526d41a14b1e02238c936824128107810ad31b8d411ba40509;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7aa0b7b3ef2ebbaa3508d265493a9e7b55ee0d67ea102af7d4e2848cdf155c8c425db3fa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h650a269ced16cb01934ea8fb6cd08c8eaf2cf53050bc2a0efd98010ef22d2eefbad1b85;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c2c2612bfd3f43c36cb42d57dab65995418849f0284df95dd397f723e6122e2bef2bb3a4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fbf6d9251fe513ac54b683770343c979355ec6155d65dd7abdd746d729885a48aff41392;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4c9f7b2260a7a2f0f00956aa43bb78adc0a9850e7792c37a3cc8fe70fefccf755c927a0f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfe332b03842d645920edf40e53498e728f4f17b98e24ee7d93615a5cfa514de3e7805a16;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he4153adde20323df1ecb1cd705ad392dd88257d013363448ed4df5ee4593f68e4948e9eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13984f0a9163652b657465607ece5957b689fdec7eb499dcef5c18e55b09e9eabc46b6269;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1617220e2268c4221ee60fa86146b481ed9a914998b179ac5f94c0d62e0cae6b18636281a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14b92ab69f9eaea7731f4311caa2935209c08728734a5865ba0e4c37707ea168fc7821331;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4fb6936abac1f296f354fa5b60bc83030ca1393df01cf08701f9ff21c335ca75cc7988a1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1916b9863505a40e0c3567731eaa2daa6f93733c556c07d5308afbc453b55a9bd38eb6ca7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haa5897ab3bd43ab345bd272aebdd4607bb0f002c06ff699e7816447c3e0bf19acc8ae298;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h636ef491179871686e6fc120d2c5f6476973a49a1655a0a7d2b1eb8cd245870a81845956;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h873acecbd478d0bed47a402048337e24329cf0f7594511da91132596063986bdbc927f87;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19bea63197c3ec4682ba58e878eca379842e482f91176203eac499743d112b7231d2b6612;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18abeb52273d23b5afddee6e3bbbb4b0b279a2aceaecee9913b53a0f9328e0aadd491abe7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10b99c08ef63a3940fa76803dd7d64924937096bc4a32006e9db8ec0df32c760a17044334;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he641fd8c43c8acdad8265b3656780374f90f467755c499a327bb203bd2e1983730f09c6c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h123dae68a6c0d503b60dde232adf4e0740bd4062be976458f5869f538aa284ecf652f5341;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h195235b0c578a059a4c06f450cddcfe59390efc5c21af38de5e71bf31e74ebabe4abd710;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hadadd10c0796961c9e6111151d62781f6936d0af6cb47931b7ea384ce338e4a6c73ffc20;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h155bdddda3d1dc8b384601091b787cbda444ecbb027d29f9d8a5c5105e781769094a6d2fe;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e4b6bfd0683555b375b8126a95c0d3670edb022f08ff251fda393803baa655cdaacc9b6d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb7d06668dc01881586443d61684b766bda0331e9fbc1483f8ec25e6bd2c82b78fabe7618;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c74d30d14fcb769d9559c86546a90ac7872cd98cb842b1cc7da2bac168000bb3fcf47379;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1db8f4147a8a503e20ece1932927d04fbebe1acfdf4bac035a6313ab8d1fe4aa2098750bf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1452e5f14e704e0e2b70a6ac8ed649a24907d1b076a5cfc81c1ebbf88fe7a7c5212bcb672;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d8c409ec023485f9ba6be5e6b3eb4a673704feb0d4bfdcc4668a16ca4f8dba57a7e374b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hebd7ae3b95917ea6fdb2f8327b387ed9e134c56d83277c44afd1e76bff46759be9effc15;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h190a94b937d68d95c246db258855f911e471760a41fac2009e941766017fc58ad79504ef6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8090cfa1c71738689877c16771cb1a6a433f81dce374b347201e97f245ca85b59e5595cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h140ed9b747185880681ea6051690fffaf1a160449d9e96bcac60d7824e5691ea303edb388;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ba5f6851cf38157f544e5bf40899d94e7142faf8472951d70c3895e4af5f0a870b13af26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h102e6f2280332e8aced48229859218b45d8528e01307427350fe41bc9e7c153ba686458f3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbc41fccac51f3c4d37ae2a47800732950c0de79b95472034f3aaeb4ec5339cce19a514f7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbaeeb05abc7d794ae03f9ff66ebe90a8885897850ae97421315182d94304af6397becec8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17779ed32c1b7ee846d6583127c82b3a26dc7c371c76c965477131cf10f4bc408fa38dda1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19394b1fc50f3539cacf1ea89191fb363e93db1d41eeadab9da60502f07306df150096871;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h5f33aaeb0ca97a4f55751e2f81aaae4a1855a1d2f6dcf13a3409d444fff8c4fa42812313;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1604628c38e50584a080dcf9e83d776b4967ad5e390c1a5871471dbfd7fcd321c2e50d8c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e20e7620996187001303f0b2ee4de99e94f45d385a3f8a57533d3737caac1a32e6226b8c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12a51923687e769da5dbfe41474efbcbef4fa1746cc2df0d6565c162ae0a49877b85a01ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h779e186c0bd8c65d8aef805f2dfdb705a47b3b6b1d6c228ef31fc7844de6cc80a0bd82e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h131535a7decb9accb9aae3ec7b7e7fb4f3c52918e982d3ae9624be032858996c9ff2f0486;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1563b5b5a169075b6a0add856d37ae08f1e03fb7b210f48061fa77a1fcc12a88fa25b1f79;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6025780c6a1dd5cd490015c75a0637158ea92b56062fc3123f2b99da107a23ff950b56ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h96f30e29de554e1d6d6e4603609bd40bf9f2aa67a5334852e143aac5a25dfddb25bf69f2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c6f1c17e6f21e314e0a5a136eceacbc027700881c4dbfe7db957cad05efb7318c6d7c24;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h71829e1242e07fccd52aa08a0e5dd172475a2bd555e29dd78c959642f2d4b6ae90045c13;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h138f965ba8741b1d5631c427c26784fcf33475d1b66d16731aa8df120e6d7d27515910bba;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1666931ed2a60a6470476d1e820b68a2bb446b94eea7cd54111defd2a6fbd0dc880623fd9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcbef50f473bcc2f1e6fbd87bdde3dcb0ac859652b8fde053f0cd735026ca1a747f5bbc55;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h187763914af7c27633295ad5257cbb29f82a9f7ddf991c16b08fe88637c2a841e1844fb3b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1926c081a417e76e33d1f2bd247a734768bbb7250436d295b50d509eb93ad4d0ebfe299df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ca6f60af95113b592479dfc679f3e4d408f1cf9af6f86cc1682f7f80730922075fc79780;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2e6181e15db1594c06cd8d46d7ba3fc6d19451034c3fe85aabfffe2d647f4fdd17520d12;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6643fef84098242daf3482f5d1ad86cf770adff7ef1847f64d8f1895669d198e0a0d48b7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1305babf3673cba5199563d5c53fa7e5b45e5b397c56b7e48af934f8cdfea0dca9887c69d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18f064e9ef4474f20bd030457f73228edf2edfae452871fc38635c7d3d27e34aba5ac0391;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7b5efd76724162964a0ec8c0d07ee1bb4507a83aef3e83e5b195c9ebb02ce6a0d97bf7cc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc50a24e56080e9e13637740dedc1d08d1bd36667a70dead1201b605ee02216f4b5be06ea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha98695364cbb2544406379d6bdcaa37c3d9bfa43490dc7d0b33eb993249c539bf548cee4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19c5cd7e0c7ffe3a678170f5e5608fa66a499ffe43bd3799b4a53e522a70eb80bd4bb2ed3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a2d569a8b583107e71858530f341cef38d993599c4cab2f75c74f6dd13652758525d49fc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18111d5667951cd4de87694c1079981e76c1a8cf8cc9097e030f0ac91d2ae0ec7894f3491;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd975ac2d9df13a22721108a7a92a2b7266095832712a15605e55729ecefb081c10354d31;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f0afeff2fd899d90aa0d35cd55f350b41e6384863b88cf48788b85cd3568783c5a4faf51;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a68cd77b66275009960f49ef5df5765f93f0b4ab4f70f21d71ef49f128c00d949fcfd3ca;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15581b4305617b047bea1743bf56edea316fd72e47f28bb25bd18ec7ce0a49d2f11441494;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf859bcd54faf9a36d0fbe3cd1aa4ebc368399bb07e52b434f0bdfb1bb43aa30908b3d018;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h160bbff1c69e9251f3987bb5c77c7a1f00c8b8ce2ffcd3cba82f01822d08c19424cd640ed;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dfde782a919cfcc33be48c39b520a4b27a4febcb3af1357540051005612dff259310ad78;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h128583a36f0a1f9c9c452528b47d37b5a3995e7c91358a1136e3f2401cefac4844d2403c7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h197e7de2cd5535762d47551e0c677b1174b45e0489d012aaddea6f85b7a33701ea8a0e3a6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h3e10cf0bdfe45e532262245024e3bfd8c56e9b843ebce63fe44b73655a02bda71aafa3df;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd9162a6c2ecbff5cfe4658df082736d92ee729f7224673fb8d0486eaed20f591405a884;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4b75f1394c12172ac015c014138a89952b94d46e4bbe9dc88e78a7adf1cb7729a6e04cdc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha10bb0608e0672b1a9b0904f6e85b58d3897657a1e14076366f750d694c5abeb6b52f2e4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h113e1c5729717d41431d58c6a89a0b56190b25b0ec63b55f9ed928e8d2d8c2f47effc2f9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11c1abe8ae77151ecbce2a0822102ef1cc0dfb210a0d75165f61eedaf3d3ad68b7d74ccb3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h195c309ba33769d842bf31fe4996f201d7f782aa2e1ec74b7ffa4a472acb425e3d617cbc9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha370a7adb9ddc53f636ae01528f4c352e8cdf715f3cf1737f2b49e1cc599d4bfe4b78db3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f2c1f72e215aa96676ec0958ed8aa8e364bb0f6723c103ac7e33618c1940eefd8f20e00;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h47346de52008fde05cd68811286ddfe802215a45977d33f1be349605035cee6af717ce3f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd9d5e059dcdb6b0d8da451a262de2fac7706ebc5db5c1a95a0c5b5b614e95de4f4fbf98e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbfd74686a675f551f767626c828e0475c7f4e0d49a0c5072c24b4ae4c86f897aa7cc9055;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a6fa0ed025b1df5c245420a68ab42f21ddd888591c2cef0ed278c1583ea27b185d5cb1ce;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h199958da438e57f1a95b0d48253450f4e05db78452d93862615bdd8cad4278bab5b0febfd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he77dd690af510a25ac72e1142c0f7d06be58ef8590ed89bfb539aad39e9d0844831b5c36;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h173811bbb1556d1abde506d1afdbcb4aa3c9a479e3008c83d6f216626e19265fb4992a3eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h352b22245bfb08caa838caf6b89efa5fb39e5af49396d9ba34506ad998a2bca148674bcb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h87c3a42962a645534e7f2048fd287d48d811bf59b210a40ca1a846355a78889160b889f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc7313ae38face9c65df3121b2c5b5b45793eec7e9df5f71202e8e5eb3bac4303fc35d1f5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a664d43482f34324072478b38b521815ff173835bf02c21109eef66ca3b33907b12a8800;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'ha1cf9ddd11c2a3db974f9851eecc3e3739ca10159aacec7d15cdd6437b047df9c388cbdf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h65a01bd3d29635be90bc9f83e5dff6499178d1dee508c38d77292f5f163deaa5a2f44218;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12f5a7af9af36f4e35cb14d7f715298d13564123d341c2894582fd0fde91b51854f926c26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7cfa08ab1273245050b2647c67b980aa317092f5919b87ccbdb07863e5c63dcc1953be59;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h31e4a10f3e468dad91dba994e9da75904aed2065c63d9eb6a96ff7261900af4e8bcd18b1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4192a7f1705a182da38709a1aeee5cef1df70bfa79a7de6627e671802585b87b5991c8f8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h102e7601120c99c70cb50f0e8694615a4f908fb4a7962b0387fc37283ecec944454128bb4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b03e283182ea87f73312c60d64cc6dd364e56a91d56d144115dca6ba4070bef254a4c59;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1041cf36a8b640ae8ad0162f72bb9db6e11b0bf53e8de6831c2d86084558eadf4dfb41d91;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd39ca6dd08c763d512f320bcee5b8087df9ee82567567ec70e636f74e73ba97315739418;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19853de04694ee3ff9866e0a0cfd3ae4d0b6a89a9c5df587a81eb11248a99f813c2b703b2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bd5f5ed87cbcaab1477e567619b1abfe67664decc97b720958c91b95607bc45deaba9969;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb9ad18668be5f601656a080d1e27b0932110aa05d0db76a76d3275f91143ce617af503ae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15085127cd0bbafdad2e937e23c6f44bc39fe40de2506421d5672140a8e73bafd6e97c5eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14318e912ad8badd1ef2b58aa23960d800a394bc1e72658c361f940ec2727e3a2688d42ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1dc88042e0d1d2291bfee98c9d6a4de76168183bd3c81c47e24766aea2a0ad97e0157cd2f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1675fc9e57428f9b881d5027d3ad622f2eaff06d2ef56231b975edd02a2db140de8895150;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4e22c3c4a2906d7b00c63db5e215f89648dbf6cd0c72213a8e9549f22f44f986ad5ed2a3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ebf6624f44c78565a969b379924ea425fdade08b47e63e18baacf1978d9b0727283abf10;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hdb4e27ad695f657f54b4a8678135c6088d6075a4fb5d60ab5f68c31419c1895b566ca2d8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hff88aa5c1dff70a926981b7a3aebd56770779a1f1831afeb642a0968266746acde846c6c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19a273fe377ab494e5cd1a43bb04a751fb2f4f1f4a638009570cf1a14d46675000217e399;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1d170b4dac0ab3677bedb9aa510c481247a3ef20d0f6a6605f1a0cd99cedb63721d42093e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ac8abb6b1dc398f564a66f7a6c1442d2f1c98572bad22dc64e45c9fa36ced0dab45b1465;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15d67574d8301ac5a3c9f8b76510180f06a0d0ca51b757be20a18d7985587a9a8f8df2d07;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4a373bee571a260f184809ca5994f55db37208ab17f11b5a344cb6ea91699353a0e1bbc8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h174260678c16906ca0bf0287ce7fa9710161bcfc498f3cd40fa6eddd093a042d0859572e1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hbf9f60ab97c8d56fbac64b80f97eb9b125ec066694e4fd4c0c7c87b7a1da9c56a78e28ee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf7c74f688d5f0c8563510b91115cd43aa084e94c7b14ecbb6f6938d88c86556a4477aa39;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'he89f598918ae3d349de2cfbb43e64135a2cbdb9650e8434d410d8f4c44d61aced18bf960;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfcacdc7638da483c4e699d4a01234bfd585c77a1986dd34eb9d7ef7acd72ed6ef6b24119;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7cc33dcd6d10eea259480e2aed2691ca980993dac0656e05db5f1b7634c3a64f76ef49cd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f5cbaef8ab46129a5325e2eeb2678cd9da3b2de84bacb35fa19a8b1f91e4262b125cdcd8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h116181349e7518fc16b453450617b4b1e0da3912c0c385157748abaa2825a9d43d79da366;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h527dbc648112b436fbde4de9372f083dc0b57a41f56545b80a6adb29ed63788b50fb6206;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14e0d6de056cf297ea41d27c9a0ddd4612db4a4a9308fc9b550c2cba7dbe719b566e89e4b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6273935bb07fe095137136f7f1dcfed8b4fa35f21991959a83bde32dc364d3dc28b7f5ab;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd5c74ef02f482bade66984b61cf43bca241a935fca8b63dbb3820bdf8692caf98ffa2c33;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h626083ceff6c0d42e02da21a39088e8c6ba4e7be6ea79f7881baafdf99460e1f2c9f5a25;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hee99d20f0521301ae737a1b36f89f1430bfeb8addfb2c01b294cbc1075e5c093acdc5f38;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13e82156a877285991f74096f5092015775d828f5344924c878e1917a4f5c89f5f3df0993;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a66078e89e248e0f5461333e08b9947166ca29335facb8b6053582bede2c259cfaa04418;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7c62e1c7f5e81deda1e0495ebb0079459214913280d827e29695e804bbf7a93ced0fe235;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h63cef47df2ccef0293558074ba1dc19b4a86f2e3b6966550c5b2c0a3ee95cf3f7e543b90;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h61ad3ab339ba2cc6c4f829678dd50aa9486356d5447baf0ff5c98602b12e8ce8c7dd78e8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc3af9f2b5cbe4e07a8ee1609dbdc45736745ce7dbd622a377d09f024e7fbc4b517ce81d6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e09d7acec4dfef68d907d33e27d9bd494edf78266d1fa9f514290a2d58e84310656bc772;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h291716d653e0918620fc7ff3580eadd63de613a9e5727cd1b47d8498325ccc2027b174db;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1bed5f7ffe313e2d8516a2e8308ff1094b2cb9e501be487a5b30a2b9e4996d20cb17a1e5d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfe68dde0cfe6dd4de5daff165d7155933e59cbc371a2e5e684cccb67d704b1b0d49ac6d8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2118309b02bf6ac18fd71905e0f5592dc333c7e9db892c17c5b35fb810123eaf9eebf517;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1297c2d2083de8354c4f7612b225b2479fdec4727fabd76ffd500f7595ae3903e48c15eea;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf505c3d70ebaa0ed4b3b7157b5dc7ee050dc20123fdaa8c9b1eac0b744f078849da7ca04;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9b1d0d64ecc17ec693846403f6bf6c6394764f26410d0355f6d6ff358e2372ca08fbce44;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15baa01a90e772aeaae99ab3b956c1dee1b1096bc2f2b6d6ad2fdce4cb77e354569b2933a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h120c0e37fc5c5b5eb81e4039194ab7f5d3ee502adada63076f665e9fc3fc1e11f441b055;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h143105216c9559e951f9b704629bdc282464b9295c6a055c5a464a1b1f202be9215b5fee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf7f4b6f66bed2c0083eab97c46470ec8a7746d8be858e448b9beb5d6b7dc5f20babb9e18;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1902cb0bbe84538b48ee811da7d2269a8a6ea3f2fea0ae265ae57323421a5dbd949cab1a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f5382c7200016f63f0ce591e0695138eb0413e3d88c3a0078370a2e6b1e67addb879c3e6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h75f62d48f6217ce271924600fc074e9588d1ec9bcc62d8fc8037da8df181367a82953ebf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc8a1b61ec5c7ee6e80b21272b554ae8bd13d9d33345dd4a8597527ba7367648a1333aa95;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb89c4efc70974439c495657104a32841b302f362487887a67de56c90cb07a51dfde54ec4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h135c6ac60a734acdaea03fdad10bcd1b2a52539f0b7a33261f2096ac4462c96a5a96cd9b2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1e9e628b9a72cdfcc49cfcbaa49cf2d788b99c88778ba652682f3fef6acebb343270f87b9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h97cf699b0f68e9b6b79abec1d26f9b82a83bfe8b61b7e6deb6319f72cbe9af9ac33c6e5c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hfc750411e50e7c141ca34320a2bf0df77a0a457324891474d0ff7f07b560759d61462848;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h11277f4ab7e4fd4f5778b2c967cd50c49dd0d0bf79f50f066c4ae43b1f886d1254991d04f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10d31c4c6479a60bc5ae533428fb20353e42c9be45ff1b3330f331f02615f9b165d67edee;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'haa8f5749650d111afd65650020f6ab83961e961471a49ca3956064f01120338932ae91cb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a1fce77652ea4c23905d0af5782e3dd6b0c2a36b8e699144e19645f05ae55c25d953466e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13230552a82ab6ca0bcd7ef7b9554fd285b79f7cbcb3f769ba1b5e6725693f3b739cc514a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'habf764aa77dda9538192bf2159e05c19f52d3a496977c03c25a93dc7ada47b72d0b11998;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ed2a7e3b58eba5568f2c4c7e3e331f64f0fe22dc765d086769dc9a18dc4cce7b8d7613ec;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9ecf7ef946a47aa52e7f0e306610e5dcad907a3a846222efee9298082fb4b4449e91d10;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1444ce30b57dafac31b5601c3be06b1ddafa4167a5c1b0ff86e752e85cef58d82c0298235;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h35dae765c9fac4471669ce29ff4bdd065cce0a292c7c61ff675966e298bba2f0dbf84f35;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf245c32f53b4fa3636daf49934c6850762ad96384838e6615d2ce0a24bcb68e4bbadf1a0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1ef81c0f5a7b4d920eb050540eb1354123f36dc4a492d0b51c661e1935b2a7e254e57984c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf08b1673ad8f51d9a70154539c0dead38e3f91724fac94ca0bef1590275cb0e78b8db928;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h187cf65213414696ec66b044877186d56ed93ea61c4a442d5b954498d0d5ec1212ba09982;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9bb620f1f902318a9eaabbe44c5ff7786aa949f99084aa491821fecebdd004995dfae615;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8168c588d2d86b26033fcb6f1afaee57d5e185f351f29d7edaa0c612aa60203f26bb86c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hcb411ced2616669386a36147ba4c59d5416ada64a97ae0f53970431baed9c16290884ef0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h16e93a96b6671a7546a8804f87abdd2e26de2abe51e93e5bdc1a1e34c3108df6e87647739;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f22cf2ab78937876e3d4c7cd65908ca82e94c49a5ab48c8fec9f46748f613e68909e5d34;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f2fb8d5b26df605813a727ed877743c07e72126a5bc7564318f5fe12d390d51032006d80;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h8bbf1f73e88770b8c4e8ae5324b8db54d9dd8e799e672849187c2bdf3638f5f692056d0a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'habfb998faa271e8b4dd1ff3d3ff7df8a641f43f5f6c18206455a78832a0bcd53f74ea31b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h18d5248583d098435d79d81e244bd1d3afdfd2609bcb7a54af11e19cc71000aed7e7ff0c2;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hf061f5777a55c422c8f22517d2f580327148a26d63773d93116e4165593f36f4054bc90f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hd9f233347b820d696c23a770d001a407c210ad0df97c2b1f7d8368537a3521323e86f7d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h100c1837435de0f9a1df70014358c12638ce7e11610cade53882092115eb6b4f21b81da7c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9831fda3d55f8d2053181e79073278e80e4a1e6b8226ccbc436a1b22e87097be897c6722;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h76f6c3b7efe63594e43da9d48568fb00fb71052e6cfb076ad11dd7f1a87ee62f3715feef;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6e55e5c8438e3e8e45045fcbb35ae16e785de527725fb608b4fb0656fec293bcb0dc4ca6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a313de3596f35232e04ce46a521148394a3ef7e8d867f8675234e407769d0f73c604f400;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14abbf5b3a6b2a146c9db3ac8dee941c9f241352cc389ac4bd07bc628c13104da6ba7d5d1;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h415a05123c27d3aabea86927d651373f251e0bd599777cceb90e8f5d695a783bce4a66b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h19d9e8ddea104c51e48007fcaaa37f08b546831720f2c0514e0518fee25d36efd4983b44a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hace4cd2eeb6f5677dcf10bb906b3833cb88298757fa297a193b7992bca174feee0a5ea1a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hafdaf4879f065d827648f602a245297a4432287005cd0ac49fd4365eb4794fa716a2a2c4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14dc91c16403de18fb597f1e01309166303a9ea04a53e4dab39b86071259f5332685f3229;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h368f76b2e68e27f7c9662a606642089be115fd63511cef2a88986f7c5618da2b923f558c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15c980137a6829e3fb96fd44ef30ca6e6037b9364497cbc4eb729b1fbcf5b7cd282bf1de3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13319a39bbc72154065781c12037c41543ee40fd45a80875c907b59008968e08d7ef7b30c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h127bcd4d43dfc6ae395cfdca3a8f719ab6dd9e586a834e4f142a7d453de0720be69732dd4;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb9c412d69a335fe634f3028f8b973046745f966bacfb8f2daee871935a7d3c2a3012fe79;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1cdf70385d5ce86a7bb3da915e0e8c646b8b46808eb5d792834f12d00d4bf47a1469f13a5;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a4bf238f4ff08690289689852d98db0cd3cdab1204ee2a121dd6963309e0a8f922f8d7d8;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1f51f2029a985338869891682b02f7bed36b9d6c4e05eaf8ccf8ad366cbb88579a00d697d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h60e10c5c54bf4e57c8dea794a8450681c4f91df579bbe290b3e63ef16220f99dee1579dc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1b7579ba8d7edd2c07acb4375d4623625f51f69c9a3425098dc0c5b112f209c4f8c6a6cbd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h446a673462d40f0bfe885df4bb3a7cef884a4740edf1df78bae76e79685eb596aa175d1c;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h17f9c3a0f780a97dbcb8e758ea6737eb7c1d91468a4b6d9edda3dcf6535fcffa7840492f6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc52085221a5a882e4cdbc79b3710e09156c9511ff0b040d3caa0cd5868453fd63753dc4e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h52b7bde32725a6857350719363bf331b53ac34f155e42989494933206281381c497f45aa;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hda417b3605ad41a338220f4688108818958e72e43b5cecfcd86b5f194f642cab45b66dbf;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h136b75aaf2fcba3d985053108e0edb1ee186adc6fa5a9aad5439eaf75f12b83c8e034de1f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h7c78297ff378192c23b08c299984554869c8c9e6f5949c299964297ced7dc067fa667b70;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h10f874f9b47d3483f8b8d2f886a5ace7f8c9da91bcbdf24345c3889fb351c05341e3ea1d;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h12b1d1f76ff1c1b318e345f34c879849d49378544a3f5c1985a2f242ce70b614a7445af97;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h146155f6d36a1bbb5424b943b379868d2266b045793f179f96bd0816fda64fe53913d8f9e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1a8e97a6cd1d8a1c2582edf7b175614de3924f064f5b0945a3aa4d85d5fcd09c0ac3eaf7;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h28e237a085ced5b32c8a107df313df2b8aa63f5898ed1434958dfa11918abd8c03bddbc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13dbad6954d1417b0de903d9f72959175bf377a601f679aaff7494953715dbdad10a9dca3;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1aac03df0204b84e4c4cdfa90da65f16c58b3bfd4d9beeb646c3dab5f9ddb3bc6883fbadc;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc5b2da4994ac0585236a3744aa23f7dfd74afd9d46c6c629d496f0024aad18efe489f4eb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h114f3e1ce9db49876da864c885d7951adf9231815590933e3cd7c79bbefa397d50861bdae;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c538d84b77ea26773e667510873f993dcbaa2a7df881b9a641d358a1518f387265238ac9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h14a7e1aae63dd484ff489d0eee6e37c9ea21b1f5373d6e45ad712afa81be3e0af6332c51b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1fac7022e8cee1ed3f70b0cc47b4919286020c40da1b11dd08bc24fa9e29604becdda4c36;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h94cffc386cd7967c0f3e8904e449a63fcc5129c551b104e499578d8701c37e03553e9bbd;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h308fcf863dd4c04da8148d5225cf10816e370ba65e982cde884359f74878dfb7fcbdf26;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h178ea1652a54a6f69e2891bf99cd1253f8e2ea6450c3ad06e7d8735de2e315faf685ba30e;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h57614c48b74cb675174c0df23673013531b353211c791bb3a87ab8ca7a57f18e72e55de0;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h4c2a8b3a150a02b65339dc550a537b306ac097fbac93fe8e9925ef073f2d046d8ef19124;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h9c0e36cf723e10ab6924dd15639114f1a9b9aa0a4069e47a501c7af745be702bfa08c958;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hc476b21112143339b6fc97a55276570ba8346ec950ce631298e2d0aae6ccc15cae88438a;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c7f7f2583be4ded08576b15b6ccde55de4d4538fb31cea6e5870e663037950f878eeb084;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h776a9eed5ea619d4027ce329eeb4cdcef2c50cca3ec33c5204ad3233e44ac3483f2d61a9;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h105acaceb64a31217ff3fa4facf1ed02cf0b51a99496ad3e359bef66e89718d396dda582b;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h13eb139c1b85b2c9fe68db63ab8d28f66abcb5cf15ae1edb076d6d8c99b2329cc3fd5b90f;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hefff00de926b3ba6a64b221919a58a53b84460a25ada0645cd966abc64f683b817983bb6;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h2215da7774d05040e3788a3b94f16823f20d3712768f873d3753d510d64a322594e92501;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h6fbdfcf9e1fb4d8d9cf65eeae30290cd0edb35e6af893921e44316052c9370c42f25c96;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h759d259a2ca2ecbe4788a88a0bc7190bc2046e7169470a37687b6e94d3b638f26f629166;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1311a17388242ce961fd181a09c6f4aaaf6f86ebe08eecf2e3b2c6d7fc338537e0da84f57;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c9d4fa8609c7f22fd9dedcbd9f6d9f5b3ded33e3ccb672992a8f2b160ed577331f7caccb;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h1c2deb9091b92e5b3ced1db3851d68687858a093160b8104843ebd33c7a2d9ebe721db839;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15305ac0dc80567100e593e8ed993f9c76a0302c8844926dab9695a633431eedb6cfbae40;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h15438bfad6ca7dda2e69ca3c435095e740ccb5f5f340d65c60de7e49a5c700d9f5c477258;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h59384a442b3a968ad9188e64bafbcc6dc09a08c82c5061025fa72b747f8c281fe3c0459;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'h177a9bb21270e6c1137a21860b6c8a57e629622ea0034618c264f6b27f9685e0282ee5386;
        #1
        {src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 289'hb1beeb3c59a58e5f75294a2f0dacaeb2540d6c2bd1f2e9c90bbe5038845568a45e348b80;
        #1
        $finish();
    end
endmodule
