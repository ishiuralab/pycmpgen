module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24);
    reg [511:0] src0;
    reg [511:0] src1;
    reg [511:0] src2;
    reg [511:0] src3;
    reg [511:0] src4;
    reg [511:0] src5;
    reg [511:0] src6;
    reg [511:0] src7;
    reg [511:0] src8;
    reg [511:0] src9;
    reg [511:0] src10;
    reg [511:0] src11;
    reg [511:0] src12;
    reg [511:0] src13;
    reg [511:0] src14;
    reg [511:0] src15;
    compressor_CLA512_16 compressor_CLA512_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24));
    initial begin
        src0 <= 512'h0;
        src1 <= 512'h0;
        src2 <= 512'h0;
        src3 <= 512'h0;
        src4 <= 512'h0;
        src5 <= 512'h0;
        src6 <= 512'h0;
        src7 <= 512'h0;
        src8 <= 512'h0;
        src9 <= 512'h0;
        src10 <= 512'h0;
        src11 <= 512'h0;
        src12 <= 512'h0;
        src13 <= 512'h0;
        src14 <= 512'h0;
        src15 <= 512'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor_CLA512_16(
    input [511:0]src0,
    input [511:0]src1,
    input [511:0]src2,
    input [511:0]src3,
    input [511:0]src4,
    input [511:0]src5,
    input [511:0]src6,
    input [511:0]src7,
    input [511:0]src8,
    input [511:0]src9,
    input [511:0]src10,
    input [511:0]src11,
    input [511:0]src12,
    input [511:0]src13,
    input [511:0]src14,
    input [511:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [0:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [0:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [0:0] comp_out24;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], 1'h0, comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], 1'h0, comp_out1[1], comp_out0[1]}),
        .dst({dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [511:0] src0,
      input wire [511:0] src1,
      input wire [511:0] src2,
      input wire [511:0] src3,
      input wire [511:0] src4,
      input wire [511:0] src5,
      input wire [511:0] src6,
      input wire [511:0] src7,
      input wire [511:0] src8,
      input wire [511:0] src9,
      input wire [511:0] src10,
      input wire [511:0] src11,
      input wire [511:0] src12,
      input wire [511:0] src13,
      input wire [511:0] src14,
      input wire [511:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [0:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [0:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [0:0] dst24);

   wire [511:0] stage0_0;
   wire [511:0] stage0_1;
   wire [511:0] stage0_2;
   wire [511:0] stage0_3;
   wire [511:0] stage0_4;
   wire [511:0] stage0_5;
   wire [511:0] stage0_6;
   wire [511:0] stage0_7;
   wire [511:0] stage0_8;
   wire [511:0] stage0_9;
   wire [511:0] stage0_10;
   wire [511:0] stage0_11;
   wire [511:0] stage0_12;
   wire [511:0] stage0_13;
   wire [511:0] stage0_14;
   wire [511:0] stage0_15;
   wire [100:0] stage1_0;
   wire [179:0] stage1_1;
   wire [172:0] stage1_2;
   wire [245:0] stage1_3;
   wire [240:0] stage1_4;
   wire [217:0] stage1_5;
   wire [206:0] stage1_6;
   wire [206:0] stage1_7;
   wire [217:0] stage1_8;
   wire [263:0] stage1_9;
   wire [209:0] stage1_10;
   wire [189:0] stage1_11;
   wire [221:0] stage1_12;
   wire [281:0] stage1_13;
   wire [244:0] stage1_14;
   wire [271:0] stage1_15;
   wire [126:0] stage1_16;
   wire [63:0] stage1_17;
   wire [22:0] stage2_0;
   wire [40:0] stage2_1;
   wire [59:0] stage2_2;
   wire [102:0] stage2_3;
   wire [116:0] stage2_4;
   wire [93:0] stage2_5;
   wire [103:0] stage2_6;
   wire [84:0] stage2_7;
   wire [86:0] stage2_8;
   wire [137:0] stage2_9;
   wire [85:0] stage2_10;
   wire [143:0] stage2_11;
   wire [84:0] stage2_12;
   wire [140:0] stage2_13;
   wire [124:0] stage2_14;
   wire [84:0] stage2_15;
   wire [104:0] stage2_16;
   wire [61:0] stage2_17;
   wire [25:0] stage2_18;
   wire [10:0] stage2_19;
   wire [5:0] stage3_0;
   wire [11:0] stage3_1;
   wire [16:0] stage3_2;
   wire [28:0] stage3_3;
   wire [39:0] stage3_4;
   wire [47:0] stage3_5;
   wire [37:0] stage3_6;
   wire [45:0] stage3_7;
   wire [40:0] stage3_8;
   wire [51:0] stage3_9;
   wire [63:0] stage3_10;
   wire [60:0] stage3_11;
   wire [52:0] stage3_12;
   wire [41:0] stage3_13;
   wire [57:0] stage3_14;
   wire [56:0] stage3_15;
   wire [49:0] stage3_16;
   wire [31:0] stage3_17;
   wire [25:0] stage3_18;
   wire [13:0] stage3_19;
   wire [5:0] stage3_20;
   wire [1:0] stage3_21;
   wire [5:0] stage4_0;
   wire [1:0] stage4_1;
   wire [10:0] stage4_2;
   wire [10:0] stage4_3;
   wire [26:0] stage4_4;
   wire [14:0] stage4_5;
   wire [21:0] stage4_6;
   wire [16:0] stage4_7;
   wire [25:0] stage4_8;
   wire [24:0] stage4_9;
   wire [37:0] stage4_10;
   wire [21:0] stage4_11;
   wire [23:0] stage4_12;
   wire [25:0] stage4_13;
   wire [18:0] stage4_14;
   wire [21:0] stage4_15;
   wire [30:0] stage4_16;
   wire [21:0] stage4_17;
   wire [12:0] stage4_18;
   wire [10:0] stage4_19;
   wire [11:0] stage4_20;
   wire [3:0] stage4_21;
   wire [5:0] stage5_0;
   wire [1:0] stage5_1;
   wire [6:0] stage5_2;
   wire [5:0] stage5_3;
   wire [12:0] stage5_4;
   wire [7:0] stage5_5;
   wire [16:0] stage5_6;
   wire [5:0] stage5_7;
   wire [9:0] stage5_8;
   wire [8:0] stage5_9;
   wire [14:0] stage5_10;
   wire [12:0] stage5_11;
   wire [13:0] stage5_12;
   wire [8:0] stage5_13;
   wire [11:0] stage5_14;
   wire [14:0] stage5_15;
   wire [16:0] stage5_16;
   wire [6:0] stage5_17;
   wire [8:0] stage5_18;
   wire [8:0] stage5_19;
   wire [5:0] stage5_20;
   wire [3:0] stage5_21;
   wire [1:0] stage5_22;
   wire [0:0] stage5_23;
   wire [5:0] stage6_0;
   wire [1:0] stage6_1;
   wire [4:0] stage6_2;
   wire [0:0] stage6_3;
   wire [6:0] stage6_4;
   wire [2:0] stage6_5;
   wire [5:0] stage6_6;
   wire [4:0] stage6_7;
   wire [3:0] stage6_8;
   wire [8:0] stage6_9;
   wire [9:0] stage6_10;
   wire [2:0] stage6_11;
   wire [3:0] stage6_12;
   wire [7:0] stage6_13;
   wire [7:0] stage6_14;
   wire [7:0] stage6_15;
   wire [5:0] stage6_16;
   wire [4:0] stage6_17;
   wire [6:0] stage6_18;
   wire [4:0] stage6_19;
   wire [7:0] stage6_20;
   wire [4:0] stage6_21;
   wire [1:0] stage6_22;
   wire [0:0] stage6_23;
   wire [5:0] stage7_0;
   wire [1:0] stage7_1;
   wire [4:0] stage7_2;
   wire [0:0] stage7_3;
   wire [6:0] stage7_4;
   wire [2:0] stage7_5;
   wire [0:0] stage7_6;
   wire [5:0] stage7_7;
   wire [0:0] stage7_8;
   wire [2:0] stage7_9;
   wire [6:0] stage7_10;
   wire [2:0] stage7_11;
   wire [1:0] stage7_12;
   wire [2:0] stage7_13;
   wire [4:0] stage7_14;
   wire [3:0] stage7_15;
   wire [1:0] stage7_16;
   wire [6:0] stage7_17;
   wire [2:0] stage7_18;
   wire [1:0] stage7_19;
   wire [3:0] stage7_20;
   wire [2:0] stage7_21;
   wire [2:0] stage7_22;
   wire [1:0] stage7_23;
   wire [1:0] stage8_0;
   wire [1:0] stage8_1;
   wire [0:0] stage8_2;
   wire [1:0] stage8_3;
   wire [1:0] stage8_4;
   wire [1:0] stage8_5;
   wire [1:0] stage8_6;
   wire [0:0] stage8_7;
   wire [1:0] stage8_8;
   wire [1:0] stage8_9;
   wire [1:0] stage8_10;
   wire [1:0] stage8_11;
   wire [1:0] stage8_12;
   wire [1:0] stage8_13;
   wire [1:0] stage8_14;
   wire [1:0] stage8_15;
   wire [1:0] stage8_16;
   wire [1:0] stage8_17;
   wire [1:0] stage8_18;
   wire [1:0] stage8_19;
   wire [1:0] stage8_20;
   wire [1:0] stage8_21;
   wire [1:0] stage8_22;
   wire [1:0] stage8_23;
   wire [0:0] stage8_24;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage8_0;
   assign dst1 = stage8_1;
   assign dst2 = stage8_2;
   assign dst3 = stage8_3;
   assign dst4 = stage8_4;
   assign dst5 = stage8_5;
   assign dst6 = stage8_6;
   assign dst7 = stage8_7;
   assign dst8 = stage8_8;
   assign dst9 = stage8_9;
   assign dst10 = stage8_10;
   assign dst11 = stage8_11;
   assign dst12 = stage8_12;
   assign dst13 = stage8_13;
   assign dst14 = stage8_14;
   assign dst15 = stage8_15;
   assign dst16 = stage8_16;
   assign dst17 = stage8_17;
   assign dst18 = stage8_18;
   assign dst19 = stage8_19;
   assign dst20 = stage8_20;
   assign dst21 = stage8_21;
   assign dst22 = stage8_22;
   assign dst23 = stage8_23;
   assign dst24 = stage8_24;

   gpc117_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6]},
      {stage0_1[0]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc117_4 gpc1 (
      {stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13]},
      {stage0_1[1]},
      {stage0_2[1]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc117_4 gpc2 (
      {stage0_0[14], stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_1[2]},
      {stage0_2[2]},
      {stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc117_4 gpc3 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27]},
      {stage0_1[3]},
      {stage0_2[3]},
      {stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc117_4 gpc4 (
      {stage0_0[28], stage0_0[29], stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[4]},
      {stage0_2[4]},
      {stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc117_4 gpc5 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_1[5]},
      {stage0_2[5]},
      {stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc117_4 gpc6 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47], stage0_0[48]},
      {stage0_1[6]},
      {stage0_2[6]},
      {stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc117_4 gpc7 (
      {stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53], stage0_0[54], stage0_0[55]},
      {stage0_1[7]},
      {stage0_2[7]},
      {stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc117_4 gpc8 (
      {stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62]},
      {stage0_1[8]},
      {stage0_2[8]},
      {stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc117_4 gpc9 (
      {stage0_0[63], stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_1[9]},
      {stage0_2[9]},
      {stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc117_4 gpc10 (
      {stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76]},
      {stage0_1[10]},
      {stage0_2[10]},
      {stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc117_4 gpc11 (
      {stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83]},
      {stage0_1[11]},
      {stage0_2[11]},
      {stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc117_4 gpc12 (
      {stage0_0[84], stage0_0[85], stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90]},
      {stage0_1[12]},
      {stage0_2[12]},
      {stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc117_4 gpc13 (
      {stage0_0[91], stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97]},
      {stage0_1[13]},
      {stage0_2[13]},
      {stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[98], stage0_0[99], stage0_0[100]},
      {stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19]},
      {stage0_2[14]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[101], stage0_0[102], stage0_0[103]},
      {stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25]},
      {stage0_2[15]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[104], stage0_0[105], stage0_0[106]},
      {stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31]},
      {stage0_2[16]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[107], stage0_0[108], stage0_0[109]},
      {stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37]},
      {stage0_2[17]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[110], stage0_0[111], stage0_0[112]},
      {stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43]},
      {stage0_2[18]},
      {stage0_3[4]},
      {stage1_4[4],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[113], stage0_0[114], stage0_0[115]},
      {stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49]},
      {stage0_2[19]},
      {stage0_3[5]},
      {stage1_4[5],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc1163_5 gpc20 (
      {stage0_0[116], stage0_0[117], stage0_0[118]},
      {stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55]},
      {stage0_2[20]},
      {stage0_3[6]},
      {stage1_4[6],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc1163_5 gpc21 (
      {stage0_0[119], stage0_0[120], stage0_0[121]},
      {stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61]},
      {stage0_2[21]},
      {stage0_3[7]},
      {stage1_4[7],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc1163_5 gpc22 (
      {stage0_0[122], stage0_0[123], stage0_0[124]},
      {stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67]},
      {stage0_2[22]},
      {stage0_3[8]},
      {stage1_4[8],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc1163_5 gpc23 (
      {stage0_0[125], stage0_0[126], stage0_0[127]},
      {stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73]},
      {stage0_2[23]},
      {stage0_3[9]},
      {stage1_4[9],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc1163_5 gpc24 (
      {stage0_0[128], stage0_0[129], stage0_0[130]},
      {stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79]},
      {stage0_2[24]},
      {stage0_3[10]},
      {stage1_4[10],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc1163_5 gpc25 (
      {stage0_0[131], stage0_0[132], stage0_0[133]},
      {stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85]},
      {stage0_2[25]},
      {stage0_3[11]},
      {stage1_4[11],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc1163_5 gpc26 (
      {stage0_0[134], stage0_0[135], stage0_0[136]},
      {stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91]},
      {stage0_2[26]},
      {stage0_3[12]},
      {stage1_4[12],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc1163_5 gpc27 (
      {stage0_0[137], stage0_0[138], stage0_0[139]},
      {stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97]},
      {stage0_2[27]},
      {stage0_3[13]},
      {stage1_4[13],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc1163_5 gpc28 (
      {stage0_0[140], stage0_0[141], stage0_0[142]},
      {stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103]},
      {stage0_2[28]},
      {stage0_3[14]},
      {stage1_4[14],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc1163_5 gpc29 (
      {stage0_0[143], stage0_0[144], stage0_0[145]},
      {stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109]},
      {stage0_2[29]},
      {stage0_3[15]},
      {stage1_4[15],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc1163_5 gpc30 (
      {stage0_0[146], stage0_0[147], stage0_0[148]},
      {stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115]},
      {stage0_2[30]},
      {stage0_3[16]},
      {stage1_4[16],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc1163_5 gpc31 (
      {stage0_0[149], stage0_0[150], stage0_0[151]},
      {stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121]},
      {stage0_2[31]},
      {stage0_3[17]},
      {stage1_4[17],stage1_3[31],stage1_2[31],stage1_1[31],stage1_0[31]}
   );
   gpc1163_5 gpc32 (
      {stage0_0[152], stage0_0[153], stage0_0[154]},
      {stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127]},
      {stage0_2[32]},
      {stage0_3[18]},
      {stage1_4[18],stage1_3[32],stage1_2[32],stage1_1[32],stage1_0[32]}
   );
   gpc1163_5 gpc33 (
      {stage0_0[155], stage0_0[156], stage0_0[157]},
      {stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131], stage0_1[132], stage0_1[133]},
      {stage0_2[33]},
      {stage0_3[19]},
      {stage1_4[19],stage1_3[33],stage1_2[33],stage1_1[33],stage1_0[33]}
   );
   gpc1163_5 gpc34 (
      {stage0_0[158], stage0_0[159], stage0_0[160]},
      {stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137], stage0_1[138], stage0_1[139]},
      {stage0_2[34]},
      {stage0_3[20]},
      {stage1_4[20],stage1_3[34],stage1_2[34],stage1_1[34],stage1_0[34]}
   );
   gpc1163_5 gpc35 (
      {stage0_0[161], stage0_0[162], stage0_0[163]},
      {stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143], stage0_1[144], stage0_1[145]},
      {stage0_2[35]},
      {stage0_3[21]},
      {stage1_4[21],stage1_3[35],stage1_2[35],stage1_1[35],stage1_0[35]}
   );
   gpc1163_5 gpc36 (
      {stage0_0[164], stage0_0[165], stage0_0[166]},
      {stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149], stage0_1[150], stage0_1[151]},
      {stage0_2[36]},
      {stage0_3[22]},
      {stage1_4[22],stage1_3[36],stage1_2[36],stage1_1[36],stage1_0[36]}
   );
   gpc1163_5 gpc37 (
      {stage0_0[167], stage0_0[168], stage0_0[169]},
      {stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155], stage0_1[156], stage0_1[157]},
      {stage0_2[37]},
      {stage0_3[23]},
      {stage1_4[23],stage1_3[37],stage1_2[37],stage1_1[37],stage1_0[37]}
   );
   gpc1163_5 gpc38 (
      {stage0_0[170], stage0_0[171], stage0_0[172]},
      {stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161], stage0_1[162], stage0_1[163]},
      {stage0_2[38]},
      {stage0_3[24]},
      {stage1_4[24],stage1_3[38],stage1_2[38],stage1_1[38],stage1_0[38]}
   );
   gpc1163_5 gpc39 (
      {stage0_0[173], stage0_0[174], stage0_0[175]},
      {stage0_1[164], stage0_1[165], stage0_1[166], stage0_1[167], stage0_1[168], stage0_1[169]},
      {stage0_2[39]},
      {stage0_3[25]},
      {stage1_4[25],stage1_3[39],stage1_2[39],stage1_1[39],stage1_0[39]}
   );
   gpc1163_5 gpc40 (
      {stage0_0[176], stage0_0[177], stage0_0[178]},
      {stage0_1[170], stage0_1[171], stage0_1[172], stage0_1[173], stage0_1[174], stage0_1[175]},
      {stage0_2[40]},
      {stage0_3[26]},
      {stage1_4[26],stage1_3[40],stage1_2[40],stage1_1[40],stage1_0[40]}
   );
   gpc1163_5 gpc41 (
      {stage0_0[179], stage0_0[180], stage0_0[181]},
      {stage0_1[176], stage0_1[177], stage0_1[178], stage0_1[179], stage0_1[180], stage0_1[181]},
      {stage0_2[41]},
      {stage0_3[27]},
      {stage1_4[27],stage1_3[41],stage1_2[41],stage1_1[41],stage1_0[41]}
   );
   gpc1163_5 gpc42 (
      {stage0_0[182], stage0_0[183], stage0_0[184]},
      {stage0_1[182], stage0_1[183], stage0_1[184], stage0_1[185], stage0_1[186], stage0_1[187]},
      {stage0_2[42]},
      {stage0_3[28]},
      {stage1_4[28],stage1_3[42],stage1_2[42],stage1_1[42],stage1_0[42]}
   );
   gpc1163_5 gpc43 (
      {stage0_0[185], stage0_0[186], stage0_0[187]},
      {stage0_1[188], stage0_1[189], stage0_1[190], stage0_1[191], stage0_1[192], stage0_1[193]},
      {stage0_2[43]},
      {stage0_3[29]},
      {stage1_4[29],stage1_3[43],stage1_2[43],stage1_1[43],stage1_0[43]}
   );
   gpc1163_5 gpc44 (
      {stage0_0[188], stage0_0[189], stage0_0[190]},
      {stage0_1[194], stage0_1[195], stage0_1[196], stage0_1[197], stage0_1[198], stage0_1[199]},
      {stage0_2[44]},
      {stage0_3[30]},
      {stage1_4[30],stage1_3[44],stage1_2[44],stage1_1[44],stage1_0[44]}
   );
   gpc606_5 gpc45 (
      {stage0_0[191], stage0_0[192], stage0_0[193], stage0_0[194], stage0_0[195], stage0_0[196]},
      {stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49], stage0_2[50]},
      {stage1_4[31],stage1_3[45],stage1_2[45],stage1_1[45],stage1_0[45]}
   );
   gpc606_5 gpc46 (
      {stage0_0[197], stage0_0[198], stage0_0[199], stage0_0[200], stage0_0[201], stage0_0[202]},
      {stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55], stage0_2[56]},
      {stage1_4[32],stage1_3[46],stage1_2[46],stage1_1[46],stage1_0[46]}
   );
   gpc606_5 gpc47 (
      {stage0_0[203], stage0_0[204], stage0_0[205], stage0_0[206], stage0_0[207], stage0_0[208]},
      {stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61], stage0_2[62]},
      {stage1_4[33],stage1_3[47],stage1_2[47],stage1_1[47],stage1_0[47]}
   );
   gpc606_5 gpc48 (
      {stage0_0[209], stage0_0[210], stage0_0[211], stage0_0[212], stage0_0[213], stage0_0[214]},
      {stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67], stage0_2[68]},
      {stage1_4[34],stage1_3[48],stage1_2[48],stage1_1[48],stage1_0[48]}
   );
   gpc606_5 gpc49 (
      {stage0_0[215], stage0_0[216], stage0_0[217], stage0_0[218], stage0_0[219], stage0_0[220]},
      {stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73], stage0_2[74]},
      {stage1_4[35],stage1_3[49],stage1_2[49],stage1_1[49],stage1_0[49]}
   );
   gpc606_5 gpc50 (
      {stage0_0[221], stage0_0[222], stage0_0[223], stage0_0[224], stage0_0[225], stage0_0[226]},
      {stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79], stage0_2[80]},
      {stage1_4[36],stage1_3[50],stage1_2[50],stage1_1[50],stage1_0[50]}
   );
   gpc606_5 gpc51 (
      {stage0_0[227], stage0_0[228], stage0_0[229], stage0_0[230], stage0_0[231], stage0_0[232]},
      {stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85], stage0_2[86]},
      {stage1_4[37],stage1_3[51],stage1_2[51],stage1_1[51],stage1_0[51]}
   );
   gpc606_5 gpc52 (
      {stage0_0[233], stage0_0[234], stage0_0[235], stage0_0[236], stage0_0[237], stage0_0[238]},
      {stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91], stage0_2[92]},
      {stage1_4[38],stage1_3[52],stage1_2[52],stage1_1[52],stage1_0[52]}
   );
   gpc606_5 gpc53 (
      {stage0_0[239], stage0_0[240], stage0_0[241], stage0_0[242], stage0_0[243], stage0_0[244]},
      {stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97], stage0_2[98]},
      {stage1_4[39],stage1_3[53],stage1_2[53],stage1_1[53],stage1_0[53]}
   );
   gpc606_5 gpc54 (
      {stage0_0[245], stage0_0[246], stage0_0[247], stage0_0[248], stage0_0[249], stage0_0[250]},
      {stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103], stage0_2[104]},
      {stage1_4[40],stage1_3[54],stage1_2[54],stage1_1[54],stage1_0[54]}
   );
   gpc606_5 gpc55 (
      {stage0_0[251], stage0_0[252], stage0_0[253], stage0_0[254], stage0_0[255], stage0_0[256]},
      {stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109], stage0_2[110]},
      {stage1_4[41],stage1_3[55],stage1_2[55],stage1_1[55],stage1_0[55]}
   );
   gpc606_5 gpc56 (
      {stage0_0[257], stage0_0[258], stage0_0[259], stage0_0[260], stage0_0[261], stage0_0[262]},
      {stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115], stage0_2[116]},
      {stage1_4[42],stage1_3[56],stage1_2[56],stage1_1[56],stage1_0[56]}
   );
   gpc606_5 gpc57 (
      {stage0_0[263], stage0_0[264], stage0_0[265], stage0_0[266], stage0_0[267], stage0_0[268]},
      {stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121], stage0_2[122]},
      {stage1_4[43],stage1_3[57],stage1_2[57],stage1_1[57],stage1_0[57]}
   );
   gpc606_5 gpc58 (
      {stage0_0[269], stage0_0[270], stage0_0[271], stage0_0[272], stage0_0[273], stage0_0[274]},
      {stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127], stage0_2[128]},
      {stage1_4[44],stage1_3[58],stage1_2[58],stage1_1[58],stage1_0[58]}
   );
   gpc606_5 gpc59 (
      {stage0_0[275], stage0_0[276], stage0_0[277], stage0_0[278], stage0_0[279], stage0_0[280]},
      {stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133], stage0_2[134]},
      {stage1_4[45],stage1_3[59],stage1_2[59],stage1_1[59],stage1_0[59]}
   );
   gpc606_5 gpc60 (
      {stage0_0[281], stage0_0[282], stage0_0[283], stage0_0[284], stage0_0[285], stage0_0[286]},
      {stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139], stage0_2[140]},
      {stage1_4[46],stage1_3[60],stage1_2[60],stage1_1[60],stage1_0[60]}
   );
   gpc606_5 gpc61 (
      {stage0_0[287], stage0_0[288], stage0_0[289], stage0_0[290], stage0_0[291], stage0_0[292]},
      {stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145], stage0_2[146]},
      {stage1_4[47],stage1_3[61],stage1_2[61],stage1_1[61],stage1_0[61]}
   );
   gpc606_5 gpc62 (
      {stage0_0[293], stage0_0[294], stage0_0[295], stage0_0[296], stage0_0[297], stage0_0[298]},
      {stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151], stage0_2[152]},
      {stage1_4[48],stage1_3[62],stage1_2[62],stage1_1[62],stage1_0[62]}
   );
   gpc606_5 gpc63 (
      {stage0_0[299], stage0_0[300], stage0_0[301], stage0_0[302], stage0_0[303], stage0_0[304]},
      {stage0_2[153], stage0_2[154], stage0_2[155], stage0_2[156], stage0_2[157], stage0_2[158]},
      {stage1_4[49],stage1_3[63],stage1_2[63],stage1_1[63],stage1_0[63]}
   );
   gpc606_5 gpc64 (
      {stage0_0[305], stage0_0[306], stage0_0[307], stage0_0[308], stage0_0[309], stage0_0[310]},
      {stage0_2[159], stage0_2[160], stage0_2[161], stage0_2[162], stage0_2[163], stage0_2[164]},
      {stage1_4[50],stage1_3[64],stage1_2[64],stage1_1[64],stage1_0[64]}
   );
   gpc606_5 gpc65 (
      {stage0_0[311], stage0_0[312], stage0_0[313], stage0_0[314], stage0_0[315], stage0_0[316]},
      {stage0_2[165], stage0_2[166], stage0_2[167], stage0_2[168], stage0_2[169], stage0_2[170]},
      {stage1_4[51],stage1_3[65],stage1_2[65],stage1_1[65],stage1_0[65]}
   );
   gpc606_5 gpc66 (
      {stage0_0[317], stage0_0[318], stage0_0[319], stage0_0[320], stage0_0[321], stage0_0[322]},
      {stage0_2[171], stage0_2[172], stage0_2[173], stage0_2[174], stage0_2[175], stage0_2[176]},
      {stage1_4[52],stage1_3[66],stage1_2[66],stage1_1[66],stage1_0[66]}
   );
   gpc606_5 gpc67 (
      {stage0_0[323], stage0_0[324], stage0_0[325], stage0_0[326], stage0_0[327], stage0_0[328]},
      {stage0_2[177], stage0_2[178], stage0_2[179], stage0_2[180], stage0_2[181], stage0_2[182]},
      {stage1_4[53],stage1_3[67],stage1_2[67],stage1_1[67],stage1_0[67]}
   );
   gpc606_5 gpc68 (
      {stage0_0[329], stage0_0[330], stage0_0[331], stage0_0[332], stage0_0[333], stage0_0[334]},
      {stage0_2[183], stage0_2[184], stage0_2[185], stage0_2[186], stage0_2[187], stage0_2[188]},
      {stage1_4[54],stage1_3[68],stage1_2[68],stage1_1[68],stage1_0[68]}
   );
   gpc606_5 gpc69 (
      {stage0_0[335], stage0_0[336], stage0_0[337], stage0_0[338], stage0_0[339], stage0_0[340]},
      {stage0_2[189], stage0_2[190], stage0_2[191], stage0_2[192], stage0_2[193], stage0_2[194]},
      {stage1_4[55],stage1_3[69],stage1_2[69],stage1_1[69],stage1_0[69]}
   );
   gpc606_5 gpc70 (
      {stage0_0[341], stage0_0[342], stage0_0[343], stage0_0[344], stage0_0[345], stage0_0[346]},
      {stage0_2[195], stage0_2[196], stage0_2[197], stage0_2[198], stage0_2[199], stage0_2[200]},
      {stage1_4[56],stage1_3[70],stage1_2[70],stage1_1[70],stage1_0[70]}
   );
   gpc606_5 gpc71 (
      {stage0_0[347], stage0_0[348], stage0_0[349], stage0_0[350], stage0_0[351], stage0_0[352]},
      {stage0_2[201], stage0_2[202], stage0_2[203], stage0_2[204], stage0_2[205], stage0_2[206]},
      {stage1_4[57],stage1_3[71],stage1_2[71],stage1_1[71],stage1_0[71]}
   );
   gpc606_5 gpc72 (
      {stage0_0[353], stage0_0[354], stage0_0[355], stage0_0[356], stage0_0[357], stage0_0[358]},
      {stage0_2[207], stage0_2[208], stage0_2[209], stage0_2[210], stage0_2[211], stage0_2[212]},
      {stage1_4[58],stage1_3[72],stage1_2[72],stage1_1[72],stage1_0[72]}
   );
   gpc606_5 gpc73 (
      {stage0_0[359], stage0_0[360], stage0_0[361], stage0_0[362], stage0_0[363], stage0_0[364]},
      {stage0_2[213], stage0_2[214], stage0_2[215], stage0_2[216], stage0_2[217], stage0_2[218]},
      {stage1_4[59],stage1_3[73],stage1_2[73],stage1_1[73],stage1_0[73]}
   );
   gpc606_5 gpc74 (
      {stage0_0[365], stage0_0[366], stage0_0[367], stage0_0[368], stage0_0[369], stage0_0[370]},
      {stage0_2[219], stage0_2[220], stage0_2[221], stage0_2[222], stage0_2[223], stage0_2[224]},
      {stage1_4[60],stage1_3[74],stage1_2[74],stage1_1[74],stage1_0[74]}
   );
   gpc606_5 gpc75 (
      {stage0_0[371], stage0_0[372], stage0_0[373], stage0_0[374], stage0_0[375], stage0_0[376]},
      {stage0_2[225], stage0_2[226], stage0_2[227], stage0_2[228], stage0_2[229], stage0_2[230]},
      {stage1_4[61],stage1_3[75],stage1_2[75],stage1_1[75],stage1_0[75]}
   );
   gpc606_5 gpc76 (
      {stage0_0[377], stage0_0[378], stage0_0[379], stage0_0[380], stage0_0[381], stage0_0[382]},
      {stage0_2[231], stage0_2[232], stage0_2[233], stage0_2[234], stage0_2[235], stage0_2[236]},
      {stage1_4[62],stage1_3[76],stage1_2[76],stage1_1[76],stage1_0[76]}
   );
   gpc606_5 gpc77 (
      {stage0_0[383], stage0_0[384], stage0_0[385], stage0_0[386], stage0_0[387], stage0_0[388]},
      {stage0_2[237], stage0_2[238], stage0_2[239], stage0_2[240], stage0_2[241], stage0_2[242]},
      {stage1_4[63],stage1_3[77],stage1_2[77],stage1_1[77],stage1_0[77]}
   );
   gpc606_5 gpc78 (
      {stage0_0[389], stage0_0[390], stage0_0[391], stage0_0[392], stage0_0[393], stage0_0[394]},
      {stage0_2[243], stage0_2[244], stage0_2[245], stage0_2[246], stage0_2[247], stage0_2[248]},
      {stage1_4[64],stage1_3[78],stage1_2[78],stage1_1[78],stage1_0[78]}
   );
   gpc606_5 gpc79 (
      {stage0_0[395], stage0_0[396], stage0_0[397], stage0_0[398], stage0_0[399], stage0_0[400]},
      {stage0_2[249], stage0_2[250], stage0_2[251], stage0_2[252], stage0_2[253], stage0_2[254]},
      {stage1_4[65],stage1_3[79],stage1_2[79],stage1_1[79],stage1_0[79]}
   );
   gpc606_5 gpc80 (
      {stage0_0[401], stage0_0[402], stage0_0[403], stage0_0[404], stage0_0[405], stage0_0[406]},
      {stage0_2[255], stage0_2[256], stage0_2[257], stage0_2[258], stage0_2[259], stage0_2[260]},
      {stage1_4[66],stage1_3[80],stage1_2[80],stage1_1[80],stage1_0[80]}
   );
   gpc606_5 gpc81 (
      {stage0_0[407], stage0_0[408], stage0_0[409], stage0_0[410], stage0_0[411], stage0_0[412]},
      {stage0_2[261], stage0_2[262], stage0_2[263], stage0_2[264], stage0_2[265], stage0_2[266]},
      {stage1_4[67],stage1_3[81],stage1_2[81],stage1_1[81],stage1_0[81]}
   );
   gpc606_5 gpc82 (
      {stage0_0[413], stage0_0[414], stage0_0[415], stage0_0[416], stage0_0[417], stage0_0[418]},
      {stage0_2[267], stage0_2[268], stage0_2[269], stage0_2[270], stage0_2[271], stage0_2[272]},
      {stage1_4[68],stage1_3[82],stage1_2[82],stage1_1[82],stage1_0[82]}
   );
   gpc606_5 gpc83 (
      {stage0_0[419], stage0_0[420], stage0_0[421], stage0_0[422], stage0_0[423], stage0_0[424]},
      {stage0_2[273], stage0_2[274], stage0_2[275], stage0_2[276], stage0_2[277], stage0_2[278]},
      {stage1_4[69],stage1_3[83],stage1_2[83],stage1_1[83],stage1_0[83]}
   );
   gpc606_5 gpc84 (
      {stage0_0[425], stage0_0[426], stage0_0[427], stage0_0[428], stage0_0[429], stage0_0[430]},
      {stage0_2[279], stage0_2[280], stage0_2[281], stage0_2[282], stage0_2[283], stage0_2[284]},
      {stage1_4[70],stage1_3[84],stage1_2[84],stage1_1[84],stage1_0[84]}
   );
   gpc606_5 gpc85 (
      {stage0_0[431], stage0_0[432], stage0_0[433], stage0_0[434], stage0_0[435], stage0_0[436]},
      {stage0_2[285], stage0_2[286], stage0_2[287], stage0_2[288], stage0_2[289], stage0_2[290]},
      {stage1_4[71],stage1_3[85],stage1_2[85],stage1_1[85],stage1_0[85]}
   );
   gpc606_5 gpc86 (
      {stage0_0[437], stage0_0[438], stage0_0[439], stage0_0[440], stage0_0[441], stage0_0[442]},
      {stage0_2[291], stage0_2[292], stage0_2[293], stage0_2[294], stage0_2[295], stage0_2[296]},
      {stage1_4[72],stage1_3[86],stage1_2[86],stage1_1[86],stage1_0[86]}
   );
   gpc606_5 gpc87 (
      {stage0_0[443], stage0_0[444], stage0_0[445], stage0_0[446], stage0_0[447], stage0_0[448]},
      {stage0_2[297], stage0_2[298], stage0_2[299], stage0_2[300], stage0_2[301], stage0_2[302]},
      {stage1_4[73],stage1_3[87],stage1_2[87],stage1_1[87],stage1_0[87]}
   );
   gpc606_5 gpc88 (
      {stage0_0[449], stage0_0[450], stage0_0[451], stage0_0[452], stage0_0[453], stage0_0[454]},
      {stage0_2[303], stage0_2[304], stage0_2[305], stage0_2[306], stage0_2[307], stage0_2[308]},
      {stage1_4[74],stage1_3[88],stage1_2[88],stage1_1[88],stage1_0[88]}
   );
   gpc606_5 gpc89 (
      {stage0_0[455], stage0_0[456], stage0_0[457], stage0_0[458], stage0_0[459], stage0_0[460]},
      {stage0_2[309], stage0_2[310], stage0_2[311], stage0_2[312], stage0_2[313], stage0_2[314]},
      {stage1_4[75],stage1_3[89],stage1_2[89],stage1_1[89],stage1_0[89]}
   );
   gpc606_5 gpc90 (
      {stage0_0[461], stage0_0[462], stage0_0[463], stage0_0[464], stage0_0[465], stage0_0[466]},
      {stage0_2[315], stage0_2[316], stage0_2[317], stage0_2[318], stage0_2[319], stage0_2[320]},
      {stage1_4[76],stage1_3[90],stage1_2[90],stage1_1[90],stage1_0[90]}
   );
   gpc606_5 gpc91 (
      {stage0_0[467], stage0_0[468], stage0_0[469], stage0_0[470], stage0_0[471], stage0_0[472]},
      {stage0_2[321], stage0_2[322], stage0_2[323], stage0_2[324], stage0_2[325], stage0_2[326]},
      {stage1_4[77],stage1_3[91],stage1_2[91],stage1_1[91],stage1_0[91]}
   );
   gpc606_5 gpc92 (
      {stage0_0[473], stage0_0[474], stage0_0[475], stage0_0[476], stage0_0[477], stage0_0[478]},
      {stage0_2[327], stage0_2[328], stage0_2[329], stage0_2[330], stage0_2[331], stage0_2[332]},
      {stage1_4[78],stage1_3[92],stage1_2[92],stage1_1[92],stage1_0[92]}
   );
   gpc606_5 gpc93 (
      {stage0_0[479], stage0_0[480], stage0_0[481], stage0_0[482], stage0_0[483], stage0_0[484]},
      {stage0_2[333], stage0_2[334], stage0_2[335], stage0_2[336], stage0_2[337], stage0_2[338]},
      {stage1_4[79],stage1_3[93],stage1_2[93],stage1_1[93],stage1_0[93]}
   );
   gpc606_5 gpc94 (
      {stage0_0[485], stage0_0[486], stage0_0[487], stage0_0[488], stage0_0[489], stage0_0[490]},
      {stage0_2[339], stage0_2[340], stage0_2[341], stage0_2[342], stage0_2[343], stage0_2[344]},
      {stage1_4[80],stage1_3[94],stage1_2[94],stage1_1[94],stage1_0[94]}
   );
   gpc606_5 gpc95 (
      {stage0_0[491], stage0_0[492], stage0_0[493], stage0_0[494], stage0_0[495], stage0_0[496]},
      {stage0_2[345], stage0_2[346], stage0_2[347], stage0_2[348], stage0_2[349], stage0_2[350]},
      {stage1_4[81],stage1_3[95],stage1_2[95],stage1_1[95],stage1_0[95]}
   );
   gpc606_5 gpc96 (
      {stage0_0[497], stage0_0[498], stage0_0[499], stage0_0[500], stage0_0[501], stage0_0[502]},
      {stage0_2[351], stage0_2[352], stage0_2[353], stage0_2[354], stage0_2[355], stage0_2[356]},
      {stage1_4[82],stage1_3[96],stage1_2[96],stage1_1[96],stage1_0[96]}
   );
   gpc606_5 gpc97 (
      {stage0_0[503], stage0_0[504], stage0_0[505], stage0_0[506], stage0_0[507], stage0_0[508]},
      {stage0_2[357], stage0_2[358], stage0_2[359], stage0_2[360], stage0_2[361], stage0_2[362]},
      {stage1_4[83],stage1_3[97],stage1_2[97],stage1_1[97],stage1_0[97]}
   );
   gpc606_5 gpc98 (
      {stage0_1[200], stage0_1[201], stage0_1[202], stage0_1[203], stage0_1[204], stage0_1[205]},
      {stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36]},
      {stage1_5[0],stage1_4[84],stage1_3[98],stage1_2[98],stage1_1[98]}
   );
   gpc606_5 gpc99 (
      {stage0_1[206], stage0_1[207], stage0_1[208], stage0_1[209], stage0_1[210], stage0_1[211]},
      {stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42]},
      {stage1_5[1],stage1_4[85],stage1_3[99],stage1_2[99],stage1_1[99]}
   );
   gpc606_5 gpc100 (
      {stage0_1[212], stage0_1[213], stage0_1[214], stage0_1[215], stage0_1[216], stage0_1[217]},
      {stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48]},
      {stage1_5[2],stage1_4[86],stage1_3[100],stage1_2[100],stage1_1[100]}
   );
   gpc606_5 gpc101 (
      {stage0_1[218], stage0_1[219], stage0_1[220], stage0_1[221], stage0_1[222], stage0_1[223]},
      {stage0_3[49], stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54]},
      {stage1_5[3],stage1_4[87],stage1_3[101],stage1_2[101],stage1_1[101]}
   );
   gpc606_5 gpc102 (
      {stage0_1[224], stage0_1[225], stage0_1[226], stage0_1[227], stage0_1[228], stage0_1[229]},
      {stage0_3[55], stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60]},
      {stage1_5[4],stage1_4[88],stage1_3[102],stage1_2[102],stage1_1[102]}
   );
   gpc606_5 gpc103 (
      {stage0_1[230], stage0_1[231], stage0_1[232], stage0_1[233], stage0_1[234], stage0_1[235]},
      {stage0_3[61], stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66]},
      {stage1_5[5],stage1_4[89],stage1_3[103],stage1_2[103],stage1_1[103]}
   );
   gpc606_5 gpc104 (
      {stage0_1[236], stage0_1[237], stage0_1[238], stage0_1[239], stage0_1[240], stage0_1[241]},
      {stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72]},
      {stage1_5[6],stage1_4[90],stage1_3[104],stage1_2[104],stage1_1[104]}
   );
   gpc606_5 gpc105 (
      {stage0_1[242], stage0_1[243], stage0_1[244], stage0_1[245], stage0_1[246], stage0_1[247]},
      {stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78]},
      {stage1_5[7],stage1_4[91],stage1_3[105],stage1_2[105],stage1_1[105]}
   );
   gpc606_5 gpc106 (
      {stage0_1[248], stage0_1[249], stage0_1[250], stage0_1[251], stage0_1[252], stage0_1[253]},
      {stage0_3[79], stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83], stage0_3[84]},
      {stage1_5[8],stage1_4[92],stage1_3[106],stage1_2[106],stage1_1[106]}
   );
   gpc606_5 gpc107 (
      {stage0_1[254], stage0_1[255], stage0_1[256], stage0_1[257], stage0_1[258], stage0_1[259]},
      {stage0_3[85], stage0_3[86], stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90]},
      {stage1_5[9],stage1_4[93],stage1_3[107],stage1_2[107],stage1_1[107]}
   );
   gpc606_5 gpc108 (
      {stage0_1[260], stage0_1[261], stage0_1[262], stage0_1[263], stage0_1[264], stage0_1[265]},
      {stage0_3[91], stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96]},
      {stage1_5[10],stage1_4[94],stage1_3[108],stage1_2[108],stage1_1[108]}
   );
   gpc606_5 gpc109 (
      {stage0_1[266], stage0_1[267], stage0_1[268], stage0_1[269], stage0_1[270], stage0_1[271]},
      {stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101], stage0_3[102]},
      {stage1_5[11],stage1_4[95],stage1_3[109],stage1_2[109],stage1_1[109]}
   );
   gpc606_5 gpc110 (
      {stage0_1[272], stage0_1[273], stage0_1[274], stage0_1[275], stage0_1[276], stage0_1[277]},
      {stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106], stage0_3[107], stage0_3[108]},
      {stage1_5[12],stage1_4[96],stage1_3[110],stage1_2[110],stage1_1[110]}
   );
   gpc606_5 gpc111 (
      {stage0_1[278], stage0_1[279], stage0_1[280], stage0_1[281], stage0_1[282], stage0_1[283]},
      {stage0_3[109], stage0_3[110], stage0_3[111], stage0_3[112], stage0_3[113], stage0_3[114]},
      {stage1_5[13],stage1_4[97],stage1_3[111],stage1_2[111],stage1_1[111]}
   );
   gpc606_5 gpc112 (
      {stage0_1[284], stage0_1[285], stage0_1[286], stage0_1[287], stage0_1[288], stage0_1[289]},
      {stage0_3[115], stage0_3[116], stage0_3[117], stage0_3[118], stage0_3[119], stage0_3[120]},
      {stage1_5[14],stage1_4[98],stage1_3[112],stage1_2[112],stage1_1[112]}
   );
   gpc606_5 gpc113 (
      {stage0_1[290], stage0_1[291], stage0_1[292], stage0_1[293], stage0_1[294], stage0_1[295]},
      {stage0_3[121], stage0_3[122], stage0_3[123], stage0_3[124], stage0_3[125], stage0_3[126]},
      {stage1_5[15],stage1_4[99],stage1_3[113],stage1_2[113],stage1_1[113]}
   );
   gpc606_5 gpc114 (
      {stage0_1[296], stage0_1[297], stage0_1[298], stage0_1[299], stage0_1[300], stage0_1[301]},
      {stage0_3[127], stage0_3[128], stage0_3[129], stage0_3[130], stage0_3[131], stage0_3[132]},
      {stage1_5[16],stage1_4[100],stage1_3[114],stage1_2[114],stage1_1[114]}
   );
   gpc606_5 gpc115 (
      {stage0_1[302], stage0_1[303], stage0_1[304], stage0_1[305], stage0_1[306], stage0_1[307]},
      {stage0_3[133], stage0_3[134], stage0_3[135], stage0_3[136], stage0_3[137], stage0_3[138]},
      {stage1_5[17],stage1_4[101],stage1_3[115],stage1_2[115],stage1_1[115]}
   );
   gpc606_5 gpc116 (
      {stage0_1[308], stage0_1[309], stage0_1[310], stage0_1[311], stage0_1[312], stage0_1[313]},
      {stage0_3[139], stage0_3[140], stage0_3[141], stage0_3[142], stage0_3[143], stage0_3[144]},
      {stage1_5[18],stage1_4[102],stage1_3[116],stage1_2[116],stage1_1[116]}
   );
   gpc606_5 gpc117 (
      {stage0_1[314], stage0_1[315], stage0_1[316], stage0_1[317], stage0_1[318], stage0_1[319]},
      {stage0_3[145], stage0_3[146], stage0_3[147], stage0_3[148], stage0_3[149], stage0_3[150]},
      {stage1_5[19],stage1_4[103],stage1_3[117],stage1_2[117],stage1_1[117]}
   );
   gpc606_5 gpc118 (
      {stage0_1[320], stage0_1[321], stage0_1[322], stage0_1[323], stage0_1[324], stage0_1[325]},
      {stage0_3[151], stage0_3[152], stage0_3[153], stage0_3[154], stage0_3[155], stage0_3[156]},
      {stage1_5[20],stage1_4[104],stage1_3[118],stage1_2[118],stage1_1[118]}
   );
   gpc606_5 gpc119 (
      {stage0_1[326], stage0_1[327], stage0_1[328], stage0_1[329], stage0_1[330], stage0_1[331]},
      {stage0_3[157], stage0_3[158], stage0_3[159], stage0_3[160], stage0_3[161], stage0_3[162]},
      {stage1_5[21],stage1_4[105],stage1_3[119],stage1_2[119],stage1_1[119]}
   );
   gpc606_5 gpc120 (
      {stage0_1[332], stage0_1[333], stage0_1[334], stage0_1[335], stage0_1[336], stage0_1[337]},
      {stage0_3[163], stage0_3[164], stage0_3[165], stage0_3[166], stage0_3[167], stage0_3[168]},
      {stage1_5[22],stage1_4[106],stage1_3[120],stage1_2[120],stage1_1[120]}
   );
   gpc606_5 gpc121 (
      {stage0_1[338], stage0_1[339], stage0_1[340], stage0_1[341], stage0_1[342], stage0_1[343]},
      {stage0_3[169], stage0_3[170], stage0_3[171], stage0_3[172], stage0_3[173], stage0_3[174]},
      {stage1_5[23],stage1_4[107],stage1_3[121],stage1_2[121],stage1_1[121]}
   );
   gpc606_5 gpc122 (
      {stage0_1[344], stage0_1[345], stage0_1[346], stage0_1[347], stage0_1[348], stage0_1[349]},
      {stage0_3[175], stage0_3[176], stage0_3[177], stage0_3[178], stage0_3[179], stage0_3[180]},
      {stage1_5[24],stage1_4[108],stage1_3[122],stage1_2[122],stage1_1[122]}
   );
   gpc606_5 gpc123 (
      {stage0_1[350], stage0_1[351], stage0_1[352], stage0_1[353], stage0_1[354], stage0_1[355]},
      {stage0_3[181], stage0_3[182], stage0_3[183], stage0_3[184], stage0_3[185], stage0_3[186]},
      {stage1_5[25],stage1_4[109],stage1_3[123],stage1_2[123],stage1_1[123]}
   );
   gpc606_5 gpc124 (
      {stage0_1[356], stage0_1[357], stage0_1[358], stage0_1[359], stage0_1[360], stage0_1[361]},
      {stage0_3[187], stage0_3[188], stage0_3[189], stage0_3[190], stage0_3[191], stage0_3[192]},
      {stage1_5[26],stage1_4[110],stage1_3[124],stage1_2[124],stage1_1[124]}
   );
   gpc606_5 gpc125 (
      {stage0_1[362], stage0_1[363], stage0_1[364], stage0_1[365], stage0_1[366], stage0_1[367]},
      {stage0_3[193], stage0_3[194], stage0_3[195], stage0_3[196], stage0_3[197], stage0_3[198]},
      {stage1_5[27],stage1_4[111],stage1_3[125],stage1_2[125],stage1_1[125]}
   );
   gpc606_5 gpc126 (
      {stage0_1[368], stage0_1[369], stage0_1[370], stage0_1[371], stage0_1[372], stage0_1[373]},
      {stage0_3[199], stage0_3[200], stage0_3[201], stage0_3[202], stage0_3[203], stage0_3[204]},
      {stage1_5[28],stage1_4[112],stage1_3[126],stage1_2[126],stage1_1[126]}
   );
   gpc606_5 gpc127 (
      {stage0_1[374], stage0_1[375], stage0_1[376], stage0_1[377], stage0_1[378], stage0_1[379]},
      {stage0_3[205], stage0_3[206], stage0_3[207], stage0_3[208], stage0_3[209], stage0_3[210]},
      {stage1_5[29],stage1_4[113],stage1_3[127],stage1_2[127],stage1_1[127]}
   );
   gpc606_5 gpc128 (
      {stage0_1[380], stage0_1[381], stage0_1[382], stage0_1[383], stage0_1[384], stage0_1[385]},
      {stage0_3[211], stage0_3[212], stage0_3[213], stage0_3[214], stage0_3[215], stage0_3[216]},
      {stage1_5[30],stage1_4[114],stage1_3[128],stage1_2[128],stage1_1[128]}
   );
   gpc606_5 gpc129 (
      {stage0_1[386], stage0_1[387], stage0_1[388], stage0_1[389], stage0_1[390], stage0_1[391]},
      {stage0_3[217], stage0_3[218], stage0_3[219], stage0_3[220], stage0_3[221], stage0_3[222]},
      {stage1_5[31],stage1_4[115],stage1_3[129],stage1_2[129],stage1_1[129]}
   );
   gpc606_5 gpc130 (
      {stage0_1[392], stage0_1[393], stage0_1[394], stage0_1[395], stage0_1[396], stage0_1[397]},
      {stage0_3[223], stage0_3[224], stage0_3[225], stage0_3[226], stage0_3[227], stage0_3[228]},
      {stage1_5[32],stage1_4[116],stage1_3[130],stage1_2[130],stage1_1[130]}
   );
   gpc606_5 gpc131 (
      {stage0_1[398], stage0_1[399], stage0_1[400], stage0_1[401], stage0_1[402], stage0_1[403]},
      {stage0_3[229], stage0_3[230], stage0_3[231], stage0_3[232], stage0_3[233], stage0_3[234]},
      {stage1_5[33],stage1_4[117],stage1_3[131],stage1_2[131],stage1_1[131]}
   );
   gpc606_5 gpc132 (
      {stage0_1[404], stage0_1[405], stage0_1[406], stage0_1[407], stage0_1[408], stage0_1[409]},
      {stage0_3[235], stage0_3[236], stage0_3[237], stage0_3[238], stage0_3[239], stage0_3[240]},
      {stage1_5[34],stage1_4[118],stage1_3[132],stage1_2[132],stage1_1[132]}
   );
   gpc606_5 gpc133 (
      {stage0_1[410], stage0_1[411], stage0_1[412], stage0_1[413], stage0_1[414], stage0_1[415]},
      {stage0_3[241], stage0_3[242], stage0_3[243], stage0_3[244], stage0_3[245], stage0_3[246]},
      {stage1_5[35],stage1_4[119],stage1_3[133],stage1_2[133],stage1_1[133]}
   );
   gpc606_5 gpc134 (
      {stage0_1[416], stage0_1[417], stage0_1[418], stage0_1[419], stage0_1[420], stage0_1[421]},
      {stage0_3[247], stage0_3[248], stage0_3[249], stage0_3[250], stage0_3[251], stage0_3[252]},
      {stage1_5[36],stage1_4[120],stage1_3[134],stage1_2[134],stage1_1[134]}
   );
   gpc606_5 gpc135 (
      {stage0_1[422], stage0_1[423], stage0_1[424], stage0_1[425], stage0_1[426], stage0_1[427]},
      {stage0_3[253], stage0_3[254], stage0_3[255], stage0_3[256], stage0_3[257], stage0_3[258]},
      {stage1_5[37],stage1_4[121],stage1_3[135],stage1_2[135],stage1_1[135]}
   );
   gpc606_5 gpc136 (
      {stage0_1[428], stage0_1[429], stage0_1[430], stage0_1[431], stage0_1[432], stage0_1[433]},
      {stage0_3[259], stage0_3[260], stage0_3[261], stage0_3[262], stage0_3[263], stage0_3[264]},
      {stage1_5[38],stage1_4[122],stage1_3[136],stage1_2[136],stage1_1[136]}
   );
   gpc606_5 gpc137 (
      {stage0_1[434], stage0_1[435], stage0_1[436], stage0_1[437], stage0_1[438], stage0_1[439]},
      {stage0_3[265], stage0_3[266], stage0_3[267], stage0_3[268], stage0_3[269], stage0_3[270]},
      {stage1_5[39],stage1_4[123],stage1_3[137],stage1_2[137],stage1_1[137]}
   );
   gpc606_5 gpc138 (
      {stage0_1[440], stage0_1[441], stage0_1[442], stage0_1[443], stage0_1[444], stage0_1[445]},
      {stage0_3[271], stage0_3[272], stage0_3[273], stage0_3[274], stage0_3[275], stage0_3[276]},
      {stage1_5[40],stage1_4[124],stage1_3[138],stage1_2[138],stage1_1[138]}
   );
   gpc606_5 gpc139 (
      {stage0_1[446], stage0_1[447], stage0_1[448], stage0_1[449], stage0_1[450], stage0_1[451]},
      {stage0_3[277], stage0_3[278], stage0_3[279], stage0_3[280], stage0_3[281], stage0_3[282]},
      {stage1_5[41],stage1_4[125],stage1_3[139],stage1_2[139],stage1_1[139]}
   );
   gpc606_5 gpc140 (
      {stage0_1[452], stage0_1[453], stage0_1[454], stage0_1[455], stage0_1[456], stage0_1[457]},
      {stage0_3[283], stage0_3[284], stage0_3[285], stage0_3[286], stage0_3[287], stage0_3[288]},
      {stage1_5[42],stage1_4[126],stage1_3[140],stage1_2[140],stage1_1[140]}
   );
   gpc606_5 gpc141 (
      {stage0_1[458], stage0_1[459], stage0_1[460], stage0_1[461], stage0_1[462], stage0_1[463]},
      {stage0_3[289], stage0_3[290], stage0_3[291], stage0_3[292], stage0_3[293], stage0_3[294]},
      {stage1_5[43],stage1_4[127],stage1_3[141],stage1_2[141],stage1_1[141]}
   );
   gpc606_5 gpc142 (
      {stage0_1[464], stage0_1[465], stage0_1[466], stage0_1[467], stage0_1[468], stage0_1[469]},
      {stage0_3[295], stage0_3[296], stage0_3[297], stage0_3[298], stage0_3[299], stage0_3[300]},
      {stage1_5[44],stage1_4[128],stage1_3[142],stage1_2[142],stage1_1[142]}
   );
   gpc606_5 gpc143 (
      {stage0_1[470], stage0_1[471], stage0_1[472], stage0_1[473], stage0_1[474], stage0_1[475]},
      {stage0_3[301], stage0_3[302], stage0_3[303], stage0_3[304], stage0_3[305], stage0_3[306]},
      {stage1_5[45],stage1_4[129],stage1_3[143],stage1_2[143],stage1_1[143]}
   );
   gpc606_5 gpc144 (
      {stage0_2[363], stage0_2[364], stage0_2[365], stage0_2[366], stage0_2[367], stage0_2[368]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[46],stage1_4[130],stage1_3[144],stage1_2[144]}
   );
   gpc606_5 gpc145 (
      {stage0_2[369], stage0_2[370], stage0_2[371], stage0_2[372], stage0_2[373], stage0_2[374]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[47],stage1_4[131],stage1_3[145],stage1_2[145]}
   );
   gpc606_5 gpc146 (
      {stage0_2[375], stage0_2[376], stage0_2[377], stage0_2[378], stage0_2[379], stage0_2[380]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[48],stage1_4[132],stage1_3[146],stage1_2[146]}
   );
   gpc606_5 gpc147 (
      {stage0_2[381], stage0_2[382], stage0_2[383], stage0_2[384], stage0_2[385], stage0_2[386]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[49],stage1_4[133],stage1_3[147],stage1_2[147]}
   );
   gpc606_5 gpc148 (
      {stage0_2[387], stage0_2[388], stage0_2[389], stage0_2[390], stage0_2[391], stage0_2[392]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[50],stage1_4[134],stage1_3[148],stage1_2[148]}
   );
   gpc615_5 gpc149 (
      {stage0_2[393], stage0_2[394], stage0_2[395], stage0_2[396], stage0_2[397]},
      {stage0_3[307]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[51],stage1_4[135],stage1_3[149],stage1_2[149]}
   );
   gpc615_5 gpc150 (
      {stage0_2[398], stage0_2[399], stage0_2[400], stage0_2[401], stage0_2[402]},
      {stage0_3[308]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[52],stage1_4[136],stage1_3[150],stage1_2[150]}
   );
   gpc615_5 gpc151 (
      {stage0_2[403], stage0_2[404], stage0_2[405], stage0_2[406], stage0_2[407]},
      {stage0_3[309]},
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage1_6[7],stage1_5[53],stage1_4[137],stage1_3[151],stage1_2[151]}
   );
   gpc615_5 gpc152 (
      {stage0_2[408], stage0_2[409], stage0_2[410], stage0_2[411], stage0_2[412]},
      {stage0_3[310]},
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage1_6[8],stage1_5[54],stage1_4[138],stage1_3[152],stage1_2[152]}
   );
   gpc615_5 gpc153 (
      {stage0_2[413], stage0_2[414], stage0_2[415], stage0_2[416], stage0_2[417]},
      {stage0_3[311]},
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage1_6[9],stage1_5[55],stage1_4[139],stage1_3[153],stage1_2[153]}
   );
   gpc615_5 gpc154 (
      {stage0_2[418], stage0_2[419], stage0_2[420], stage0_2[421], stage0_2[422]},
      {stage0_3[312]},
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage1_6[10],stage1_5[56],stage1_4[140],stage1_3[154],stage1_2[154]}
   );
   gpc615_5 gpc155 (
      {stage0_2[423], stage0_2[424], stage0_2[425], stage0_2[426], stage0_2[427]},
      {stage0_3[313]},
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage1_6[11],stage1_5[57],stage1_4[141],stage1_3[155],stage1_2[155]}
   );
   gpc615_5 gpc156 (
      {stage0_2[428], stage0_2[429], stage0_2[430], stage0_2[431], stage0_2[432]},
      {stage0_3[314]},
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage1_6[12],stage1_5[58],stage1_4[142],stage1_3[156],stage1_2[156]}
   );
   gpc615_5 gpc157 (
      {stage0_2[433], stage0_2[434], stage0_2[435], stage0_2[436], stage0_2[437]},
      {stage0_3[315]},
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage1_6[13],stage1_5[59],stage1_4[143],stage1_3[157],stage1_2[157]}
   );
   gpc615_5 gpc158 (
      {stage0_2[438], stage0_2[439], stage0_2[440], stage0_2[441], stage0_2[442]},
      {stage0_3[316]},
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage1_6[14],stage1_5[60],stage1_4[144],stage1_3[158],stage1_2[158]}
   );
   gpc615_5 gpc159 (
      {stage0_2[443], stage0_2[444], stage0_2[445], stage0_2[446], stage0_2[447]},
      {stage0_3[317]},
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage1_6[15],stage1_5[61],stage1_4[145],stage1_3[159],stage1_2[159]}
   );
   gpc615_5 gpc160 (
      {stage0_2[448], stage0_2[449], stage0_2[450], stage0_2[451], stage0_2[452]},
      {stage0_3[318]},
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage1_6[16],stage1_5[62],stage1_4[146],stage1_3[160],stage1_2[160]}
   );
   gpc615_5 gpc161 (
      {stage0_2[453], stage0_2[454], stage0_2[455], stage0_2[456], stage0_2[457]},
      {stage0_3[319]},
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage1_6[17],stage1_5[63],stage1_4[147],stage1_3[161],stage1_2[161]}
   );
   gpc615_5 gpc162 (
      {stage0_2[458], stage0_2[459], stage0_2[460], stage0_2[461], stage0_2[462]},
      {stage0_3[320]},
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage1_6[18],stage1_5[64],stage1_4[148],stage1_3[162],stage1_2[162]}
   );
   gpc615_5 gpc163 (
      {stage0_2[463], stage0_2[464], stage0_2[465], stage0_2[466], stage0_2[467]},
      {stage0_3[321]},
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage1_6[19],stage1_5[65],stage1_4[149],stage1_3[163],stage1_2[163]}
   );
   gpc615_5 gpc164 (
      {stage0_2[468], stage0_2[469], stage0_2[470], stage0_2[471], stage0_2[472]},
      {stage0_3[322]},
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage1_6[20],stage1_5[66],stage1_4[150],stage1_3[164],stage1_2[164]}
   );
   gpc615_5 gpc165 (
      {stage0_2[473], stage0_2[474], stage0_2[475], stage0_2[476], stage0_2[477]},
      {stage0_3[323]},
      {stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131]},
      {stage1_6[21],stage1_5[67],stage1_4[151],stage1_3[165],stage1_2[165]}
   );
   gpc615_5 gpc166 (
      {stage0_2[478], stage0_2[479], stage0_2[480], stage0_2[481], stage0_2[482]},
      {stage0_3[324]},
      {stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137]},
      {stage1_6[22],stage1_5[68],stage1_4[152],stage1_3[166],stage1_2[166]}
   );
   gpc615_5 gpc167 (
      {stage0_2[483], stage0_2[484], stage0_2[485], stage0_2[486], stage0_2[487]},
      {stage0_3[325]},
      {stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143]},
      {stage1_6[23],stage1_5[69],stage1_4[153],stage1_3[167],stage1_2[167]}
   );
   gpc615_5 gpc168 (
      {stage0_2[488], stage0_2[489], stage0_2[490], stage0_2[491], stage0_2[492]},
      {stage0_3[326]},
      {stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149]},
      {stage1_6[24],stage1_5[70],stage1_4[154],stage1_3[168],stage1_2[168]}
   );
   gpc615_5 gpc169 (
      {stage0_2[493], stage0_2[494], stage0_2[495], stage0_2[496], stage0_2[497]},
      {stage0_3[327]},
      {stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155]},
      {stage1_6[25],stage1_5[71],stage1_4[155],stage1_3[169],stage1_2[169]}
   );
   gpc615_5 gpc170 (
      {stage0_2[498], stage0_2[499], stage0_2[500], stage0_2[501], stage0_2[502]},
      {stage0_3[328]},
      {stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161]},
      {stage1_6[26],stage1_5[72],stage1_4[156],stage1_3[170],stage1_2[170]}
   );
   gpc615_5 gpc171 (
      {stage0_2[503], stage0_2[504], stage0_2[505], stage0_2[506], stage0_2[507]},
      {stage0_3[329]},
      {stage0_4[162], stage0_4[163], stage0_4[164], stage0_4[165], stage0_4[166], stage0_4[167]},
      {stage1_6[27],stage1_5[73],stage1_4[157],stage1_3[171],stage1_2[171]}
   );
   gpc615_5 gpc172 (
      {stage0_2[508], stage0_2[509], stage0_2[510], stage0_2[511], 1'b0},
      {stage0_3[330]},
      {stage0_4[168], stage0_4[169], stage0_4[170], stage0_4[171], stage0_4[172], stage0_4[173]},
      {stage1_6[28],stage1_5[74],stage1_4[158],stage1_3[172],stage1_2[172]}
   );
   gpc615_5 gpc173 (
      {stage0_3[331], stage0_3[332], stage0_3[333], stage0_3[334], stage0_3[335]},
      {stage0_4[174]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[29],stage1_5[75],stage1_4[159],stage1_3[173]}
   );
   gpc615_5 gpc174 (
      {stage0_3[336], stage0_3[337], stage0_3[338], stage0_3[339], stage0_3[340]},
      {stage0_4[175]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[30],stage1_5[76],stage1_4[160],stage1_3[174]}
   );
   gpc615_5 gpc175 (
      {stage0_3[341], stage0_3[342], stage0_3[343], stage0_3[344], stage0_3[345]},
      {stage0_4[176]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[31],stage1_5[77],stage1_4[161],stage1_3[175]}
   );
   gpc615_5 gpc176 (
      {stage0_3[346], stage0_3[347], stage0_3[348], stage0_3[349], stage0_3[350]},
      {stage0_4[177]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[32],stage1_5[78],stage1_4[162],stage1_3[176]}
   );
   gpc615_5 gpc177 (
      {stage0_3[351], stage0_3[352], stage0_3[353], stage0_3[354], stage0_3[355]},
      {stage0_4[178]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[33],stage1_5[79],stage1_4[163],stage1_3[177]}
   );
   gpc615_5 gpc178 (
      {stage0_3[356], stage0_3[357], stage0_3[358], stage0_3[359], stage0_3[360]},
      {stage0_4[179]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[34],stage1_5[80],stage1_4[164],stage1_3[178]}
   );
   gpc615_5 gpc179 (
      {stage0_3[361], stage0_3[362], stage0_3[363], stage0_3[364], stage0_3[365]},
      {stage0_4[180]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[35],stage1_5[81],stage1_4[165],stage1_3[179]}
   );
   gpc615_5 gpc180 (
      {stage0_3[366], stage0_3[367], stage0_3[368], stage0_3[369], stage0_3[370]},
      {stage0_4[181]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[36],stage1_5[82],stage1_4[166],stage1_3[180]}
   );
   gpc615_5 gpc181 (
      {stage0_3[371], stage0_3[372], stage0_3[373], stage0_3[374], stage0_3[375]},
      {stage0_4[182]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[37],stage1_5[83],stage1_4[167],stage1_3[181]}
   );
   gpc615_5 gpc182 (
      {stage0_3[376], stage0_3[377], stage0_3[378], stage0_3[379], stage0_3[380]},
      {stage0_4[183]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[38],stage1_5[84],stage1_4[168],stage1_3[182]}
   );
   gpc615_5 gpc183 (
      {stage0_3[381], stage0_3[382], stage0_3[383], stage0_3[384], stage0_3[385]},
      {stage0_4[184]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[39],stage1_5[85],stage1_4[169],stage1_3[183]}
   );
   gpc615_5 gpc184 (
      {stage0_3[386], stage0_3[387], stage0_3[388], stage0_3[389], stage0_3[390]},
      {stage0_4[185]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[40],stage1_5[86],stage1_4[170],stage1_3[184]}
   );
   gpc615_5 gpc185 (
      {stage0_3[391], stage0_3[392], stage0_3[393], stage0_3[394], stage0_3[395]},
      {stage0_4[186]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[41],stage1_5[87],stage1_4[171],stage1_3[185]}
   );
   gpc615_5 gpc186 (
      {stage0_3[396], stage0_3[397], stage0_3[398], stage0_3[399], stage0_3[400]},
      {stage0_4[187]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[42],stage1_5[88],stage1_4[172],stage1_3[186]}
   );
   gpc615_5 gpc187 (
      {stage0_3[401], stage0_3[402], stage0_3[403], stage0_3[404], stage0_3[405]},
      {stage0_4[188]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[43],stage1_5[89],stage1_4[173],stage1_3[187]}
   );
   gpc615_5 gpc188 (
      {stage0_3[406], stage0_3[407], stage0_3[408], stage0_3[409], stage0_3[410]},
      {stage0_4[189]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[44],stage1_5[90],stage1_4[174],stage1_3[188]}
   );
   gpc615_5 gpc189 (
      {stage0_3[411], stage0_3[412], stage0_3[413], stage0_3[414], stage0_3[415]},
      {stage0_4[190]},
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage1_7[16],stage1_6[45],stage1_5[91],stage1_4[175],stage1_3[189]}
   );
   gpc615_5 gpc190 (
      {stage0_3[416], stage0_3[417], stage0_3[418], stage0_3[419], stage0_3[420]},
      {stage0_4[191]},
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage1_7[17],stage1_6[46],stage1_5[92],stage1_4[176],stage1_3[190]}
   );
   gpc615_5 gpc191 (
      {stage0_3[421], stage0_3[422], stage0_3[423], stage0_3[424], stage0_3[425]},
      {stage0_4[192]},
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage1_7[18],stage1_6[47],stage1_5[93],stage1_4[177],stage1_3[191]}
   );
   gpc615_5 gpc192 (
      {stage0_3[426], stage0_3[427], stage0_3[428], stage0_3[429], stage0_3[430]},
      {stage0_4[193]},
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage1_7[19],stage1_6[48],stage1_5[94],stage1_4[178],stage1_3[192]}
   );
   gpc615_5 gpc193 (
      {stage0_3[431], stage0_3[432], stage0_3[433], stage0_3[434], stage0_3[435]},
      {stage0_4[194]},
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage1_7[20],stage1_6[49],stage1_5[95],stage1_4[179],stage1_3[193]}
   );
   gpc615_5 gpc194 (
      {stage0_3[436], stage0_3[437], stage0_3[438], stage0_3[439], stage0_3[440]},
      {stage0_4[195]},
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage1_7[21],stage1_6[50],stage1_5[96],stage1_4[180],stage1_3[194]}
   );
   gpc615_5 gpc195 (
      {stage0_3[441], stage0_3[442], stage0_3[443], stage0_3[444], stage0_3[445]},
      {stage0_4[196]},
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage1_7[22],stage1_6[51],stage1_5[97],stage1_4[181],stage1_3[195]}
   );
   gpc615_5 gpc196 (
      {stage0_3[446], stage0_3[447], stage0_3[448], stage0_3[449], stage0_3[450]},
      {stage0_4[197]},
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage1_7[23],stage1_6[52],stage1_5[98],stage1_4[182],stage1_3[196]}
   );
   gpc615_5 gpc197 (
      {stage0_3[451], stage0_3[452], stage0_3[453], stage0_3[454], stage0_3[455]},
      {stage0_4[198]},
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage1_7[24],stage1_6[53],stage1_5[99],stage1_4[183],stage1_3[197]}
   );
   gpc615_5 gpc198 (
      {stage0_3[456], stage0_3[457], stage0_3[458], stage0_3[459], stage0_3[460]},
      {stage0_4[199]},
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage1_7[25],stage1_6[54],stage1_5[100],stage1_4[184],stage1_3[198]}
   );
   gpc615_5 gpc199 (
      {stage0_3[461], stage0_3[462], stage0_3[463], stage0_3[464], stage0_3[465]},
      {stage0_4[200]},
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage1_7[26],stage1_6[55],stage1_5[101],stage1_4[185],stage1_3[199]}
   );
   gpc606_5 gpc200 (
      {stage0_4[201], stage0_4[202], stage0_4[203], stage0_4[204], stage0_4[205], stage0_4[206]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[27],stage1_6[56],stage1_5[102],stage1_4[186]}
   );
   gpc606_5 gpc201 (
      {stage0_4[207], stage0_4[208], stage0_4[209], stage0_4[210], stage0_4[211], stage0_4[212]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[28],stage1_6[57],stage1_5[103],stage1_4[187]}
   );
   gpc606_5 gpc202 (
      {stage0_4[213], stage0_4[214], stage0_4[215], stage0_4[216], stage0_4[217], stage0_4[218]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[29],stage1_6[58],stage1_5[104],stage1_4[188]}
   );
   gpc606_5 gpc203 (
      {stage0_4[219], stage0_4[220], stage0_4[221], stage0_4[222], stage0_4[223], stage0_4[224]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[30],stage1_6[59],stage1_5[105],stage1_4[189]}
   );
   gpc606_5 gpc204 (
      {stage0_4[225], stage0_4[226], stage0_4[227], stage0_4[228], stage0_4[229], stage0_4[230]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[31],stage1_6[60],stage1_5[106],stage1_4[190]}
   );
   gpc606_5 gpc205 (
      {stage0_4[231], stage0_4[232], stage0_4[233], stage0_4[234], stage0_4[235], stage0_4[236]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[32],stage1_6[61],stage1_5[107],stage1_4[191]}
   );
   gpc606_5 gpc206 (
      {stage0_4[237], stage0_4[238], stage0_4[239], stage0_4[240], stage0_4[241], stage0_4[242]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[33],stage1_6[62],stage1_5[108],stage1_4[192]}
   );
   gpc606_5 gpc207 (
      {stage0_4[243], stage0_4[244], stage0_4[245], stage0_4[246], stage0_4[247], stage0_4[248]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[34],stage1_6[63],stage1_5[109],stage1_4[193]}
   );
   gpc606_5 gpc208 (
      {stage0_4[249], stage0_4[250], stage0_4[251], stage0_4[252], stage0_4[253], stage0_4[254]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[35],stage1_6[64],stage1_5[110],stage1_4[194]}
   );
   gpc606_5 gpc209 (
      {stage0_4[255], stage0_4[256], stage0_4[257], stage0_4[258], stage0_4[259], stage0_4[260]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[36],stage1_6[65],stage1_5[111],stage1_4[195]}
   );
   gpc606_5 gpc210 (
      {stage0_4[261], stage0_4[262], stage0_4[263], stage0_4[264], stage0_4[265], stage0_4[266]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[37],stage1_6[66],stage1_5[112],stage1_4[196]}
   );
   gpc606_5 gpc211 (
      {stage0_4[267], stage0_4[268], stage0_4[269], stage0_4[270], stage0_4[271], stage0_4[272]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[38],stage1_6[67],stage1_5[113],stage1_4[197]}
   );
   gpc606_5 gpc212 (
      {stage0_4[273], stage0_4[274], stage0_4[275], stage0_4[276], stage0_4[277], stage0_4[278]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[39],stage1_6[68],stage1_5[114],stage1_4[198]}
   );
   gpc606_5 gpc213 (
      {stage0_4[279], stage0_4[280], stage0_4[281], stage0_4[282], stage0_4[283], stage0_4[284]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[40],stage1_6[69],stage1_5[115],stage1_4[199]}
   );
   gpc606_5 gpc214 (
      {stage0_4[285], stage0_4[286], stage0_4[287], stage0_4[288], stage0_4[289], stage0_4[290]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[41],stage1_6[70],stage1_5[116],stage1_4[200]}
   );
   gpc606_5 gpc215 (
      {stage0_4[291], stage0_4[292], stage0_4[293], stage0_4[294], stage0_4[295], stage0_4[296]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[42],stage1_6[71],stage1_5[117],stage1_4[201]}
   );
   gpc606_5 gpc216 (
      {stage0_4[297], stage0_4[298], stage0_4[299], stage0_4[300], stage0_4[301], stage0_4[302]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[43],stage1_6[72],stage1_5[118],stage1_4[202]}
   );
   gpc606_5 gpc217 (
      {stage0_4[303], stage0_4[304], stage0_4[305], stage0_4[306], stage0_4[307], stage0_4[308]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[44],stage1_6[73],stage1_5[119],stage1_4[203]}
   );
   gpc606_5 gpc218 (
      {stage0_4[309], stage0_4[310], stage0_4[311], stage0_4[312], stage0_4[313], stage0_4[314]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[45],stage1_6[74],stage1_5[120],stage1_4[204]}
   );
   gpc606_5 gpc219 (
      {stage0_4[315], stage0_4[316], stage0_4[317], stage0_4[318], stage0_4[319], stage0_4[320]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[46],stage1_6[75],stage1_5[121],stage1_4[205]}
   );
   gpc606_5 gpc220 (
      {stage0_4[321], stage0_4[322], stage0_4[323], stage0_4[324], stage0_4[325], stage0_4[326]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[47],stage1_6[76],stage1_5[122],stage1_4[206]}
   );
   gpc606_5 gpc221 (
      {stage0_4[327], stage0_4[328], stage0_4[329], stage0_4[330], stage0_4[331], stage0_4[332]},
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage1_8[21],stage1_7[48],stage1_6[77],stage1_5[123],stage1_4[207]}
   );
   gpc606_5 gpc222 (
      {stage0_4[333], stage0_4[334], stage0_4[335], stage0_4[336], stage0_4[337], stage0_4[338]},
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage1_8[22],stage1_7[49],stage1_6[78],stage1_5[124],stage1_4[208]}
   );
   gpc606_5 gpc223 (
      {stage0_4[339], stage0_4[340], stage0_4[341], stage0_4[342], stage0_4[343], stage0_4[344]},
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage1_8[23],stage1_7[50],stage1_6[79],stage1_5[125],stage1_4[209]}
   );
   gpc606_5 gpc224 (
      {stage0_4[345], stage0_4[346], stage0_4[347], stage0_4[348], stage0_4[349], stage0_4[350]},
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage1_8[24],stage1_7[51],stage1_6[80],stage1_5[126],stage1_4[210]}
   );
   gpc606_5 gpc225 (
      {stage0_4[351], stage0_4[352], stage0_4[353], stage0_4[354], stage0_4[355], stage0_4[356]},
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage1_8[25],stage1_7[52],stage1_6[81],stage1_5[127],stage1_4[211]}
   );
   gpc606_5 gpc226 (
      {stage0_4[357], stage0_4[358], stage0_4[359], stage0_4[360], stage0_4[361], stage0_4[362]},
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage1_8[26],stage1_7[53],stage1_6[82],stage1_5[128],stage1_4[212]}
   );
   gpc606_5 gpc227 (
      {stage0_4[363], stage0_4[364], stage0_4[365], stage0_4[366], stage0_4[367], stage0_4[368]},
      {stage0_6[162], stage0_6[163], stage0_6[164], stage0_6[165], stage0_6[166], stage0_6[167]},
      {stage1_8[27],stage1_7[54],stage1_6[83],stage1_5[129],stage1_4[213]}
   );
   gpc606_5 gpc228 (
      {stage0_4[369], stage0_4[370], stage0_4[371], stage0_4[372], stage0_4[373], stage0_4[374]},
      {stage0_6[168], stage0_6[169], stage0_6[170], stage0_6[171], stage0_6[172], stage0_6[173]},
      {stage1_8[28],stage1_7[55],stage1_6[84],stage1_5[130],stage1_4[214]}
   );
   gpc606_5 gpc229 (
      {stage0_4[375], stage0_4[376], stage0_4[377], stage0_4[378], stage0_4[379], stage0_4[380]},
      {stage0_6[174], stage0_6[175], stage0_6[176], stage0_6[177], stage0_6[178], stage0_6[179]},
      {stage1_8[29],stage1_7[56],stage1_6[85],stage1_5[131],stage1_4[215]}
   );
   gpc606_5 gpc230 (
      {stage0_4[381], stage0_4[382], stage0_4[383], stage0_4[384], stage0_4[385], stage0_4[386]},
      {stage0_6[180], stage0_6[181], stage0_6[182], stage0_6[183], stage0_6[184], stage0_6[185]},
      {stage1_8[30],stage1_7[57],stage1_6[86],stage1_5[132],stage1_4[216]}
   );
   gpc606_5 gpc231 (
      {stage0_4[387], stage0_4[388], stage0_4[389], stage0_4[390], stage0_4[391], stage0_4[392]},
      {stage0_6[186], stage0_6[187], stage0_6[188], stage0_6[189], stage0_6[190], stage0_6[191]},
      {stage1_8[31],stage1_7[58],stage1_6[87],stage1_5[133],stage1_4[217]}
   );
   gpc606_5 gpc232 (
      {stage0_4[393], stage0_4[394], stage0_4[395], stage0_4[396], stage0_4[397], stage0_4[398]},
      {stage0_6[192], stage0_6[193], stage0_6[194], stage0_6[195], stage0_6[196], stage0_6[197]},
      {stage1_8[32],stage1_7[59],stage1_6[88],stage1_5[134],stage1_4[218]}
   );
   gpc606_5 gpc233 (
      {stage0_4[399], stage0_4[400], stage0_4[401], stage0_4[402], stage0_4[403], stage0_4[404]},
      {stage0_6[198], stage0_6[199], stage0_6[200], stage0_6[201], stage0_6[202], stage0_6[203]},
      {stage1_8[33],stage1_7[60],stage1_6[89],stage1_5[135],stage1_4[219]}
   );
   gpc606_5 gpc234 (
      {stage0_4[405], stage0_4[406], stage0_4[407], stage0_4[408], stage0_4[409], stage0_4[410]},
      {stage0_6[204], stage0_6[205], stage0_6[206], stage0_6[207], stage0_6[208], stage0_6[209]},
      {stage1_8[34],stage1_7[61],stage1_6[90],stage1_5[136],stage1_4[220]}
   );
   gpc606_5 gpc235 (
      {stage0_4[411], stage0_4[412], stage0_4[413], stage0_4[414], stage0_4[415], stage0_4[416]},
      {stage0_6[210], stage0_6[211], stage0_6[212], stage0_6[213], stage0_6[214], stage0_6[215]},
      {stage1_8[35],stage1_7[62],stage1_6[91],stage1_5[137],stage1_4[221]}
   );
   gpc615_5 gpc236 (
      {stage0_4[417], stage0_4[418], stage0_4[419], stage0_4[420], stage0_4[421]},
      {stage0_5[162]},
      {stage0_6[216], stage0_6[217], stage0_6[218], stage0_6[219], stage0_6[220], stage0_6[221]},
      {stage1_8[36],stage1_7[63],stage1_6[92],stage1_5[138],stage1_4[222]}
   );
   gpc615_5 gpc237 (
      {stage0_4[422], stage0_4[423], stage0_4[424], stage0_4[425], stage0_4[426]},
      {stage0_5[163]},
      {stage0_6[222], stage0_6[223], stage0_6[224], stage0_6[225], stage0_6[226], stage0_6[227]},
      {stage1_8[37],stage1_7[64],stage1_6[93],stage1_5[139],stage1_4[223]}
   );
   gpc615_5 gpc238 (
      {stage0_4[427], stage0_4[428], stage0_4[429], stage0_4[430], stage0_4[431]},
      {stage0_5[164]},
      {stage0_6[228], stage0_6[229], stage0_6[230], stage0_6[231], stage0_6[232], stage0_6[233]},
      {stage1_8[38],stage1_7[65],stage1_6[94],stage1_5[140],stage1_4[224]}
   );
   gpc615_5 gpc239 (
      {stage0_4[432], stage0_4[433], stage0_4[434], stage0_4[435], stage0_4[436]},
      {stage0_5[165]},
      {stage0_6[234], stage0_6[235], stage0_6[236], stage0_6[237], stage0_6[238], stage0_6[239]},
      {stage1_8[39],stage1_7[66],stage1_6[95],stage1_5[141],stage1_4[225]}
   );
   gpc615_5 gpc240 (
      {stage0_4[437], stage0_4[438], stage0_4[439], stage0_4[440], stage0_4[441]},
      {stage0_5[166]},
      {stage0_6[240], stage0_6[241], stage0_6[242], stage0_6[243], stage0_6[244], stage0_6[245]},
      {stage1_8[40],stage1_7[67],stage1_6[96],stage1_5[142],stage1_4[226]}
   );
   gpc615_5 gpc241 (
      {stage0_4[442], stage0_4[443], stage0_4[444], stage0_4[445], stage0_4[446]},
      {stage0_5[167]},
      {stage0_6[246], stage0_6[247], stage0_6[248], stage0_6[249], stage0_6[250], stage0_6[251]},
      {stage1_8[41],stage1_7[68],stage1_6[97],stage1_5[143],stage1_4[227]}
   );
   gpc615_5 gpc242 (
      {stage0_4[447], stage0_4[448], stage0_4[449], stage0_4[450], stage0_4[451]},
      {stage0_5[168]},
      {stage0_6[252], stage0_6[253], stage0_6[254], stage0_6[255], stage0_6[256], stage0_6[257]},
      {stage1_8[42],stage1_7[69],stage1_6[98],stage1_5[144],stage1_4[228]}
   );
   gpc615_5 gpc243 (
      {stage0_4[452], stage0_4[453], stage0_4[454], stage0_4[455], stage0_4[456]},
      {stage0_5[169]},
      {stage0_6[258], stage0_6[259], stage0_6[260], stage0_6[261], stage0_6[262], stage0_6[263]},
      {stage1_8[43],stage1_7[70],stage1_6[99],stage1_5[145],stage1_4[229]}
   );
   gpc615_5 gpc244 (
      {stage0_4[457], stage0_4[458], stage0_4[459], stage0_4[460], stage0_4[461]},
      {stage0_5[170]},
      {stage0_6[264], stage0_6[265], stage0_6[266], stage0_6[267], stage0_6[268], stage0_6[269]},
      {stage1_8[44],stage1_7[71],stage1_6[100],stage1_5[146],stage1_4[230]}
   );
   gpc615_5 gpc245 (
      {stage0_4[462], stage0_4[463], stage0_4[464], stage0_4[465], stage0_4[466]},
      {stage0_5[171]},
      {stage0_6[270], stage0_6[271], stage0_6[272], stage0_6[273], stage0_6[274], stage0_6[275]},
      {stage1_8[45],stage1_7[72],stage1_6[101],stage1_5[147],stage1_4[231]}
   );
   gpc615_5 gpc246 (
      {stage0_4[467], stage0_4[468], stage0_4[469], stage0_4[470], stage0_4[471]},
      {stage0_5[172]},
      {stage0_6[276], stage0_6[277], stage0_6[278], stage0_6[279], stage0_6[280], stage0_6[281]},
      {stage1_8[46],stage1_7[73],stage1_6[102],stage1_5[148],stage1_4[232]}
   );
   gpc615_5 gpc247 (
      {stage0_4[472], stage0_4[473], stage0_4[474], stage0_4[475], stage0_4[476]},
      {stage0_5[173]},
      {stage0_6[282], stage0_6[283], stage0_6[284], stage0_6[285], stage0_6[286], stage0_6[287]},
      {stage1_8[47],stage1_7[74],stage1_6[103],stage1_5[149],stage1_4[233]}
   );
   gpc615_5 gpc248 (
      {stage0_4[477], stage0_4[478], stage0_4[479], stage0_4[480], stage0_4[481]},
      {stage0_5[174]},
      {stage0_6[288], stage0_6[289], stage0_6[290], stage0_6[291], stage0_6[292], stage0_6[293]},
      {stage1_8[48],stage1_7[75],stage1_6[104],stage1_5[150],stage1_4[234]}
   );
   gpc615_5 gpc249 (
      {stage0_4[482], stage0_4[483], stage0_4[484], stage0_4[485], stage0_4[486]},
      {stage0_5[175]},
      {stage0_6[294], stage0_6[295], stage0_6[296], stage0_6[297], stage0_6[298], stage0_6[299]},
      {stage1_8[49],stage1_7[76],stage1_6[105],stage1_5[151],stage1_4[235]}
   );
   gpc615_5 gpc250 (
      {stage0_4[487], stage0_4[488], stage0_4[489], stage0_4[490], stage0_4[491]},
      {stage0_5[176]},
      {stage0_6[300], stage0_6[301], stage0_6[302], stage0_6[303], stage0_6[304], stage0_6[305]},
      {stage1_8[50],stage1_7[77],stage1_6[106],stage1_5[152],stage1_4[236]}
   );
   gpc615_5 gpc251 (
      {stage0_4[492], stage0_4[493], stage0_4[494], stage0_4[495], stage0_4[496]},
      {stage0_5[177]},
      {stage0_6[306], stage0_6[307], stage0_6[308], stage0_6[309], stage0_6[310], stage0_6[311]},
      {stage1_8[51],stage1_7[78],stage1_6[107],stage1_5[153],stage1_4[237]}
   );
   gpc615_5 gpc252 (
      {stage0_4[497], stage0_4[498], stage0_4[499], stage0_4[500], stage0_4[501]},
      {stage0_5[178]},
      {stage0_6[312], stage0_6[313], stage0_6[314], stage0_6[315], stage0_6[316], stage0_6[317]},
      {stage1_8[52],stage1_7[79],stage1_6[108],stage1_5[154],stage1_4[238]}
   );
   gpc615_5 gpc253 (
      {stage0_4[502], stage0_4[503], stage0_4[504], stage0_4[505], stage0_4[506]},
      {stage0_5[179]},
      {stage0_6[318], stage0_6[319], stage0_6[320], stage0_6[321], stage0_6[322], stage0_6[323]},
      {stage1_8[53],stage1_7[80],stage1_6[109],stage1_5[155],stage1_4[239]}
   );
   gpc615_5 gpc254 (
      {stage0_4[507], stage0_4[508], stage0_4[509], stage0_4[510], stage0_4[511]},
      {stage0_5[180]},
      {stage0_6[324], stage0_6[325], stage0_6[326], stage0_6[327], stage0_6[328], stage0_6[329]},
      {stage1_8[54],stage1_7[81],stage1_6[110],stage1_5[156],stage1_4[240]}
   );
   gpc606_5 gpc255 (
      {stage0_5[181], stage0_5[182], stage0_5[183], stage0_5[184], stage0_5[185], stage0_5[186]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[55],stage1_7[82],stage1_6[111],stage1_5[157]}
   );
   gpc606_5 gpc256 (
      {stage0_5[187], stage0_5[188], stage0_5[189], stage0_5[190], stage0_5[191], stage0_5[192]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[56],stage1_7[83],stage1_6[112],stage1_5[158]}
   );
   gpc606_5 gpc257 (
      {stage0_5[193], stage0_5[194], stage0_5[195], stage0_5[196], stage0_5[197], stage0_5[198]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[57],stage1_7[84],stage1_6[113],stage1_5[159]}
   );
   gpc606_5 gpc258 (
      {stage0_5[199], stage0_5[200], stage0_5[201], stage0_5[202], stage0_5[203], stage0_5[204]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[58],stage1_7[85],stage1_6[114],stage1_5[160]}
   );
   gpc606_5 gpc259 (
      {stage0_5[205], stage0_5[206], stage0_5[207], stage0_5[208], stage0_5[209], stage0_5[210]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[59],stage1_7[86],stage1_6[115],stage1_5[161]}
   );
   gpc606_5 gpc260 (
      {stage0_5[211], stage0_5[212], stage0_5[213], stage0_5[214], stage0_5[215], stage0_5[216]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[60],stage1_7[87],stage1_6[116],stage1_5[162]}
   );
   gpc606_5 gpc261 (
      {stage0_5[217], stage0_5[218], stage0_5[219], stage0_5[220], stage0_5[221], stage0_5[222]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[61],stage1_7[88],stage1_6[117],stage1_5[163]}
   );
   gpc606_5 gpc262 (
      {stage0_5[223], stage0_5[224], stage0_5[225], stage0_5[226], stage0_5[227], stage0_5[228]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[62],stage1_7[89],stage1_6[118],stage1_5[164]}
   );
   gpc606_5 gpc263 (
      {stage0_5[229], stage0_5[230], stage0_5[231], stage0_5[232], stage0_5[233], stage0_5[234]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[63],stage1_7[90],stage1_6[119],stage1_5[165]}
   );
   gpc606_5 gpc264 (
      {stage0_5[235], stage0_5[236], stage0_5[237], stage0_5[238], stage0_5[239], stage0_5[240]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[64],stage1_7[91],stage1_6[120],stage1_5[166]}
   );
   gpc606_5 gpc265 (
      {stage0_5[241], stage0_5[242], stage0_5[243], stage0_5[244], stage0_5[245], stage0_5[246]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[65],stage1_7[92],stage1_6[121],stage1_5[167]}
   );
   gpc606_5 gpc266 (
      {stage0_5[247], stage0_5[248], stage0_5[249], stage0_5[250], stage0_5[251], stage0_5[252]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[66],stage1_7[93],stage1_6[122],stage1_5[168]}
   );
   gpc606_5 gpc267 (
      {stage0_5[253], stage0_5[254], stage0_5[255], stage0_5[256], stage0_5[257], stage0_5[258]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[67],stage1_7[94],stage1_6[123],stage1_5[169]}
   );
   gpc606_5 gpc268 (
      {stage0_5[259], stage0_5[260], stage0_5[261], stage0_5[262], stage0_5[263], stage0_5[264]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[68],stage1_7[95],stage1_6[124],stage1_5[170]}
   );
   gpc606_5 gpc269 (
      {stage0_5[265], stage0_5[266], stage0_5[267], stage0_5[268], stage0_5[269], stage0_5[270]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[69],stage1_7[96],stage1_6[125],stage1_5[171]}
   );
   gpc606_5 gpc270 (
      {stage0_5[271], stage0_5[272], stage0_5[273], stage0_5[274], stage0_5[275], stage0_5[276]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[70],stage1_7[97],stage1_6[126],stage1_5[172]}
   );
   gpc606_5 gpc271 (
      {stage0_5[277], stage0_5[278], stage0_5[279], stage0_5[280], stage0_5[281], stage0_5[282]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[71],stage1_7[98],stage1_6[127],stage1_5[173]}
   );
   gpc606_5 gpc272 (
      {stage0_5[283], stage0_5[284], stage0_5[285], stage0_5[286], stage0_5[287], stage0_5[288]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[72],stage1_7[99],stage1_6[128],stage1_5[174]}
   );
   gpc606_5 gpc273 (
      {stage0_5[289], stage0_5[290], stage0_5[291], stage0_5[292], stage0_5[293], stage0_5[294]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[73],stage1_7[100],stage1_6[129],stage1_5[175]}
   );
   gpc606_5 gpc274 (
      {stage0_5[295], stage0_5[296], stage0_5[297], stage0_5[298], stage0_5[299], stage0_5[300]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[74],stage1_7[101],stage1_6[130],stage1_5[176]}
   );
   gpc606_5 gpc275 (
      {stage0_5[301], stage0_5[302], stage0_5[303], stage0_5[304], stage0_5[305], stage0_5[306]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[75],stage1_7[102],stage1_6[131],stage1_5[177]}
   );
   gpc606_5 gpc276 (
      {stage0_5[307], stage0_5[308], stage0_5[309], stage0_5[310], stage0_5[311], stage0_5[312]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[76],stage1_7[103],stage1_6[132],stage1_5[178]}
   );
   gpc606_5 gpc277 (
      {stage0_5[313], stage0_5[314], stage0_5[315], stage0_5[316], stage0_5[317], stage0_5[318]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[77],stage1_7[104],stage1_6[133],stage1_5[179]}
   );
   gpc606_5 gpc278 (
      {stage0_5[319], stage0_5[320], stage0_5[321], stage0_5[322], stage0_5[323], stage0_5[324]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[78],stage1_7[105],stage1_6[134],stage1_5[180]}
   );
   gpc606_5 gpc279 (
      {stage0_5[325], stage0_5[326], stage0_5[327], stage0_5[328], stage0_5[329], stage0_5[330]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[79],stage1_7[106],stage1_6[135],stage1_5[181]}
   );
   gpc606_5 gpc280 (
      {stage0_5[331], stage0_5[332], stage0_5[333], stage0_5[334], stage0_5[335], stage0_5[336]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[80],stage1_7[107],stage1_6[136],stage1_5[182]}
   );
   gpc606_5 gpc281 (
      {stage0_5[337], stage0_5[338], stage0_5[339], stage0_5[340], stage0_5[341], stage0_5[342]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[81],stage1_7[108],stage1_6[137],stage1_5[183]}
   );
   gpc606_5 gpc282 (
      {stage0_5[343], stage0_5[344], stage0_5[345], stage0_5[346], stage0_5[347], stage0_5[348]},
      {stage0_7[162], stage0_7[163], stage0_7[164], stage0_7[165], stage0_7[166], stage0_7[167]},
      {stage1_9[27],stage1_8[82],stage1_7[109],stage1_6[138],stage1_5[184]}
   );
   gpc606_5 gpc283 (
      {stage0_5[349], stage0_5[350], stage0_5[351], stage0_5[352], stage0_5[353], stage0_5[354]},
      {stage0_7[168], stage0_7[169], stage0_7[170], stage0_7[171], stage0_7[172], stage0_7[173]},
      {stage1_9[28],stage1_8[83],stage1_7[110],stage1_6[139],stage1_5[185]}
   );
   gpc606_5 gpc284 (
      {stage0_5[355], stage0_5[356], stage0_5[357], stage0_5[358], stage0_5[359], stage0_5[360]},
      {stage0_7[174], stage0_7[175], stage0_7[176], stage0_7[177], stage0_7[178], stage0_7[179]},
      {stage1_9[29],stage1_8[84],stage1_7[111],stage1_6[140],stage1_5[186]}
   );
   gpc606_5 gpc285 (
      {stage0_5[361], stage0_5[362], stage0_5[363], stage0_5[364], stage0_5[365], stage0_5[366]},
      {stage0_7[180], stage0_7[181], stage0_7[182], stage0_7[183], stage0_7[184], stage0_7[185]},
      {stage1_9[30],stage1_8[85],stage1_7[112],stage1_6[141],stage1_5[187]}
   );
   gpc606_5 gpc286 (
      {stage0_5[367], stage0_5[368], stage0_5[369], stage0_5[370], stage0_5[371], stage0_5[372]},
      {stage0_7[186], stage0_7[187], stage0_7[188], stage0_7[189], stage0_7[190], stage0_7[191]},
      {stage1_9[31],stage1_8[86],stage1_7[113],stage1_6[142],stage1_5[188]}
   );
   gpc606_5 gpc287 (
      {stage0_5[373], stage0_5[374], stage0_5[375], stage0_5[376], stage0_5[377], stage0_5[378]},
      {stage0_7[192], stage0_7[193], stage0_7[194], stage0_7[195], stage0_7[196], stage0_7[197]},
      {stage1_9[32],stage1_8[87],stage1_7[114],stage1_6[143],stage1_5[189]}
   );
   gpc606_5 gpc288 (
      {stage0_5[379], stage0_5[380], stage0_5[381], stage0_5[382], stage0_5[383], stage0_5[384]},
      {stage0_7[198], stage0_7[199], stage0_7[200], stage0_7[201], stage0_7[202], stage0_7[203]},
      {stage1_9[33],stage1_8[88],stage1_7[115],stage1_6[144],stage1_5[190]}
   );
   gpc606_5 gpc289 (
      {stage0_5[385], stage0_5[386], stage0_5[387], stage0_5[388], stage0_5[389], stage0_5[390]},
      {stage0_7[204], stage0_7[205], stage0_7[206], stage0_7[207], stage0_7[208], stage0_7[209]},
      {stage1_9[34],stage1_8[89],stage1_7[116],stage1_6[145],stage1_5[191]}
   );
   gpc606_5 gpc290 (
      {stage0_5[391], stage0_5[392], stage0_5[393], stage0_5[394], stage0_5[395], stage0_5[396]},
      {stage0_7[210], stage0_7[211], stage0_7[212], stage0_7[213], stage0_7[214], stage0_7[215]},
      {stage1_9[35],stage1_8[90],stage1_7[117],stage1_6[146],stage1_5[192]}
   );
   gpc606_5 gpc291 (
      {stage0_5[397], stage0_5[398], stage0_5[399], stage0_5[400], stage0_5[401], stage0_5[402]},
      {stage0_7[216], stage0_7[217], stage0_7[218], stage0_7[219], stage0_7[220], stage0_7[221]},
      {stage1_9[36],stage1_8[91],stage1_7[118],stage1_6[147],stage1_5[193]}
   );
   gpc606_5 gpc292 (
      {stage0_5[403], stage0_5[404], stage0_5[405], stage0_5[406], stage0_5[407], stage0_5[408]},
      {stage0_7[222], stage0_7[223], stage0_7[224], stage0_7[225], stage0_7[226], stage0_7[227]},
      {stage1_9[37],stage1_8[92],stage1_7[119],stage1_6[148],stage1_5[194]}
   );
   gpc606_5 gpc293 (
      {stage0_5[409], stage0_5[410], stage0_5[411], stage0_5[412], stage0_5[413], stage0_5[414]},
      {stage0_7[228], stage0_7[229], stage0_7[230], stage0_7[231], stage0_7[232], stage0_7[233]},
      {stage1_9[38],stage1_8[93],stage1_7[120],stage1_6[149],stage1_5[195]}
   );
   gpc606_5 gpc294 (
      {stage0_5[415], stage0_5[416], stage0_5[417], stage0_5[418], stage0_5[419], stage0_5[420]},
      {stage0_7[234], stage0_7[235], stage0_7[236], stage0_7[237], stage0_7[238], stage0_7[239]},
      {stage1_9[39],stage1_8[94],stage1_7[121],stage1_6[150],stage1_5[196]}
   );
   gpc606_5 gpc295 (
      {stage0_5[421], stage0_5[422], stage0_5[423], stage0_5[424], stage0_5[425], stage0_5[426]},
      {stage0_7[240], stage0_7[241], stage0_7[242], stage0_7[243], stage0_7[244], stage0_7[245]},
      {stage1_9[40],stage1_8[95],stage1_7[122],stage1_6[151],stage1_5[197]}
   );
   gpc606_5 gpc296 (
      {stage0_5[427], stage0_5[428], stage0_5[429], stage0_5[430], stage0_5[431], stage0_5[432]},
      {stage0_7[246], stage0_7[247], stage0_7[248], stage0_7[249], stage0_7[250], stage0_7[251]},
      {stage1_9[41],stage1_8[96],stage1_7[123],stage1_6[152],stage1_5[198]}
   );
   gpc606_5 gpc297 (
      {stage0_5[433], stage0_5[434], stage0_5[435], stage0_5[436], stage0_5[437], stage0_5[438]},
      {stage0_7[252], stage0_7[253], stage0_7[254], stage0_7[255], stage0_7[256], stage0_7[257]},
      {stage1_9[42],stage1_8[97],stage1_7[124],stage1_6[153],stage1_5[199]}
   );
   gpc606_5 gpc298 (
      {stage0_5[439], stage0_5[440], stage0_5[441], stage0_5[442], stage0_5[443], stage0_5[444]},
      {stage0_7[258], stage0_7[259], stage0_7[260], stage0_7[261], stage0_7[262], stage0_7[263]},
      {stage1_9[43],stage1_8[98],stage1_7[125],stage1_6[154],stage1_5[200]}
   );
   gpc606_5 gpc299 (
      {stage0_5[445], stage0_5[446], stage0_5[447], stage0_5[448], stage0_5[449], stage0_5[450]},
      {stage0_7[264], stage0_7[265], stage0_7[266], stage0_7[267], stage0_7[268], stage0_7[269]},
      {stage1_9[44],stage1_8[99],stage1_7[126],stage1_6[155],stage1_5[201]}
   );
   gpc606_5 gpc300 (
      {stage0_5[451], stage0_5[452], stage0_5[453], stage0_5[454], stage0_5[455], stage0_5[456]},
      {stage0_7[270], stage0_7[271], stage0_7[272], stage0_7[273], stage0_7[274], stage0_7[275]},
      {stage1_9[45],stage1_8[100],stage1_7[127],stage1_6[156],stage1_5[202]}
   );
   gpc606_5 gpc301 (
      {stage0_5[457], stage0_5[458], stage0_5[459], stage0_5[460], stage0_5[461], stage0_5[462]},
      {stage0_7[276], stage0_7[277], stage0_7[278], stage0_7[279], stage0_7[280], stage0_7[281]},
      {stage1_9[46],stage1_8[101],stage1_7[128],stage1_6[157],stage1_5[203]}
   );
   gpc606_5 gpc302 (
      {stage0_5[463], stage0_5[464], stage0_5[465], stage0_5[466], stage0_5[467], stage0_5[468]},
      {stage0_7[282], stage0_7[283], stage0_7[284], stage0_7[285], stage0_7[286], stage0_7[287]},
      {stage1_9[47],stage1_8[102],stage1_7[129],stage1_6[158],stage1_5[204]}
   );
   gpc606_5 gpc303 (
      {stage0_5[469], stage0_5[470], stage0_5[471], stage0_5[472], stage0_5[473], stage0_5[474]},
      {stage0_7[288], stage0_7[289], stage0_7[290], stage0_7[291], stage0_7[292], stage0_7[293]},
      {stage1_9[48],stage1_8[103],stage1_7[130],stage1_6[159],stage1_5[205]}
   );
   gpc606_5 gpc304 (
      {stage0_5[475], stage0_5[476], stage0_5[477], stage0_5[478], stage0_5[479], stage0_5[480]},
      {stage0_7[294], stage0_7[295], stage0_7[296], stage0_7[297], stage0_7[298], stage0_7[299]},
      {stage1_9[49],stage1_8[104],stage1_7[131],stage1_6[160],stage1_5[206]}
   );
   gpc606_5 gpc305 (
      {stage0_5[481], stage0_5[482], stage0_5[483], stage0_5[484], stage0_5[485], stage0_5[486]},
      {stage0_7[300], stage0_7[301], stage0_7[302], stage0_7[303], stage0_7[304], stage0_7[305]},
      {stage1_9[50],stage1_8[105],stage1_7[132],stage1_6[161],stage1_5[207]}
   );
   gpc606_5 gpc306 (
      {stage0_5[487], stage0_5[488], stage0_5[489], stage0_5[490], stage0_5[491], stage0_5[492]},
      {stage0_7[306], stage0_7[307], stage0_7[308], stage0_7[309], stage0_7[310], stage0_7[311]},
      {stage1_9[51],stage1_8[106],stage1_7[133],stage1_6[162],stage1_5[208]}
   );
   gpc606_5 gpc307 (
      {stage0_5[493], stage0_5[494], stage0_5[495], stage0_5[496], stage0_5[497], stage0_5[498]},
      {stage0_7[312], stage0_7[313], stage0_7[314], stage0_7[315], stage0_7[316], stage0_7[317]},
      {stage1_9[52],stage1_8[107],stage1_7[134],stage1_6[163],stage1_5[209]}
   );
   gpc606_5 gpc308 (
      {stage0_5[499], stage0_5[500], stage0_5[501], stage0_5[502], stage0_5[503], stage0_5[504]},
      {stage0_7[318], stage0_7[319], stage0_7[320], stage0_7[321], stage0_7[322], stage0_7[323]},
      {stage1_9[53],stage1_8[108],stage1_7[135],stage1_6[164],stage1_5[210]}
   );
   gpc615_5 gpc309 (
      {stage0_6[330], stage0_6[331], stage0_6[332], stage0_6[333], stage0_6[334]},
      {stage0_7[324]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[54],stage1_8[109],stage1_7[136],stage1_6[165]}
   );
   gpc615_5 gpc310 (
      {stage0_6[335], stage0_6[336], stage0_6[337], stage0_6[338], stage0_6[339]},
      {stage0_7[325]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[55],stage1_8[110],stage1_7[137],stage1_6[166]}
   );
   gpc615_5 gpc311 (
      {stage0_6[340], stage0_6[341], stage0_6[342], stage0_6[343], stage0_6[344]},
      {stage0_7[326]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[56],stage1_8[111],stage1_7[138],stage1_6[167]}
   );
   gpc615_5 gpc312 (
      {stage0_6[345], stage0_6[346], stage0_6[347], stage0_6[348], stage0_6[349]},
      {stage0_7[327]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[57],stage1_8[112],stage1_7[139],stage1_6[168]}
   );
   gpc615_5 gpc313 (
      {stage0_6[350], stage0_6[351], stage0_6[352], stage0_6[353], stage0_6[354]},
      {stage0_7[328]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[58],stage1_8[113],stage1_7[140],stage1_6[169]}
   );
   gpc615_5 gpc314 (
      {stage0_6[355], stage0_6[356], stage0_6[357], stage0_6[358], stage0_6[359]},
      {stage0_7[329]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[59],stage1_8[114],stage1_7[141],stage1_6[170]}
   );
   gpc615_5 gpc315 (
      {stage0_6[360], stage0_6[361], stage0_6[362], stage0_6[363], stage0_6[364]},
      {stage0_7[330]},
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage1_10[6],stage1_9[60],stage1_8[115],stage1_7[142],stage1_6[171]}
   );
   gpc615_5 gpc316 (
      {stage0_6[365], stage0_6[366], stage0_6[367], stage0_6[368], stage0_6[369]},
      {stage0_7[331]},
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage1_10[7],stage1_9[61],stage1_8[116],stage1_7[143],stage1_6[172]}
   );
   gpc615_5 gpc317 (
      {stage0_6[370], stage0_6[371], stage0_6[372], stage0_6[373], stage0_6[374]},
      {stage0_7[332]},
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage1_10[8],stage1_9[62],stage1_8[117],stage1_7[144],stage1_6[173]}
   );
   gpc615_5 gpc318 (
      {stage0_6[375], stage0_6[376], stage0_6[377], stage0_6[378], stage0_6[379]},
      {stage0_7[333]},
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage1_10[9],stage1_9[63],stage1_8[118],stage1_7[145],stage1_6[174]}
   );
   gpc615_5 gpc319 (
      {stage0_6[380], stage0_6[381], stage0_6[382], stage0_6[383], stage0_6[384]},
      {stage0_7[334]},
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage1_10[10],stage1_9[64],stage1_8[119],stage1_7[146],stage1_6[175]}
   );
   gpc615_5 gpc320 (
      {stage0_6[385], stage0_6[386], stage0_6[387], stage0_6[388], stage0_6[389]},
      {stage0_7[335]},
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage1_10[11],stage1_9[65],stage1_8[120],stage1_7[147],stage1_6[176]}
   );
   gpc615_5 gpc321 (
      {stage0_6[390], stage0_6[391], stage0_6[392], stage0_6[393], stage0_6[394]},
      {stage0_7[336]},
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77]},
      {stage1_10[12],stage1_9[66],stage1_8[121],stage1_7[148],stage1_6[177]}
   );
   gpc615_5 gpc322 (
      {stage0_6[395], stage0_6[396], stage0_6[397], stage0_6[398], stage0_6[399]},
      {stage0_7[337]},
      {stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83]},
      {stage1_10[13],stage1_9[67],stage1_8[122],stage1_7[149],stage1_6[178]}
   );
   gpc615_5 gpc323 (
      {stage0_6[400], stage0_6[401], stage0_6[402], stage0_6[403], stage0_6[404]},
      {stage0_7[338]},
      {stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89]},
      {stage1_10[14],stage1_9[68],stage1_8[123],stage1_7[150],stage1_6[179]}
   );
   gpc615_5 gpc324 (
      {stage0_6[405], stage0_6[406], stage0_6[407], stage0_6[408], stage0_6[409]},
      {stage0_7[339]},
      {stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95]},
      {stage1_10[15],stage1_9[69],stage1_8[124],stage1_7[151],stage1_6[180]}
   );
   gpc615_5 gpc325 (
      {stage0_6[410], stage0_6[411], stage0_6[412], stage0_6[413], stage0_6[414]},
      {stage0_7[340]},
      {stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage1_10[16],stage1_9[70],stage1_8[125],stage1_7[152],stage1_6[181]}
   );
   gpc615_5 gpc326 (
      {stage0_6[415], stage0_6[416], stage0_6[417], stage0_6[418], stage0_6[419]},
      {stage0_7[341]},
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107]},
      {stage1_10[17],stage1_9[71],stage1_8[126],stage1_7[153],stage1_6[182]}
   );
   gpc615_5 gpc327 (
      {stage0_6[420], stage0_6[421], stage0_6[422], stage0_6[423], stage0_6[424]},
      {stage0_7[342]},
      {stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111], stage0_8[112], stage0_8[113]},
      {stage1_10[18],stage1_9[72],stage1_8[127],stage1_7[154],stage1_6[183]}
   );
   gpc615_5 gpc328 (
      {stage0_6[425], stage0_6[426], stage0_6[427], stage0_6[428], stage0_6[429]},
      {stage0_7[343]},
      {stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117], stage0_8[118], stage0_8[119]},
      {stage1_10[19],stage1_9[73],stage1_8[128],stage1_7[155],stage1_6[184]}
   );
   gpc615_5 gpc329 (
      {stage0_6[430], stage0_6[431], stage0_6[432], stage0_6[433], stage0_6[434]},
      {stage0_7[344]},
      {stage0_8[120], stage0_8[121], stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125]},
      {stage1_10[20],stage1_9[74],stage1_8[129],stage1_7[156],stage1_6[185]}
   );
   gpc615_5 gpc330 (
      {stage0_6[435], stage0_6[436], stage0_6[437], stage0_6[438], stage0_6[439]},
      {stage0_7[345]},
      {stage0_8[126], stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage1_10[21],stage1_9[75],stage1_8[130],stage1_7[157],stage1_6[186]}
   );
   gpc615_5 gpc331 (
      {stage0_6[440], stage0_6[441], stage0_6[442], stage0_6[443], stage0_6[444]},
      {stage0_7[346]},
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136], stage0_8[137]},
      {stage1_10[22],stage1_9[76],stage1_8[131],stage1_7[158],stage1_6[187]}
   );
   gpc615_5 gpc332 (
      {stage0_6[445], stage0_6[446], stage0_6[447], stage0_6[448], stage0_6[449]},
      {stage0_7[347]},
      {stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141], stage0_8[142], stage0_8[143]},
      {stage1_10[23],stage1_9[77],stage1_8[132],stage1_7[159],stage1_6[188]}
   );
   gpc615_5 gpc333 (
      {stage0_6[450], stage0_6[451], stage0_6[452], stage0_6[453], stage0_6[454]},
      {stage0_7[348]},
      {stage0_8[144], stage0_8[145], stage0_8[146], stage0_8[147], stage0_8[148], stage0_8[149]},
      {stage1_10[24],stage1_9[78],stage1_8[133],stage1_7[160],stage1_6[189]}
   );
   gpc615_5 gpc334 (
      {stage0_6[455], stage0_6[456], stage0_6[457], stage0_6[458], stage0_6[459]},
      {stage0_7[349]},
      {stage0_8[150], stage0_8[151], stage0_8[152], stage0_8[153], stage0_8[154], stage0_8[155]},
      {stage1_10[25],stage1_9[79],stage1_8[134],stage1_7[161],stage1_6[190]}
   );
   gpc615_5 gpc335 (
      {stage0_6[460], stage0_6[461], stage0_6[462], stage0_6[463], stage0_6[464]},
      {stage0_7[350]},
      {stage0_8[156], stage0_8[157], stage0_8[158], stage0_8[159], stage0_8[160], stage0_8[161]},
      {stage1_10[26],stage1_9[80],stage1_8[135],stage1_7[162],stage1_6[191]}
   );
   gpc615_5 gpc336 (
      {stage0_6[465], stage0_6[466], stage0_6[467], stage0_6[468], stage0_6[469]},
      {stage0_7[351]},
      {stage0_8[162], stage0_8[163], stage0_8[164], stage0_8[165], stage0_8[166], stage0_8[167]},
      {stage1_10[27],stage1_9[81],stage1_8[136],stage1_7[163],stage1_6[192]}
   );
   gpc615_5 gpc337 (
      {stage0_6[470], stage0_6[471], stage0_6[472], stage0_6[473], stage0_6[474]},
      {stage0_7[352]},
      {stage0_8[168], stage0_8[169], stage0_8[170], stage0_8[171], stage0_8[172], stage0_8[173]},
      {stage1_10[28],stage1_9[82],stage1_8[137],stage1_7[164],stage1_6[193]}
   );
   gpc615_5 gpc338 (
      {stage0_6[475], stage0_6[476], stage0_6[477], stage0_6[478], stage0_6[479]},
      {stage0_7[353]},
      {stage0_8[174], stage0_8[175], stage0_8[176], stage0_8[177], stage0_8[178], stage0_8[179]},
      {stage1_10[29],stage1_9[83],stage1_8[138],stage1_7[165],stage1_6[194]}
   );
   gpc615_5 gpc339 (
      {stage0_6[480], stage0_6[481], stage0_6[482], stage0_6[483], stage0_6[484]},
      {stage0_7[354]},
      {stage0_8[180], stage0_8[181], stage0_8[182], stage0_8[183], stage0_8[184], stage0_8[185]},
      {stage1_10[30],stage1_9[84],stage1_8[139],stage1_7[166],stage1_6[195]}
   );
   gpc615_5 gpc340 (
      {stage0_6[485], stage0_6[486], stage0_6[487], stage0_6[488], stage0_6[489]},
      {stage0_7[355]},
      {stage0_8[186], stage0_8[187], stage0_8[188], stage0_8[189], stage0_8[190], stage0_8[191]},
      {stage1_10[31],stage1_9[85],stage1_8[140],stage1_7[167],stage1_6[196]}
   );
   gpc615_5 gpc341 (
      {stage0_6[490], stage0_6[491], stage0_6[492], stage0_6[493], stage0_6[494]},
      {stage0_7[356]},
      {stage0_8[192], stage0_8[193], stage0_8[194], stage0_8[195], stage0_8[196], stage0_8[197]},
      {stage1_10[32],stage1_9[86],stage1_8[141],stage1_7[168],stage1_6[197]}
   );
   gpc615_5 gpc342 (
      {stage0_6[495], stage0_6[496], stage0_6[497], stage0_6[498], stage0_6[499]},
      {stage0_7[357]},
      {stage0_8[198], stage0_8[199], stage0_8[200], stage0_8[201], stage0_8[202], stage0_8[203]},
      {stage1_10[33],stage1_9[87],stage1_8[142],stage1_7[169],stage1_6[198]}
   );
   gpc615_5 gpc343 (
      {stage0_6[500], stage0_6[501], stage0_6[502], stage0_6[503], stage0_6[504]},
      {stage0_7[358]},
      {stage0_8[204], stage0_8[205], stage0_8[206], stage0_8[207], stage0_8[208], stage0_8[209]},
      {stage1_10[34],stage1_9[88],stage1_8[143],stage1_7[170],stage1_6[199]}
   );
   gpc606_5 gpc344 (
      {stage0_7[359], stage0_7[360], stage0_7[361], stage0_7[362], stage0_7[363], stage0_7[364]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[35],stage1_9[89],stage1_8[144],stage1_7[171]}
   );
   gpc606_5 gpc345 (
      {stage0_7[365], stage0_7[366], stage0_7[367], stage0_7[368], stage0_7[369], stage0_7[370]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[36],stage1_9[90],stage1_8[145],stage1_7[172]}
   );
   gpc606_5 gpc346 (
      {stage0_7[371], stage0_7[372], stage0_7[373], stage0_7[374], stage0_7[375], stage0_7[376]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[37],stage1_9[91],stage1_8[146],stage1_7[173]}
   );
   gpc606_5 gpc347 (
      {stage0_7[377], stage0_7[378], stage0_7[379], stage0_7[380], stage0_7[381], stage0_7[382]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[38],stage1_9[92],stage1_8[147],stage1_7[174]}
   );
   gpc606_5 gpc348 (
      {stage0_7[383], stage0_7[384], stage0_7[385], stage0_7[386], stage0_7[387], stage0_7[388]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[39],stage1_9[93],stage1_8[148],stage1_7[175]}
   );
   gpc606_5 gpc349 (
      {stage0_7[389], stage0_7[390], stage0_7[391], stage0_7[392], stage0_7[393], stage0_7[394]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[40],stage1_9[94],stage1_8[149],stage1_7[176]}
   );
   gpc606_5 gpc350 (
      {stage0_7[395], stage0_7[396], stage0_7[397], stage0_7[398], stage0_7[399], stage0_7[400]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[41],stage1_9[95],stage1_8[150],stage1_7[177]}
   );
   gpc606_5 gpc351 (
      {stage0_7[401], stage0_7[402], stage0_7[403], stage0_7[404], stage0_7[405], stage0_7[406]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[42],stage1_9[96],stage1_8[151],stage1_7[178]}
   );
   gpc606_5 gpc352 (
      {stage0_7[407], stage0_7[408], stage0_7[409], stage0_7[410], stage0_7[411], stage0_7[412]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[43],stage1_9[97],stage1_8[152],stage1_7[179]}
   );
   gpc606_5 gpc353 (
      {stage0_7[413], stage0_7[414], stage0_7[415], stage0_7[416], stage0_7[417], stage0_7[418]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[44],stage1_9[98],stage1_8[153],stage1_7[180]}
   );
   gpc606_5 gpc354 (
      {stage0_7[419], stage0_7[420], stage0_7[421], stage0_7[422], stage0_7[423], stage0_7[424]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[45],stage1_9[99],stage1_8[154],stage1_7[181]}
   );
   gpc606_5 gpc355 (
      {stage0_7[425], stage0_7[426], stage0_7[427], stage0_7[428], stage0_7[429], stage0_7[430]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[46],stage1_9[100],stage1_8[155],stage1_7[182]}
   );
   gpc606_5 gpc356 (
      {stage0_7[431], stage0_7[432], stage0_7[433], stage0_7[434], stage0_7[435], stage0_7[436]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[47],stage1_9[101],stage1_8[156],stage1_7[183]}
   );
   gpc606_5 gpc357 (
      {stage0_7[437], stage0_7[438], stage0_7[439], stage0_7[440], stage0_7[441], stage0_7[442]},
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83]},
      {stage1_11[13],stage1_10[48],stage1_9[102],stage1_8[157],stage1_7[184]}
   );
   gpc606_5 gpc358 (
      {stage0_7[443], stage0_7[444], stage0_7[445], stage0_7[446], stage0_7[447], stage0_7[448]},
      {stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89]},
      {stage1_11[14],stage1_10[49],stage1_9[103],stage1_8[158],stage1_7[185]}
   );
   gpc606_5 gpc359 (
      {stage0_7[449], stage0_7[450], stage0_7[451], stage0_7[452], stage0_7[453], stage0_7[454]},
      {stage0_9[90], stage0_9[91], stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95]},
      {stage1_11[15],stage1_10[50],stage1_9[104],stage1_8[159],stage1_7[186]}
   );
   gpc606_5 gpc360 (
      {stage0_7[455], stage0_7[456], stage0_7[457], stage0_7[458], stage0_7[459], stage0_7[460]},
      {stage0_9[96], stage0_9[97], stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101]},
      {stage1_11[16],stage1_10[51],stage1_9[105],stage1_8[160],stage1_7[187]}
   );
   gpc615_5 gpc361 (
      {stage0_7[461], stage0_7[462], stage0_7[463], stage0_7[464], stage0_7[465]},
      {stage0_8[210]},
      {stage0_9[102], stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage1_11[17],stage1_10[52],stage1_9[106],stage1_8[161],stage1_7[188]}
   );
   gpc615_5 gpc362 (
      {stage0_7[466], stage0_7[467], stage0_7[468], stage0_7[469], stage0_7[470]},
      {stage0_8[211]},
      {stage0_9[108], stage0_9[109], stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113]},
      {stage1_11[18],stage1_10[53],stage1_9[107],stage1_8[162],stage1_7[189]}
   );
   gpc615_5 gpc363 (
      {stage0_7[471], stage0_7[472], stage0_7[473], stage0_7[474], stage0_7[475]},
      {stage0_8[212]},
      {stage0_9[114], stage0_9[115], stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119]},
      {stage1_11[19],stage1_10[54],stage1_9[108],stage1_8[163],stage1_7[190]}
   );
   gpc615_5 gpc364 (
      {stage0_7[476], stage0_7[477], stage0_7[478], stage0_7[479], stage0_7[480]},
      {stage0_8[213]},
      {stage0_9[120], stage0_9[121], stage0_9[122], stage0_9[123], stage0_9[124], stage0_9[125]},
      {stage1_11[20],stage1_10[55],stage1_9[109],stage1_8[164],stage1_7[191]}
   );
   gpc615_5 gpc365 (
      {stage0_7[481], stage0_7[482], stage0_7[483], stage0_7[484], stage0_7[485]},
      {stage0_8[214]},
      {stage0_9[126], stage0_9[127], stage0_9[128], stage0_9[129], stage0_9[130], stage0_9[131]},
      {stage1_11[21],stage1_10[56],stage1_9[110],stage1_8[165],stage1_7[192]}
   );
   gpc615_5 gpc366 (
      {stage0_7[486], stage0_7[487], stage0_7[488], stage0_7[489], stage0_7[490]},
      {stage0_8[215]},
      {stage0_9[132], stage0_9[133], stage0_9[134], stage0_9[135], stage0_9[136], stage0_9[137]},
      {stage1_11[22],stage1_10[57],stage1_9[111],stage1_8[166],stage1_7[193]}
   );
   gpc615_5 gpc367 (
      {stage0_7[491], stage0_7[492], stage0_7[493], stage0_7[494], stage0_7[495]},
      {stage0_8[216]},
      {stage0_9[138], stage0_9[139], stage0_9[140], stage0_9[141], stage0_9[142], stage0_9[143]},
      {stage1_11[23],stage1_10[58],stage1_9[112],stage1_8[167],stage1_7[194]}
   );
   gpc615_5 gpc368 (
      {stage0_7[496], stage0_7[497], stage0_7[498], stage0_7[499], stage0_7[500]},
      {stage0_8[217]},
      {stage0_9[144], stage0_9[145], stage0_9[146], stage0_9[147], stage0_9[148], stage0_9[149]},
      {stage1_11[24],stage1_10[59],stage1_9[113],stage1_8[168],stage1_7[195]}
   );
   gpc606_5 gpc369 (
      {stage0_8[218], stage0_8[219], stage0_8[220], stage0_8[221], stage0_8[222], stage0_8[223]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[25],stage1_10[60],stage1_9[114],stage1_8[169]}
   );
   gpc606_5 gpc370 (
      {stage0_8[224], stage0_8[225], stage0_8[226], stage0_8[227], stage0_8[228], stage0_8[229]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[26],stage1_10[61],stage1_9[115],stage1_8[170]}
   );
   gpc606_5 gpc371 (
      {stage0_8[230], stage0_8[231], stage0_8[232], stage0_8[233], stage0_8[234], stage0_8[235]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[27],stage1_10[62],stage1_9[116],stage1_8[171]}
   );
   gpc606_5 gpc372 (
      {stage0_8[236], stage0_8[237], stage0_8[238], stage0_8[239], stage0_8[240], stage0_8[241]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[28],stage1_10[63],stage1_9[117],stage1_8[172]}
   );
   gpc606_5 gpc373 (
      {stage0_8[242], stage0_8[243], stage0_8[244], stage0_8[245], stage0_8[246], stage0_8[247]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[29],stage1_10[64],stage1_9[118],stage1_8[173]}
   );
   gpc606_5 gpc374 (
      {stage0_8[248], stage0_8[249], stage0_8[250], stage0_8[251], stage0_8[252], stage0_8[253]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[30],stage1_10[65],stage1_9[119],stage1_8[174]}
   );
   gpc606_5 gpc375 (
      {stage0_8[254], stage0_8[255], stage0_8[256], stage0_8[257], stage0_8[258], stage0_8[259]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[31],stage1_10[66],stage1_9[120],stage1_8[175]}
   );
   gpc606_5 gpc376 (
      {stage0_8[260], stage0_8[261], stage0_8[262], stage0_8[263], stage0_8[264], stage0_8[265]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[32],stage1_10[67],stage1_9[121],stage1_8[176]}
   );
   gpc606_5 gpc377 (
      {stage0_8[266], stage0_8[267], stage0_8[268], stage0_8[269], stage0_8[270], stage0_8[271]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[33],stage1_10[68],stage1_9[122],stage1_8[177]}
   );
   gpc606_5 gpc378 (
      {stage0_8[272], stage0_8[273], stage0_8[274], stage0_8[275], stage0_8[276], stage0_8[277]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[34],stage1_10[69],stage1_9[123],stage1_8[178]}
   );
   gpc606_5 gpc379 (
      {stage0_8[278], stage0_8[279], stage0_8[280], stage0_8[281], stage0_8[282], stage0_8[283]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[35],stage1_10[70],stage1_9[124],stage1_8[179]}
   );
   gpc606_5 gpc380 (
      {stage0_8[284], stage0_8[285], stage0_8[286], stage0_8[287], stage0_8[288], stage0_8[289]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[36],stage1_10[71],stage1_9[125],stage1_8[180]}
   );
   gpc606_5 gpc381 (
      {stage0_8[290], stage0_8[291], stage0_8[292], stage0_8[293], stage0_8[294], stage0_8[295]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[37],stage1_10[72],stage1_9[126],stage1_8[181]}
   );
   gpc606_5 gpc382 (
      {stage0_8[296], stage0_8[297], stage0_8[298], stage0_8[299], stage0_8[300], stage0_8[301]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[38],stage1_10[73],stage1_9[127],stage1_8[182]}
   );
   gpc606_5 gpc383 (
      {stage0_8[302], stage0_8[303], stage0_8[304], stage0_8[305], stage0_8[306], stage0_8[307]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[39],stage1_10[74],stage1_9[128],stage1_8[183]}
   );
   gpc606_5 gpc384 (
      {stage0_8[308], stage0_8[309], stage0_8[310], stage0_8[311], stage0_8[312], stage0_8[313]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[40],stage1_10[75],stage1_9[129],stage1_8[184]}
   );
   gpc606_5 gpc385 (
      {stage0_8[314], stage0_8[315], stage0_8[316], stage0_8[317], stage0_8[318], stage0_8[319]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[41],stage1_10[76],stage1_9[130],stage1_8[185]}
   );
   gpc606_5 gpc386 (
      {stage0_8[320], stage0_8[321], stage0_8[322], stage0_8[323], stage0_8[324], stage0_8[325]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[42],stage1_10[77],stage1_9[131],stage1_8[186]}
   );
   gpc606_5 gpc387 (
      {stage0_8[326], stage0_8[327], stage0_8[328], stage0_8[329], stage0_8[330], stage0_8[331]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[43],stage1_10[78],stage1_9[132],stage1_8[187]}
   );
   gpc606_5 gpc388 (
      {stage0_8[332], stage0_8[333], stage0_8[334], stage0_8[335], stage0_8[336], stage0_8[337]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[44],stage1_10[79],stage1_9[133],stage1_8[188]}
   );
   gpc606_5 gpc389 (
      {stage0_8[338], stage0_8[339], stage0_8[340], stage0_8[341], stage0_8[342], stage0_8[343]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[45],stage1_10[80],stage1_9[134],stage1_8[189]}
   );
   gpc606_5 gpc390 (
      {stage0_8[344], stage0_8[345], stage0_8[346], stage0_8[347], stage0_8[348], stage0_8[349]},
      {stage0_10[126], stage0_10[127], stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131]},
      {stage1_12[21],stage1_11[46],stage1_10[81],stage1_9[135],stage1_8[190]}
   );
   gpc606_5 gpc391 (
      {stage0_8[350], stage0_8[351], stage0_8[352], stage0_8[353], stage0_8[354], stage0_8[355]},
      {stage0_10[132], stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage1_12[22],stage1_11[47],stage1_10[82],stage1_9[136],stage1_8[191]}
   );
   gpc606_5 gpc392 (
      {stage0_8[356], stage0_8[357], stage0_8[358], stage0_8[359], stage0_8[360], stage0_8[361]},
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142], stage0_10[143]},
      {stage1_12[23],stage1_11[48],stage1_10[83],stage1_9[137],stage1_8[192]}
   );
   gpc606_5 gpc393 (
      {stage0_8[362], stage0_8[363], stage0_8[364], stage0_8[365], stage0_8[366], stage0_8[367]},
      {stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147], stage0_10[148], stage0_10[149]},
      {stage1_12[24],stage1_11[49],stage1_10[84],stage1_9[138],stage1_8[193]}
   );
   gpc606_5 gpc394 (
      {stage0_8[368], stage0_8[369], stage0_8[370], stage0_8[371], stage0_8[372], stage0_8[373]},
      {stage0_10[150], stage0_10[151], stage0_10[152], stage0_10[153], stage0_10[154], stage0_10[155]},
      {stage1_12[25],stage1_11[50],stage1_10[85],stage1_9[139],stage1_8[194]}
   );
   gpc606_5 gpc395 (
      {stage0_8[374], stage0_8[375], stage0_8[376], stage0_8[377], stage0_8[378], stage0_8[379]},
      {stage0_10[156], stage0_10[157], stage0_10[158], stage0_10[159], stage0_10[160], stage0_10[161]},
      {stage1_12[26],stage1_11[51],stage1_10[86],stage1_9[140],stage1_8[195]}
   );
   gpc606_5 gpc396 (
      {stage0_8[380], stage0_8[381], stage0_8[382], stage0_8[383], stage0_8[384], stage0_8[385]},
      {stage0_10[162], stage0_10[163], stage0_10[164], stage0_10[165], stage0_10[166], stage0_10[167]},
      {stage1_12[27],stage1_11[52],stage1_10[87],stage1_9[141],stage1_8[196]}
   );
   gpc606_5 gpc397 (
      {stage0_8[386], stage0_8[387], stage0_8[388], stage0_8[389], stage0_8[390], stage0_8[391]},
      {stage0_10[168], stage0_10[169], stage0_10[170], stage0_10[171], stage0_10[172], stage0_10[173]},
      {stage1_12[28],stage1_11[53],stage1_10[88],stage1_9[142],stage1_8[197]}
   );
   gpc606_5 gpc398 (
      {stage0_8[392], stage0_8[393], stage0_8[394], stage0_8[395], stage0_8[396], stage0_8[397]},
      {stage0_10[174], stage0_10[175], stage0_10[176], stage0_10[177], stage0_10[178], stage0_10[179]},
      {stage1_12[29],stage1_11[54],stage1_10[89],stage1_9[143],stage1_8[198]}
   );
   gpc606_5 gpc399 (
      {stage0_8[398], stage0_8[399], stage0_8[400], stage0_8[401], stage0_8[402], stage0_8[403]},
      {stage0_10[180], stage0_10[181], stage0_10[182], stage0_10[183], stage0_10[184], stage0_10[185]},
      {stage1_12[30],stage1_11[55],stage1_10[90],stage1_9[144],stage1_8[199]}
   );
   gpc606_5 gpc400 (
      {stage0_8[404], stage0_8[405], stage0_8[406], stage0_8[407], stage0_8[408], stage0_8[409]},
      {stage0_10[186], stage0_10[187], stage0_10[188], stage0_10[189], stage0_10[190], stage0_10[191]},
      {stage1_12[31],stage1_11[56],stage1_10[91],stage1_9[145],stage1_8[200]}
   );
   gpc606_5 gpc401 (
      {stage0_8[410], stage0_8[411], stage0_8[412], stage0_8[413], stage0_8[414], stage0_8[415]},
      {stage0_10[192], stage0_10[193], stage0_10[194], stage0_10[195], stage0_10[196], stage0_10[197]},
      {stage1_12[32],stage1_11[57],stage1_10[92],stage1_9[146],stage1_8[201]}
   );
   gpc606_5 gpc402 (
      {stage0_8[416], stage0_8[417], stage0_8[418], stage0_8[419], stage0_8[420], stage0_8[421]},
      {stage0_10[198], stage0_10[199], stage0_10[200], stage0_10[201], stage0_10[202], stage0_10[203]},
      {stage1_12[33],stage1_11[58],stage1_10[93],stage1_9[147],stage1_8[202]}
   );
   gpc606_5 gpc403 (
      {stage0_8[422], stage0_8[423], stage0_8[424], stage0_8[425], stage0_8[426], stage0_8[427]},
      {stage0_10[204], stage0_10[205], stage0_10[206], stage0_10[207], stage0_10[208], stage0_10[209]},
      {stage1_12[34],stage1_11[59],stage1_10[94],stage1_9[148],stage1_8[203]}
   );
   gpc606_5 gpc404 (
      {stage0_8[428], stage0_8[429], stage0_8[430], stage0_8[431], stage0_8[432], stage0_8[433]},
      {stage0_10[210], stage0_10[211], stage0_10[212], stage0_10[213], stage0_10[214], stage0_10[215]},
      {stage1_12[35],stage1_11[60],stage1_10[95],stage1_9[149],stage1_8[204]}
   );
   gpc606_5 gpc405 (
      {stage0_8[434], stage0_8[435], stage0_8[436], stage0_8[437], stage0_8[438], stage0_8[439]},
      {stage0_10[216], stage0_10[217], stage0_10[218], stage0_10[219], stage0_10[220], stage0_10[221]},
      {stage1_12[36],stage1_11[61],stage1_10[96],stage1_9[150],stage1_8[205]}
   );
   gpc606_5 gpc406 (
      {stage0_8[440], stage0_8[441], stage0_8[442], stage0_8[443], stage0_8[444], stage0_8[445]},
      {stage0_10[222], stage0_10[223], stage0_10[224], stage0_10[225], stage0_10[226], stage0_10[227]},
      {stage1_12[37],stage1_11[62],stage1_10[97],stage1_9[151],stage1_8[206]}
   );
   gpc606_5 gpc407 (
      {stage0_8[446], stage0_8[447], stage0_8[448], stage0_8[449], stage0_8[450], stage0_8[451]},
      {stage0_10[228], stage0_10[229], stage0_10[230], stage0_10[231], stage0_10[232], stage0_10[233]},
      {stage1_12[38],stage1_11[63],stage1_10[98],stage1_9[152],stage1_8[207]}
   );
   gpc606_5 gpc408 (
      {stage0_8[452], stage0_8[453], stage0_8[454], stage0_8[455], stage0_8[456], stage0_8[457]},
      {stage0_10[234], stage0_10[235], stage0_10[236], stage0_10[237], stage0_10[238], stage0_10[239]},
      {stage1_12[39],stage1_11[64],stage1_10[99],stage1_9[153],stage1_8[208]}
   );
   gpc606_5 gpc409 (
      {stage0_8[458], stage0_8[459], stage0_8[460], stage0_8[461], stage0_8[462], stage0_8[463]},
      {stage0_10[240], stage0_10[241], stage0_10[242], stage0_10[243], stage0_10[244], stage0_10[245]},
      {stage1_12[40],stage1_11[65],stage1_10[100],stage1_9[154],stage1_8[209]}
   );
   gpc606_5 gpc410 (
      {stage0_8[464], stage0_8[465], stage0_8[466], stage0_8[467], stage0_8[468], stage0_8[469]},
      {stage0_10[246], stage0_10[247], stage0_10[248], stage0_10[249], stage0_10[250], stage0_10[251]},
      {stage1_12[41],stage1_11[66],stage1_10[101],stage1_9[155],stage1_8[210]}
   );
   gpc606_5 gpc411 (
      {stage0_8[470], stage0_8[471], stage0_8[472], stage0_8[473], stage0_8[474], stage0_8[475]},
      {stage0_10[252], stage0_10[253], stage0_10[254], stage0_10[255], stage0_10[256], stage0_10[257]},
      {stage1_12[42],stage1_11[67],stage1_10[102],stage1_9[156],stage1_8[211]}
   );
   gpc606_5 gpc412 (
      {stage0_8[476], stage0_8[477], stage0_8[478], stage0_8[479], stage0_8[480], stage0_8[481]},
      {stage0_10[258], stage0_10[259], stage0_10[260], stage0_10[261], stage0_10[262], stage0_10[263]},
      {stage1_12[43],stage1_11[68],stage1_10[103],stage1_9[157],stage1_8[212]}
   );
   gpc606_5 gpc413 (
      {stage0_8[482], stage0_8[483], stage0_8[484], stage0_8[485], stage0_8[486], stage0_8[487]},
      {stage0_10[264], stage0_10[265], stage0_10[266], stage0_10[267], stage0_10[268], stage0_10[269]},
      {stage1_12[44],stage1_11[69],stage1_10[104],stage1_9[158],stage1_8[213]}
   );
   gpc606_5 gpc414 (
      {stage0_8[488], stage0_8[489], stage0_8[490], stage0_8[491], stage0_8[492], stage0_8[493]},
      {stage0_10[270], stage0_10[271], stage0_10[272], stage0_10[273], stage0_10[274], stage0_10[275]},
      {stage1_12[45],stage1_11[70],stage1_10[105],stage1_9[159],stage1_8[214]}
   );
   gpc606_5 gpc415 (
      {stage0_8[494], stage0_8[495], stage0_8[496], stage0_8[497], stage0_8[498], stage0_8[499]},
      {stage0_10[276], stage0_10[277], stage0_10[278], stage0_10[279], stage0_10[280], stage0_10[281]},
      {stage1_12[46],stage1_11[71],stage1_10[106],stage1_9[160],stage1_8[215]}
   );
   gpc606_5 gpc416 (
      {stage0_8[500], stage0_8[501], stage0_8[502], stage0_8[503], stage0_8[504], stage0_8[505]},
      {stage0_10[282], stage0_10[283], stage0_10[284], stage0_10[285], stage0_10[286], stage0_10[287]},
      {stage1_12[47],stage1_11[72],stage1_10[107],stage1_9[161],stage1_8[216]}
   );
   gpc606_5 gpc417 (
      {stage0_8[506], stage0_8[507], stage0_8[508], stage0_8[509], stage0_8[510], stage0_8[511]},
      {stage0_10[288], stage0_10[289], stage0_10[290], stage0_10[291], stage0_10[292], stage0_10[293]},
      {stage1_12[48],stage1_11[73],stage1_10[108],stage1_9[162],stage1_8[217]}
   );
   gpc606_5 gpc418 (
      {stage0_9[150], stage0_9[151], stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[49],stage1_11[74],stage1_10[109],stage1_9[163]}
   );
   gpc615_5 gpc419 (
      {stage0_9[156], stage0_9[157], stage0_9[158], stage0_9[159], stage0_9[160]},
      {stage0_10[294]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[50],stage1_11[75],stage1_10[110],stage1_9[164]}
   );
   gpc615_5 gpc420 (
      {stage0_9[161], stage0_9[162], stage0_9[163], stage0_9[164], stage0_9[165]},
      {stage0_10[295]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[51],stage1_11[76],stage1_10[111],stage1_9[165]}
   );
   gpc615_5 gpc421 (
      {stage0_9[166], stage0_9[167], stage0_9[168], stage0_9[169], stage0_9[170]},
      {stage0_10[296]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[52],stage1_11[77],stage1_10[112],stage1_9[166]}
   );
   gpc615_5 gpc422 (
      {stage0_9[171], stage0_9[172], stage0_9[173], stage0_9[174], stage0_9[175]},
      {stage0_10[297]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[53],stage1_11[78],stage1_10[113],stage1_9[167]}
   );
   gpc615_5 gpc423 (
      {stage0_9[176], stage0_9[177], stage0_9[178], stage0_9[179], stage0_9[180]},
      {stage0_10[298]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[54],stage1_11[79],stage1_10[114],stage1_9[168]}
   );
   gpc615_5 gpc424 (
      {stage0_9[181], stage0_9[182], stage0_9[183], stage0_9[184], stage0_9[185]},
      {stage0_10[299]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[55],stage1_11[80],stage1_10[115],stage1_9[169]}
   );
   gpc615_5 gpc425 (
      {stage0_9[186], stage0_9[187], stage0_9[188], stage0_9[189], stage0_9[190]},
      {stage0_10[300]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[56],stage1_11[81],stage1_10[116],stage1_9[170]}
   );
   gpc615_5 gpc426 (
      {stage0_9[191], stage0_9[192], stage0_9[193], stage0_9[194], stage0_9[195]},
      {stage0_10[301]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[57],stage1_11[82],stage1_10[117],stage1_9[171]}
   );
   gpc615_5 gpc427 (
      {stage0_9[196], stage0_9[197], stage0_9[198], stage0_9[199], stage0_9[200]},
      {stage0_10[302]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[58],stage1_11[83],stage1_10[118],stage1_9[172]}
   );
   gpc615_5 gpc428 (
      {stage0_9[201], stage0_9[202], stage0_9[203], stage0_9[204], stage0_9[205]},
      {stage0_10[303]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[59],stage1_11[84],stage1_10[119],stage1_9[173]}
   );
   gpc615_5 gpc429 (
      {stage0_9[206], stage0_9[207], stage0_9[208], stage0_9[209], stage0_9[210]},
      {stage0_10[304]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[60],stage1_11[85],stage1_10[120],stage1_9[174]}
   );
   gpc615_5 gpc430 (
      {stage0_9[211], stage0_9[212], stage0_9[213], stage0_9[214], stage0_9[215]},
      {stage0_10[305]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[61],stage1_11[86],stage1_10[121],stage1_9[175]}
   );
   gpc615_5 gpc431 (
      {stage0_9[216], stage0_9[217], stage0_9[218], stage0_9[219], stage0_9[220]},
      {stage0_10[306]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[62],stage1_11[87],stage1_10[122],stage1_9[176]}
   );
   gpc615_5 gpc432 (
      {stage0_9[221], stage0_9[222], stage0_9[223], stage0_9[224], stage0_9[225]},
      {stage0_10[307]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[63],stage1_11[88],stage1_10[123],stage1_9[177]}
   );
   gpc615_5 gpc433 (
      {stage0_9[226], stage0_9[227], stage0_9[228], stage0_9[229], stage0_9[230]},
      {stage0_10[308]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[64],stage1_11[89],stage1_10[124],stage1_9[178]}
   );
   gpc615_5 gpc434 (
      {stage0_9[231], stage0_9[232], stage0_9[233], stage0_9[234], stage0_9[235]},
      {stage0_10[309]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[65],stage1_11[90],stage1_10[125],stage1_9[179]}
   );
   gpc615_5 gpc435 (
      {stage0_9[236], stage0_9[237], stage0_9[238], stage0_9[239], stage0_9[240]},
      {stage0_10[310]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[66],stage1_11[91],stage1_10[126],stage1_9[180]}
   );
   gpc615_5 gpc436 (
      {stage0_9[241], stage0_9[242], stage0_9[243], stage0_9[244], stage0_9[245]},
      {stage0_10[311]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[67],stage1_11[92],stage1_10[127],stage1_9[181]}
   );
   gpc615_5 gpc437 (
      {stage0_9[246], stage0_9[247], stage0_9[248], stage0_9[249], stage0_9[250]},
      {stage0_10[312]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[68],stage1_11[93],stage1_10[128],stage1_9[182]}
   );
   gpc615_5 gpc438 (
      {stage0_9[251], stage0_9[252], stage0_9[253], stage0_9[254], stage0_9[255]},
      {stage0_10[313]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[69],stage1_11[94],stage1_10[129],stage1_9[183]}
   );
   gpc615_5 gpc439 (
      {stage0_9[256], stage0_9[257], stage0_9[258], stage0_9[259], stage0_9[260]},
      {stage0_10[314]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[70],stage1_11[95],stage1_10[130],stage1_9[184]}
   );
   gpc615_5 gpc440 (
      {stage0_9[261], stage0_9[262], stage0_9[263], stage0_9[264], stage0_9[265]},
      {stage0_10[315]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[71],stage1_11[96],stage1_10[131],stage1_9[185]}
   );
   gpc615_5 gpc441 (
      {stage0_9[266], stage0_9[267], stage0_9[268], stage0_9[269], stage0_9[270]},
      {stage0_10[316]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[72],stage1_11[97],stage1_10[132],stage1_9[186]}
   );
   gpc615_5 gpc442 (
      {stage0_9[271], stage0_9[272], stage0_9[273], stage0_9[274], stage0_9[275]},
      {stage0_10[317]},
      {stage0_11[144], stage0_11[145], stage0_11[146], stage0_11[147], stage0_11[148], stage0_11[149]},
      {stage1_13[24],stage1_12[73],stage1_11[98],stage1_10[133],stage1_9[187]}
   );
   gpc615_5 gpc443 (
      {stage0_9[276], stage0_9[277], stage0_9[278], stage0_9[279], stage0_9[280]},
      {stage0_10[318]},
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage1_13[25],stage1_12[74],stage1_11[99],stage1_10[134],stage1_9[188]}
   );
   gpc615_5 gpc444 (
      {stage0_9[281], stage0_9[282], stage0_9[283], stage0_9[284], stage0_9[285]},
      {stage0_10[319]},
      {stage0_11[156], stage0_11[157], stage0_11[158], stage0_11[159], stage0_11[160], stage0_11[161]},
      {stage1_13[26],stage1_12[75],stage1_11[100],stage1_10[135],stage1_9[189]}
   );
   gpc615_5 gpc445 (
      {stage0_9[286], stage0_9[287], stage0_9[288], stage0_9[289], stage0_9[290]},
      {stage0_10[320]},
      {stage0_11[162], stage0_11[163], stage0_11[164], stage0_11[165], stage0_11[166], stage0_11[167]},
      {stage1_13[27],stage1_12[76],stage1_11[101],stage1_10[136],stage1_9[190]}
   );
   gpc615_5 gpc446 (
      {stage0_9[291], stage0_9[292], stage0_9[293], stage0_9[294], stage0_9[295]},
      {stage0_10[321]},
      {stage0_11[168], stage0_11[169], stage0_11[170], stage0_11[171], stage0_11[172], stage0_11[173]},
      {stage1_13[28],stage1_12[77],stage1_11[102],stage1_10[137],stage1_9[191]}
   );
   gpc615_5 gpc447 (
      {stage0_9[296], stage0_9[297], stage0_9[298], stage0_9[299], stage0_9[300]},
      {stage0_10[322]},
      {stage0_11[174], stage0_11[175], stage0_11[176], stage0_11[177], stage0_11[178], stage0_11[179]},
      {stage1_13[29],stage1_12[78],stage1_11[103],stage1_10[138],stage1_9[192]}
   );
   gpc615_5 gpc448 (
      {stage0_9[301], stage0_9[302], stage0_9[303], stage0_9[304], stage0_9[305]},
      {stage0_10[323]},
      {stage0_11[180], stage0_11[181], stage0_11[182], stage0_11[183], stage0_11[184], stage0_11[185]},
      {stage1_13[30],stage1_12[79],stage1_11[104],stage1_10[139],stage1_9[193]}
   );
   gpc615_5 gpc449 (
      {stage0_9[306], stage0_9[307], stage0_9[308], stage0_9[309], stage0_9[310]},
      {stage0_10[324]},
      {stage0_11[186], stage0_11[187], stage0_11[188], stage0_11[189], stage0_11[190], stage0_11[191]},
      {stage1_13[31],stage1_12[80],stage1_11[105],stage1_10[140],stage1_9[194]}
   );
   gpc615_5 gpc450 (
      {stage0_9[311], stage0_9[312], stage0_9[313], stage0_9[314], stage0_9[315]},
      {stage0_10[325]},
      {stage0_11[192], stage0_11[193], stage0_11[194], stage0_11[195], stage0_11[196], stage0_11[197]},
      {stage1_13[32],stage1_12[81],stage1_11[106],stage1_10[141],stage1_9[195]}
   );
   gpc615_5 gpc451 (
      {stage0_9[316], stage0_9[317], stage0_9[318], stage0_9[319], stage0_9[320]},
      {stage0_10[326]},
      {stage0_11[198], stage0_11[199], stage0_11[200], stage0_11[201], stage0_11[202], stage0_11[203]},
      {stage1_13[33],stage1_12[82],stage1_11[107],stage1_10[142],stage1_9[196]}
   );
   gpc615_5 gpc452 (
      {stage0_9[321], stage0_9[322], stage0_9[323], stage0_9[324], stage0_9[325]},
      {stage0_10[327]},
      {stage0_11[204], stage0_11[205], stage0_11[206], stage0_11[207], stage0_11[208], stage0_11[209]},
      {stage1_13[34],stage1_12[83],stage1_11[108],stage1_10[143],stage1_9[197]}
   );
   gpc615_5 gpc453 (
      {stage0_9[326], stage0_9[327], stage0_9[328], stage0_9[329], stage0_9[330]},
      {stage0_10[328]},
      {stage0_11[210], stage0_11[211], stage0_11[212], stage0_11[213], stage0_11[214], stage0_11[215]},
      {stage1_13[35],stage1_12[84],stage1_11[109],stage1_10[144],stage1_9[198]}
   );
   gpc615_5 gpc454 (
      {stage0_9[331], stage0_9[332], stage0_9[333], stage0_9[334], stage0_9[335]},
      {stage0_10[329]},
      {stage0_11[216], stage0_11[217], stage0_11[218], stage0_11[219], stage0_11[220], stage0_11[221]},
      {stage1_13[36],stage1_12[85],stage1_11[110],stage1_10[145],stage1_9[199]}
   );
   gpc615_5 gpc455 (
      {stage0_9[336], stage0_9[337], stage0_9[338], stage0_9[339], stage0_9[340]},
      {stage0_10[330]},
      {stage0_11[222], stage0_11[223], stage0_11[224], stage0_11[225], stage0_11[226], stage0_11[227]},
      {stage1_13[37],stage1_12[86],stage1_11[111],stage1_10[146],stage1_9[200]}
   );
   gpc615_5 gpc456 (
      {stage0_9[341], stage0_9[342], stage0_9[343], stage0_9[344], stage0_9[345]},
      {stage0_10[331]},
      {stage0_11[228], stage0_11[229], stage0_11[230], stage0_11[231], stage0_11[232], stage0_11[233]},
      {stage1_13[38],stage1_12[87],stage1_11[112],stage1_10[147],stage1_9[201]}
   );
   gpc615_5 gpc457 (
      {stage0_9[346], stage0_9[347], stage0_9[348], stage0_9[349], stage0_9[350]},
      {stage0_10[332]},
      {stage0_11[234], stage0_11[235], stage0_11[236], stage0_11[237], stage0_11[238], stage0_11[239]},
      {stage1_13[39],stage1_12[88],stage1_11[113],stage1_10[148],stage1_9[202]}
   );
   gpc615_5 gpc458 (
      {stage0_9[351], stage0_9[352], stage0_9[353], stage0_9[354], stage0_9[355]},
      {stage0_10[333]},
      {stage0_11[240], stage0_11[241], stage0_11[242], stage0_11[243], stage0_11[244], stage0_11[245]},
      {stage1_13[40],stage1_12[89],stage1_11[114],stage1_10[149],stage1_9[203]}
   );
   gpc615_5 gpc459 (
      {stage0_9[356], stage0_9[357], stage0_9[358], stage0_9[359], stage0_9[360]},
      {stage0_10[334]},
      {stage0_11[246], stage0_11[247], stage0_11[248], stage0_11[249], stage0_11[250], stage0_11[251]},
      {stage1_13[41],stage1_12[90],stage1_11[115],stage1_10[150],stage1_9[204]}
   );
   gpc615_5 gpc460 (
      {stage0_9[361], stage0_9[362], stage0_9[363], stage0_9[364], stage0_9[365]},
      {stage0_10[335]},
      {stage0_11[252], stage0_11[253], stage0_11[254], stage0_11[255], stage0_11[256], stage0_11[257]},
      {stage1_13[42],stage1_12[91],stage1_11[116],stage1_10[151],stage1_9[205]}
   );
   gpc615_5 gpc461 (
      {stage0_9[366], stage0_9[367], stage0_9[368], stage0_9[369], stage0_9[370]},
      {stage0_10[336]},
      {stage0_11[258], stage0_11[259], stage0_11[260], stage0_11[261], stage0_11[262], stage0_11[263]},
      {stage1_13[43],stage1_12[92],stage1_11[117],stage1_10[152],stage1_9[206]}
   );
   gpc615_5 gpc462 (
      {stage0_9[371], stage0_9[372], stage0_9[373], stage0_9[374], stage0_9[375]},
      {stage0_10[337]},
      {stage0_11[264], stage0_11[265], stage0_11[266], stage0_11[267], stage0_11[268], stage0_11[269]},
      {stage1_13[44],stage1_12[93],stage1_11[118],stage1_10[153],stage1_9[207]}
   );
   gpc615_5 gpc463 (
      {stage0_9[376], stage0_9[377], stage0_9[378], stage0_9[379], stage0_9[380]},
      {stage0_10[338]},
      {stage0_11[270], stage0_11[271], stage0_11[272], stage0_11[273], stage0_11[274], stage0_11[275]},
      {stage1_13[45],stage1_12[94],stage1_11[119],stage1_10[154],stage1_9[208]}
   );
   gpc615_5 gpc464 (
      {stage0_9[381], stage0_9[382], stage0_9[383], stage0_9[384], stage0_9[385]},
      {stage0_10[339]},
      {stage0_11[276], stage0_11[277], stage0_11[278], stage0_11[279], stage0_11[280], stage0_11[281]},
      {stage1_13[46],stage1_12[95],stage1_11[120],stage1_10[155],stage1_9[209]}
   );
   gpc615_5 gpc465 (
      {stage0_9[386], stage0_9[387], stage0_9[388], stage0_9[389], stage0_9[390]},
      {stage0_10[340]},
      {stage0_11[282], stage0_11[283], stage0_11[284], stage0_11[285], stage0_11[286], stage0_11[287]},
      {stage1_13[47],stage1_12[96],stage1_11[121],stage1_10[156],stage1_9[210]}
   );
   gpc615_5 gpc466 (
      {stage0_9[391], stage0_9[392], stage0_9[393], stage0_9[394], stage0_9[395]},
      {stage0_10[341]},
      {stage0_11[288], stage0_11[289], stage0_11[290], stage0_11[291], stage0_11[292], stage0_11[293]},
      {stage1_13[48],stage1_12[97],stage1_11[122],stage1_10[157],stage1_9[211]}
   );
   gpc615_5 gpc467 (
      {stage0_9[396], stage0_9[397], stage0_9[398], stage0_9[399], stage0_9[400]},
      {stage0_10[342]},
      {stage0_11[294], stage0_11[295], stage0_11[296], stage0_11[297], stage0_11[298], stage0_11[299]},
      {stage1_13[49],stage1_12[98],stage1_11[123],stage1_10[158],stage1_9[212]}
   );
   gpc615_5 gpc468 (
      {stage0_9[401], stage0_9[402], stage0_9[403], stage0_9[404], stage0_9[405]},
      {stage0_10[343]},
      {stage0_11[300], stage0_11[301], stage0_11[302], stage0_11[303], stage0_11[304], stage0_11[305]},
      {stage1_13[50],stage1_12[99],stage1_11[124],stage1_10[159],stage1_9[213]}
   );
   gpc615_5 gpc469 (
      {stage0_9[406], stage0_9[407], stage0_9[408], stage0_9[409], stage0_9[410]},
      {stage0_10[344]},
      {stage0_11[306], stage0_11[307], stage0_11[308], stage0_11[309], stage0_11[310], stage0_11[311]},
      {stage1_13[51],stage1_12[100],stage1_11[125],stage1_10[160],stage1_9[214]}
   );
   gpc615_5 gpc470 (
      {stage0_9[411], stage0_9[412], stage0_9[413], stage0_9[414], stage0_9[415]},
      {stage0_10[345]},
      {stage0_11[312], stage0_11[313], stage0_11[314], stage0_11[315], stage0_11[316], stage0_11[317]},
      {stage1_13[52],stage1_12[101],stage1_11[126],stage1_10[161],stage1_9[215]}
   );
   gpc615_5 gpc471 (
      {stage0_9[416], stage0_9[417], stage0_9[418], stage0_9[419], stage0_9[420]},
      {stage0_10[346]},
      {stage0_11[318], stage0_11[319], stage0_11[320], stage0_11[321], stage0_11[322], stage0_11[323]},
      {stage1_13[53],stage1_12[102],stage1_11[127],stage1_10[162],stage1_9[216]}
   );
   gpc615_5 gpc472 (
      {stage0_9[421], stage0_9[422], stage0_9[423], stage0_9[424], stage0_9[425]},
      {stage0_10[347]},
      {stage0_11[324], stage0_11[325], stage0_11[326], stage0_11[327], stage0_11[328], stage0_11[329]},
      {stage1_13[54],stage1_12[103],stage1_11[128],stage1_10[163],stage1_9[217]}
   );
   gpc615_5 gpc473 (
      {stage0_9[426], stage0_9[427], stage0_9[428], stage0_9[429], stage0_9[430]},
      {stage0_10[348]},
      {stage0_11[330], stage0_11[331], stage0_11[332], stage0_11[333], stage0_11[334], stage0_11[335]},
      {stage1_13[55],stage1_12[104],stage1_11[129],stage1_10[164],stage1_9[218]}
   );
   gpc615_5 gpc474 (
      {stage0_9[431], stage0_9[432], stage0_9[433], stage0_9[434], stage0_9[435]},
      {stage0_10[349]},
      {stage0_11[336], stage0_11[337], stage0_11[338], stage0_11[339], stage0_11[340], stage0_11[341]},
      {stage1_13[56],stage1_12[105],stage1_11[130],stage1_10[165],stage1_9[219]}
   );
   gpc615_5 gpc475 (
      {stage0_9[436], stage0_9[437], stage0_9[438], stage0_9[439], stage0_9[440]},
      {stage0_10[350]},
      {stage0_11[342], stage0_11[343], stage0_11[344], stage0_11[345], stage0_11[346], stage0_11[347]},
      {stage1_13[57],stage1_12[106],stage1_11[131],stage1_10[166],stage1_9[220]}
   );
   gpc615_5 gpc476 (
      {stage0_9[441], stage0_9[442], stage0_9[443], stage0_9[444], stage0_9[445]},
      {stage0_10[351]},
      {stage0_11[348], stage0_11[349], stage0_11[350], stage0_11[351], stage0_11[352], stage0_11[353]},
      {stage1_13[58],stage1_12[107],stage1_11[132],stage1_10[167],stage1_9[221]}
   );
   gpc615_5 gpc477 (
      {stage0_9[446], stage0_9[447], stage0_9[448], stage0_9[449], stage0_9[450]},
      {stage0_10[352]},
      {stage0_11[354], stage0_11[355], stage0_11[356], stage0_11[357], stage0_11[358], stage0_11[359]},
      {stage1_13[59],stage1_12[108],stage1_11[133],stage1_10[168],stage1_9[222]}
   );
   gpc615_5 gpc478 (
      {stage0_9[451], stage0_9[452], stage0_9[453], stage0_9[454], stage0_9[455]},
      {stage0_10[353]},
      {stage0_11[360], stage0_11[361], stage0_11[362], stage0_11[363], stage0_11[364], stage0_11[365]},
      {stage1_13[60],stage1_12[109],stage1_11[134],stage1_10[169],stage1_9[223]}
   );
   gpc615_5 gpc479 (
      {stage0_9[456], stage0_9[457], stage0_9[458], stage0_9[459], stage0_9[460]},
      {stage0_10[354]},
      {stage0_11[366], stage0_11[367], stage0_11[368], stage0_11[369], stage0_11[370], stage0_11[371]},
      {stage1_13[61],stage1_12[110],stage1_11[135],stage1_10[170],stage1_9[224]}
   );
   gpc615_5 gpc480 (
      {stage0_9[461], stage0_9[462], stage0_9[463], stage0_9[464], stage0_9[465]},
      {stage0_10[355]},
      {stage0_11[372], stage0_11[373], stage0_11[374], stage0_11[375], stage0_11[376], stage0_11[377]},
      {stage1_13[62],stage1_12[111],stage1_11[136],stage1_10[171],stage1_9[225]}
   );
   gpc615_5 gpc481 (
      {stage0_9[466], stage0_9[467], stage0_9[468], stage0_9[469], stage0_9[470]},
      {stage0_10[356]},
      {stage0_11[378], stage0_11[379], stage0_11[380], stage0_11[381], stage0_11[382], stage0_11[383]},
      {stage1_13[63],stage1_12[112],stage1_11[137],stage1_10[172],stage1_9[226]}
   );
   gpc615_5 gpc482 (
      {stage0_9[471], stage0_9[472], stage0_9[473], stage0_9[474], stage0_9[475]},
      {stage0_10[357]},
      {stage0_11[384], stage0_11[385], stage0_11[386], stage0_11[387], stage0_11[388], stage0_11[389]},
      {stage1_13[64],stage1_12[113],stage1_11[138],stage1_10[173],stage1_9[227]}
   );
   gpc606_5 gpc483 (
      {stage0_10[358], stage0_10[359], stage0_10[360], stage0_10[361], stage0_10[362], stage0_10[363]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[65],stage1_12[114],stage1_11[139],stage1_10[174]}
   );
   gpc606_5 gpc484 (
      {stage0_10[364], stage0_10[365], stage0_10[366], stage0_10[367], stage0_10[368], stage0_10[369]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[66],stage1_12[115],stage1_11[140],stage1_10[175]}
   );
   gpc606_5 gpc485 (
      {stage0_10[370], stage0_10[371], stage0_10[372], stage0_10[373], stage0_10[374], stage0_10[375]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[67],stage1_12[116],stage1_11[141],stage1_10[176]}
   );
   gpc606_5 gpc486 (
      {stage0_10[376], stage0_10[377], stage0_10[378], stage0_10[379], stage0_10[380], stage0_10[381]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[68],stage1_12[117],stage1_11[142],stage1_10[177]}
   );
   gpc606_5 gpc487 (
      {stage0_10[382], stage0_10[383], stage0_10[384], stage0_10[385], stage0_10[386], stage0_10[387]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[69],stage1_12[118],stage1_11[143],stage1_10[178]}
   );
   gpc606_5 gpc488 (
      {stage0_10[388], stage0_10[389], stage0_10[390], stage0_10[391], stage0_10[392], stage0_10[393]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[70],stage1_12[119],stage1_11[144],stage1_10[179]}
   );
   gpc615_5 gpc489 (
      {stage0_10[394], stage0_10[395], stage0_10[396], stage0_10[397], stage0_10[398]},
      {stage0_11[390]},
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage1_14[6],stage1_13[71],stage1_12[120],stage1_11[145],stage1_10[180]}
   );
   gpc615_5 gpc490 (
      {stage0_10[399], stage0_10[400], stage0_10[401], stage0_10[402], stage0_10[403]},
      {stage0_11[391]},
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage1_14[7],stage1_13[72],stage1_12[121],stage1_11[146],stage1_10[181]}
   );
   gpc615_5 gpc491 (
      {stage0_10[404], stage0_10[405], stage0_10[406], stage0_10[407], stage0_10[408]},
      {stage0_11[392]},
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage1_14[8],stage1_13[73],stage1_12[122],stage1_11[147],stage1_10[182]}
   );
   gpc615_5 gpc492 (
      {stage0_10[409], stage0_10[410], stage0_10[411], stage0_10[412], stage0_10[413]},
      {stage0_11[393]},
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage1_14[9],stage1_13[74],stage1_12[123],stage1_11[148],stage1_10[183]}
   );
   gpc615_5 gpc493 (
      {stage0_10[414], stage0_10[415], stage0_10[416], stage0_10[417], stage0_10[418]},
      {stage0_11[394]},
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage1_14[10],stage1_13[75],stage1_12[124],stage1_11[149],stage1_10[184]}
   );
   gpc615_5 gpc494 (
      {stage0_10[419], stage0_10[420], stage0_10[421], stage0_10[422], stage0_10[423]},
      {stage0_11[395]},
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage1_14[11],stage1_13[76],stage1_12[125],stage1_11[150],stage1_10[185]}
   );
   gpc615_5 gpc495 (
      {stage0_10[424], stage0_10[425], stage0_10[426], stage0_10[427], stage0_10[428]},
      {stage0_11[396]},
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage1_14[12],stage1_13[77],stage1_12[126],stage1_11[151],stage1_10[186]}
   );
   gpc615_5 gpc496 (
      {stage0_10[429], stage0_10[430], stage0_10[431], stage0_10[432], stage0_10[433]},
      {stage0_11[397]},
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage1_14[13],stage1_13[78],stage1_12[127],stage1_11[152],stage1_10[187]}
   );
   gpc615_5 gpc497 (
      {stage0_10[434], stage0_10[435], stage0_10[436], stage0_10[437], stage0_10[438]},
      {stage0_11[398]},
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage1_14[14],stage1_13[79],stage1_12[128],stage1_11[153],stage1_10[188]}
   );
   gpc615_5 gpc498 (
      {stage0_10[439], stage0_10[440], stage0_10[441], stage0_10[442], stage0_10[443]},
      {stage0_11[399]},
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage1_14[15],stage1_13[80],stage1_12[129],stage1_11[154],stage1_10[189]}
   );
   gpc615_5 gpc499 (
      {stage0_10[444], stage0_10[445], stage0_10[446], stage0_10[447], stage0_10[448]},
      {stage0_11[400]},
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage1_14[16],stage1_13[81],stage1_12[130],stage1_11[155],stage1_10[190]}
   );
   gpc615_5 gpc500 (
      {stage0_10[449], stage0_10[450], stage0_10[451], stage0_10[452], stage0_10[453]},
      {stage0_11[401]},
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage1_14[17],stage1_13[82],stage1_12[131],stage1_11[156],stage1_10[191]}
   );
   gpc615_5 gpc501 (
      {stage0_10[454], stage0_10[455], stage0_10[456], stage0_10[457], stage0_10[458]},
      {stage0_11[402]},
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage1_14[18],stage1_13[83],stage1_12[132],stage1_11[157],stage1_10[192]}
   );
   gpc615_5 gpc502 (
      {stage0_10[459], stage0_10[460], stage0_10[461], stage0_10[462], stage0_10[463]},
      {stage0_11[403]},
      {stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage1_14[19],stage1_13[84],stage1_12[133],stage1_11[158],stage1_10[193]}
   );
   gpc615_5 gpc503 (
      {stage0_10[464], stage0_10[465], stage0_10[466], stage0_10[467], stage0_10[468]},
      {stage0_11[404]},
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125]},
      {stage1_14[20],stage1_13[85],stage1_12[134],stage1_11[159],stage1_10[194]}
   );
   gpc615_5 gpc504 (
      {stage0_10[469], stage0_10[470], stage0_10[471], stage0_10[472], stage0_10[473]},
      {stage0_11[405]},
      {stage0_12[126], stage0_12[127], stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131]},
      {stage1_14[21],stage1_13[86],stage1_12[135],stage1_11[160],stage1_10[195]}
   );
   gpc615_5 gpc505 (
      {stage0_10[474], stage0_10[475], stage0_10[476], stage0_10[477], stage0_10[478]},
      {stage0_11[406]},
      {stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137]},
      {stage1_14[22],stage1_13[87],stage1_12[136],stage1_11[161],stage1_10[196]}
   );
   gpc615_5 gpc506 (
      {stage0_10[479], stage0_10[480], stage0_10[481], stage0_10[482], stage0_10[483]},
      {stage0_11[407]},
      {stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141], stage0_12[142], stage0_12[143]},
      {stage1_14[23],stage1_13[88],stage1_12[137],stage1_11[162],stage1_10[197]}
   );
   gpc615_5 gpc507 (
      {stage0_10[484], stage0_10[485], stage0_10[486], stage0_10[487], stage0_10[488]},
      {stage0_11[408]},
      {stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147], stage0_12[148], stage0_12[149]},
      {stage1_14[24],stage1_13[89],stage1_12[138],stage1_11[163],stage1_10[198]}
   );
   gpc615_5 gpc508 (
      {stage0_10[489], stage0_10[490], stage0_10[491], stage0_10[492], stage0_10[493]},
      {stage0_11[409]},
      {stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155]},
      {stage1_14[25],stage1_13[90],stage1_12[139],stage1_11[164],stage1_10[199]}
   );
   gpc615_5 gpc509 (
      {stage0_10[494], stage0_10[495], stage0_10[496], stage0_10[497], stage0_10[498]},
      {stage0_11[410]},
      {stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage1_14[26],stage1_13[91],stage1_12[140],stage1_11[165],stage1_10[200]}
   );
   gpc615_5 gpc510 (
      {stage0_10[499], stage0_10[500], stage0_10[501], stage0_10[502], stage0_10[503]},
      {stage0_11[411]},
      {stage0_12[162], stage0_12[163], stage0_12[164], stage0_12[165], stage0_12[166], stage0_12[167]},
      {stage1_14[27],stage1_13[92],stage1_12[141],stage1_11[166],stage1_10[201]}
   );
   gpc606_5 gpc511 (
      {stage0_11[412], stage0_11[413], stage0_11[414], stage0_11[415], stage0_11[416], stage0_11[417]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[28],stage1_13[93],stage1_12[142],stage1_11[167]}
   );
   gpc606_5 gpc512 (
      {stage0_11[418], stage0_11[419], stage0_11[420], stage0_11[421], stage0_11[422], stage0_11[423]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[29],stage1_13[94],stage1_12[143],stage1_11[168]}
   );
   gpc606_5 gpc513 (
      {stage0_11[424], stage0_11[425], stage0_11[426], stage0_11[427], stage0_11[428], stage0_11[429]},
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage1_15[2],stage1_14[30],stage1_13[95],stage1_12[144],stage1_11[169]}
   );
   gpc606_5 gpc514 (
      {stage0_11[430], stage0_11[431], stage0_11[432], stage0_11[433], stage0_11[434], stage0_11[435]},
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage1_15[3],stage1_14[31],stage1_13[96],stage1_12[145],stage1_11[170]}
   );
   gpc606_5 gpc515 (
      {stage0_11[436], stage0_11[437], stage0_11[438], stage0_11[439], stage0_11[440], stage0_11[441]},
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage1_15[4],stage1_14[32],stage1_13[97],stage1_12[146],stage1_11[171]}
   );
   gpc606_5 gpc516 (
      {stage0_11[442], stage0_11[443], stage0_11[444], stage0_11[445], stage0_11[446], stage0_11[447]},
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage1_15[5],stage1_14[33],stage1_13[98],stage1_12[147],stage1_11[172]}
   );
   gpc606_5 gpc517 (
      {stage0_11[448], stage0_11[449], stage0_11[450], stage0_11[451], stage0_11[452], stage0_11[453]},
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage1_15[6],stage1_14[34],stage1_13[99],stage1_12[148],stage1_11[173]}
   );
   gpc606_5 gpc518 (
      {stage0_11[454], stage0_11[455], stage0_11[456], stage0_11[457], stage0_11[458], stage0_11[459]},
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage1_15[7],stage1_14[35],stage1_13[100],stage1_12[149],stage1_11[174]}
   );
   gpc606_5 gpc519 (
      {stage0_11[460], stage0_11[461], stage0_11[462], stage0_11[463], stage0_11[464], stage0_11[465]},
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage1_15[8],stage1_14[36],stage1_13[101],stage1_12[150],stage1_11[175]}
   );
   gpc615_5 gpc520 (
      {stage0_11[466], stage0_11[467], stage0_11[468], stage0_11[469], stage0_11[470]},
      {stage0_12[168]},
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage1_15[9],stage1_14[37],stage1_13[102],stage1_12[151],stage1_11[176]}
   );
   gpc615_5 gpc521 (
      {stage0_11[471], stage0_11[472], stage0_11[473], stage0_11[474], stage0_11[475]},
      {stage0_12[169]},
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage1_15[10],stage1_14[38],stage1_13[103],stage1_12[152],stage1_11[177]}
   );
   gpc615_5 gpc522 (
      {stage0_11[476], stage0_11[477], stage0_11[478], stage0_11[479], stage0_11[480]},
      {stage0_12[170]},
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage1_15[11],stage1_14[39],stage1_13[104],stage1_12[153],stage1_11[178]}
   );
   gpc615_5 gpc523 (
      {stage0_11[481], stage0_11[482], stage0_11[483], stage0_11[484], stage0_11[485]},
      {stage0_12[171]},
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage1_15[12],stage1_14[40],stage1_13[105],stage1_12[154],stage1_11[179]}
   );
   gpc615_5 gpc524 (
      {stage0_11[486], stage0_11[487], stage0_11[488], stage0_11[489], stage0_11[490]},
      {stage0_12[172]},
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage1_15[13],stage1_14[41],stage1_13[106],stage1_12[155],stage1_11[180]}
   );
   gpc615_5 gpc525 (
      {stage0_11[491], stage0_11[492], stage0_11[493], stage0_11[494], stage0_11[495]},
      {stage0_12[173]},
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage1_15[14],stage1_14[42],stage1_13[107],stage1_12[156],stage1_11[181]}
   );
   gpc615_5 gpc526 (
      {stage0_11[496], stage0_11[497], stage0_11[498], stage0_11[499], stage0_11[500]},
      {stage0_12[174]},
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage1_15[15],stage1_14[43],stage1_13[108],stage1_12[157],stage1_11[182]}
   );
   gpc615_5 gpc527 (
      {stage0_11[501], stage0_11[502], stage0_11[503], stage0_11[504], stage0_11[505]},
      {stage0_12[175]},
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage1_15[16],stage1_14[44],stage1_13[109],stage1_12[158],stage1_11[183]}
   );
   gpc606_5 gpc528 (
      {stage0_12[176], stage0_12[177], stage0_12[178], stage0_12[179], stage0_12[180], stage0_12[181]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[17],stage1_14[45],stage1_13[110],stage1_12[159]}
   );
   gpc606_5 gpc529 (
      {stage0_12[182], stage0_12[183], stage0_12[184], stage0_12[185], stage0_12[186], stage0_12[187]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[18],stage1_14[46],stage1_13[111],stage1_12[160]}
   );
   gpc606_5 gpc530 (
      {stage0_12[188], stage0_12[189], stage0_12[190], stage0_12[191], stage0_12[192], stage0_12[193]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[19],stage1_14[47],stage1_13[112],stage1_12[161]}
   );
   gpc606_5 gpc531 (
      {stage0_12[194], stage0_12[195], stage0_12[196], stage0_12[197], stage0_12[198], stage0_12[199]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[20],stage1_14[48],stage1_13[113],stage1_12[162]}
   );
   gpc606_5 gpc532 (
      {stage0_12[200], stage0_12[201], stage0_12[202], stage0_12[203], stage0_12[204], stage0_12[205]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[21],stage1_14[49],stage1_13[114],stage1_12[163]}
   );
   gpc606_5 gpc533 (
      {stage0_12[206], stage0_12[207], stage0_12[208], stage0_12[209], stage0_12[210], stage0_12[211]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[22],stage1_14[50],stage1_13[115],stage1_12[164]}
   );
   gpc606_5 gpc534 (
      {stage0_12[212], stage0_12[213], stage0_12[214], stage0_12[215], stage0_12[216], stage0_12[217]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[23],stage1_14[51],stage1_13[116],stage1_12[165]}
   );
   gpc606_5 gpc535 (
      {stage0_12[218], stage0_12[219], stage0_12[220], stage0_12[221], stage0_12[222], stage0_12[223]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[24],stage1_14[52],stage1_13[117],stage1_12[166]}
   );
   gpc606_5 gpc536 (
      {stage0_12[224], stage0_12[225], stage0_12[226], stage0_12[227], stage0_12[228], stage0_12[229]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[25],stage1_14[53],stage1_13[118],stage1_12[167]}
   );
   gpc606_5 gpc537 (
      {stage0_12[230], stage0_12[231], stage0_12[232], stage0_12[233], stage0_12[234], stage0_12[235]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[26],stage1_14[54],stage1_13[119],stage1_12[168]}
   );
   gpc606_5 gpc538 (
      {stage0_12[236], stage0_12[237], stage0_12[238], stage0_12[239], stage0_12[240], stage0_12[241]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[27],stage1_14[55],stage1_13[120],stage1_12[169]}
   );
   gpc606_5 gpc539 (
      {stage0_12[242], stage0_12[243], stage0_12[244], stage0_12[245], stage0_12[246], stage0_12[247]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[28],stage1_14[56],stage1_13[121],stage1_12[170]}
   );
   gpc606_5 gpc540 (
      {stage0_12[248], stage0_12[249], stage0_12[250], stage0_12[251], stage0_12[252], stage0_12[253]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[29],stage1_14[57],stage1_13[122],stage1_12[171]}
   );
   gpc606_5 gpc541 (
      {stage0_12[254], stage0_12[255], stage0_12[256], stage0_12[257], stage0_12[258], stage0_12[259]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[30],stage1_14[58],stage1_13[123],stage1_12[172]}
   );
   gpc606_5 gpc542 (
      {stage0_12[260], stage0_12[261], stage0_12[262], stage0_12[263], stage0_12[264], stage0_12[265]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[31],stage1_14[59],stage1_13[124],stage1_12[173]}
   );
   gpc606_5 gpc543 (
      {stage0_12[266], stage0_12[267], stage0_12[268], stage0_12[269], stage0_12[270], stage0_12[271]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[32],stage1_14[60],stage1_13[125],stage1_12[174]}
   );
   gpc606_5 gpc544 (
      {stage0_12[272], stage0_12[273], stage0_12[274], stage0_12[275], stage0_12[276], stage0_12[277]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[33],stage1_14[61],stage1_13[126],stage1_12[175]}
   );
   gpc606_5 gpc545 (
      {stage0_12[278], stage0_12[279], stage0_12[280], stage0_12[281], stage0_12[282], stage0_12[283]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[34],stage1_14[62],stage1_13[127],stage1_12[176]}
   );
   gpc606_5 gpc546 (
      {stage0_12[284], stage0_12[285], stage0_12[286], stage0_12[287], stage0_12[288], stage0_12[289]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[35],stage1_14[63],stage1_13[128],stage1_12[177]}
   );
   gpc606_5 gpc547 (
      {stage0_12[290], stage0_12[291], stage0_12[292], stage0_12[293], stage0_12[294], stage0_12[295]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[36],stage1_14[64],stage1_13[129],stage1_12[178]}
   );
   gpc606_5 gpc548 (
      {stage0_12[296], stage0_12[297], stage0_12[298], stage0_12[299], stage0_12[300], stage0_12[301]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[37],stage1_14[65],stage1_13[130],stage1_12[179]}
   );
   gpc615_5 gpc549 (
      {stage0_12[302], stage0_12[303], stage0_12[304], stage0_12[305], stage0_12[306]},
      {stage0_13[102]},
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131]},
      {stage1_16[21],stage1_15[38],stage1_14[66],stage1_13[131],stage1_12[180]}
   );
   gpc615_5 gpc550 (
      {stage0_12[307], stage0_12[308], stage0_12[309], stage0_12[310], stage0_12[311]},
      {stage0_13[103]},
      {stage0_14[132], stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137]},
      {stage1_16[22],stage1_15[39],stage1_14[67],stage1_13[132],stage1_12[181]}
   );
   gpc615_5 gpc551 (
      {stage0_12[312], stage0_12[313], stage0_12[314], stage0_12[315], stage0_12[316]},
      {stage0_13[104]},
      {stage0_14[138], stage0_14[139], stage0_14[140], stage0_14[141], stage0_14[142], stage0_14[143]},
      {stage1_16[23],stage1_15[40],stage1_14[68],stage1_13[133],stage1_12[182]}
   );
   gpc615_5 gpc552 (
      {stage0_12[317], stage0_12[318], stage0_12[319], stage0_12[320], stage0_12[321]},
      {stage0_13[105]},
      {stage0_14[144], stage0_14[145], stage0_14[146], stage0_14[147], stage0_14[148], stage0_14[149]},
      {stage1_16[24],stage1_15[41],stage1_14[69],stage1_13[134],stage1_12[183]}
   );
   gpc615_5 gpc553 (
      {stage0_12[322], stage0_12[323], stage0_12[324], stage0_12[325], stage0_12[326]},
      {stage0_13[106]},
      {stage0_14[150], stage0_14[151], stage0_14[152], stage0_14[153], stage0_14[154], stage0_14[155]},
      {stage1_16[25],stage1_15[42],stage1_14[70],stage1_13[135],stage1_12[184]}
   );
   gpc615_5 gpc554 (
      {stage0_12[327], stage0_12[328], stage0_12[329], stage0_12[330], stage0_12[331]},
      {stage0_13[107]},
      {stage0_14[156], stage0_14[157], stage0_14[158], stage0_14[159], stage0_14[160], stage0_14[161]},
      {stage1_16[26],stage1_15[43],stage1_14[71],stage1_13[136],stage1_12[185]}
   );
   gpc615_5 gpc555 (
      {stage0_12[332], stage0_12[333], stage0_12[334], stage0_12[335], stage0_12[336]},
      {stage0_13[108]},
      {stage0_14[162], stage0_14[163], stage0_14[164], stage0_14[165], stage0_14[166], stage0_14[167]},
      {stage1_16[27],stage1_15[44],stage1_14[72],stage1_13[137],stage1_12[186]}
   );
   gpc615_5 gpc556 (
      {stage0_12[337], stage0_12[338], stage0_12[339], stage0_12[340], stage0_12[341]},
      {stage0_13[109]},
      {stage0_14[168], stage0_14[169], stage0_14[170], stage0_14[171], stage0_14[172], stage0_14[173]},
      {stage1_16[28],stage1_15[45],stage1_14[73],stage1_13[138],stage1_12[187]}
   );
   gpc615_5 gpc557 (
      {stage0_12[342], stage0_12[343], stage0_12[344], stage0_12[345], stage0_12[346]},
      {stage0_13[110]},
      {stage0_14[174], stage0_14[175], stage0_14[176], stage0_14[177], stage0_14[178], stage0_14[179]},
      {stage1_16[29],stage1_15[46],stage1_14[74],stage1_13[139],stage1_12[188]}
   );
   gpc615_5 gpc558 (
      {stage0_12[347], stage0_12[348], stage0_12[349], stage0_12[350], stage0_12[351]},
      {stage0_13[111]},
      {stage0_14[180], stage0_14[181], stage0_14[182], stage0_14[183], stage0_14[184], stage0_14[185]},
      {stage1_16[30],stage1_15[47],stage1_14[75],stage1_13[140],stage1_12[189]}
   );
   gpc615_5 gpc559 (
      {stage0_12[352], stage0_12[353], stage0_12[354], stage0_12[355], stage0_12[356]},
      {stage0_13[112]},
      {stage0_14[186], stage0_14[187], stage0_14[188], stage0_14[189], stage0_14[190], stage0_14[191]},
      {stage1_16[31],stage1_15[48],stage1_14[76],stage1_13[141],stage1_12[190]}
   );
   gpc615_5 gpc560 (
      {stage0_12[357], stage0_12[358], stage0_12[359], stage0_12[360], stage0_12[361]},
      {stage0_13[113]},
      {stage0_14[192], stage0_14[193], stage0_14[194], stage0_14[195], stage0_14[196], stage0_14[197]},
      {stage1_16[32],stage1_15[49],stage1_14[77],stage1_13[142],stage1_12[191]}
   );
   gpc615_5 gpc561 (
      {stage0_12[362], stage0_12[363], stage0_12[364], stage0_12[365], stage0_12[366]},
      {stage0_13[114]},
      {stage0_14[198], stage0_14[199], stage0_14[200], stage0_14[201], stage0_14[202], stage0_14[203]},
      {stage1_16[33],stage1_15[50],stage1_14[78],stage1_13[143],stage1_12[192]}
   );
   gpc615_5 gpc562 (
      {stage0_12[367], stage0_12[368], stage0_12[369], stage0_12[370], stage0_12[371]},
      {stage0_13[115]},
      {stage0_14[204], stage0_14[205], stage0_14[206], stage0_14[207], stage0_14[208], stage0_14[209]},
      {stage1_16[34],stage1_15[51],stage1_14[79],stage1_13[144],stage1_12[193]}
   );
   gpc615_5 gpc563 (
      {stage0_12[372], stage0_12[373], stage0_12[374], stage0_12[375], stage0_12[376]},
      {stage0_13[116]},
      {stage0_14[210], stage0_14[211], stage0_14[212], stage0_14[213], stage0_14[214], stage0_14[215]},
      {stage1_16[35],stage1_15[52],stage1_14[80],stage1_13[145],stage1_12[194]}
   );
   gpc615_5 gpc564 (
      {stage0_12[377], stage0_12[378], stage0_12[379], stage0_12[380], stage0_12[381]},
      {stage0_13[117]},
      {stage0_14[216], stage0_14[217], stage0_14[218], stage0_14[219], stage0_14[220], stage0_14[221]},
      {stage1_16[36],stage1_15[53],stage1_14[81],stage1_13[146],stage1_12[195]}
   );
   gpc615_5 gpc565 (
      {stage0_12[382], stage0_12[383], stage0_12[384], stage0_12[385], stage0_12[386]},
      {stage0_13[118]},
      {stage0_14[222], stage0_14[223], stage0_14[224], stage0_14[225], stage0_14[226], stage0_14[227]},
      {stage1_16[37],stage1_15[54],stage1_14[82],stage1_13[147],stage1_12[196]}
   );
   gpc615_5 gpc566 (
      {stage0_12[387], stage0_12[388], stage0_12[389], stage0_12[390], stage0_12[391]},
      {stage0_13[119]},
      {stage0_14[228], stage0_14[229], stage0_14[230], stage0_14[231], stage0_14[232], stage0_14[233]},
      {stage1_16[38],stage1_15[55],stage1_14[83],stage1_13[148],stage1_12[197]}
   );
   gpc615_5 gpc567 (
      {stage0_12[392], stage0_12[393], stage0_12[394], stage0_12[395], stage0_12[396]},
      {stage0_13[120]},
      {stage0_14[234], stage0_14[235], stage0_14[236], stage0_14[237], stage0_14[238], stage0_14[239]},
      {stage1_16[39],stage1_15[56],stage1_14[84],stage1_13[149],stage1_12[198]}
   );
   gpc615_5 gpc568 (
      {stage0_12[397], stage0_12[398], stage0_12[399], stage0_12[400], stage0_12[401]},
      {stage0_13[121]},
      {stage0_14[240], stage0_14[241], stage0_14[242], stage0_14[243], stage0_14[244], stage0_14[245]},
      {stage1_16[40],stage1_15[57],stage1_14[85],stage1_13[150],stage1_12[199]}
   );
   gpc615_5 gpc569 (
      {stage0_12[402], stage0_12[403], stage0_12[404], stage0_12[405], stage0_12[406]},
      {stage0_13[122]},
      {stage0_14[246], stage0_14[247], stage0_14[248], stage0_14[249], stage0_14[250], stage0_14[251]},
      {stage1_16[41],stage1_15[58],stage1_14[86],stage1_13[151],stage1_12[200]}
   );
   gpc615_5 gpc570 (
      {stage0_12[407], stage0_12[408], stage0_12[409], stage0_12[410], stage0_12[411]},
      {stage0_13[123]},
      {stage0_14[252], stage0_14[253], stage0_14[254], stage0_14[255], stage0_14[256], stage0_14[257]},
      {stage1_16[42],stage1_15[59],stage1_14[87],stage1_13[152],stage1_12[201]}
   );
   gpc615_5 gpc571 (
      {stage0_12[412], stage0_12[413], stage0_12[414], stage0_12[415], stage0_12[416]},
      {stage0_13[124]},
      {stage0_14[258], stage0_14[259], stage0_14[260], stage0_14[261], stage0_14[262], stage0_14[263]},
      {stage1_16[43],stage1_15[60],stage1_14[88],stage1_13[153],stage1_12[202]}
   );
   gpc615_5 gpc572 (
      {stage0_12[417], stage0_12[418], stage0_12[419], stage0_12[420], stage0_12[421]},
      {stage0_13[125]},
      {stage0_14[264], stage0_14[265], stage0_14[266], stage0_14[267], stage0_14[268], stage0_14[269]},
      {stage1_16[44],stage1_15[61],stage1_14[89],stage1_13[154],stage1_12[203]}
   );
   gpc615_5 gpc573 (
      {stage0_12[422], stage0_12[423], stage0_12[424], stage0_12[425], stage0_12[426]},
      {stage0_13[126]},
      {stage0_14[270], stage0_14[271], stage0_14[272], stage0_14[273], stage0_14[274], stage0_14[275]},
      {stage1_16[45],stage1_15[62],stage1_14[90],stage1_13[155],stage1_12[204]}
   );
   gpc615_5 gpc574 (
      {stage0_12[427], stage0_12[428], stage0_12[429], stage0_12[430], stage0_12[431]},
      {stage0_13[127]},
      {stage0_14[276], stage0_14[277], stage0_14[278], stage0_14[279], stage0_14[280], stage0_14[281]},
      {stage1_16[46],stage1_15[63],stage1_14[91],stage1_13[156],stage1_12[205]}
   );
   gpc615_5 gpc575 (
      {stage0_12[432], stage0_12[433], stage0_12[434], stage0_12[435], stage0_12[436]},
      {stage0_13[128]},
      {stage0_14[282], stage0_14[283], stage0_14[284], stage0_14[285], stage0_14[286], stage0_14[287]},
      {stage1_16[47],stage1_15[64],stage1_14[92],stage1_13[157],stage1_12[206]}
   );
   gpc615_5 gpc576 (
      {stage0_12[437], stage0_12[438], stage0_12[439], stage0_12[440], stage0_12[441]},
      {stage0_13[129]},
      {stage0_14[288], stage0_14[289], stage0_14[290], stage0_14[291], stage0_14[292], stage0_14[293]},
      {stage1_16[48],stage1_15[65],stage1_14[93],stage1_13[158],stage1_12[207]}
   );
   gpc615_5 gpc577 (
      {stage0_12[442], stage0_12[443], stage0_12[444], stage0_12[445], stage0_12[446]},
      {stage0_13[130]},
      {stage0_14[294], stage0_14[295], stage0_14[296], stage0_14[297], stage0_14[298], stage0_14[299]},
      {stage1_16[49],stage1_15[66],stage1_14[94],stage1_13[159],stage1_12[208]}
   );
   gpc615_5 gpc578 (
      {stage0_12[447], stage0_12[448], stage0_12[449], stage0_12[450], stage0_12[451]},
      {stage0_13[131]},
      {stage0_14[300], stage0_14[301], stage0_14[302], stage0_14[303], stage0_14[304], stage0_14[305]},
      {stage1_16[50],stage1_15[67],stage1_14[95],stage1_13[160],stage1_12[209]}
   );
   gpc615_5 gpc579 (
      {stage0_12[452], stage0_12[453], stage0_12[454], stage0_12[455], stage0_12[456]},
      {stage0_13[132]},
      {stage0_14[306], stage0_14[307], stage0_14[308], stage0_14[309], stage0_14[310], stage0_14[311]},
      {stage1_16[51],stage1_15[68],stage1_14[96],stage1_13[161],stage1_12[210]}
   );
   gpc615_5 gpc580 (
      {stage0_12[457], stage0_12[458], stage0_12[459], stage0_12[460], stage0_12[461]},
      {stage0_13[133]},
      {stage0_14[312], stage0_14[313], stage0_14[314], stage0_14[315], stage0_14[316], stage0_14[317]},
      {stage1_16[52],stage1_15[69],stage1_14[97],stage1_13[162],stage1_12[211]}
   );
   gpc615_5 gpc581 (
      {stage0_12[462], stage0_12[463], stage0_12[464], stage0_12[465], stage0_12[466]},
      {stage0_13[134]},
      {stage0_14[318], stage0_14[319], stage0_14[320], stage0_14[321], stage0_14[322], stage0_14[323]},
      {stage1_16[53],stage1_15[70],stage1_14[98],stage1_13[163],stage1_12[212]}
   );
   gpc615_5 gpc582 (
      {stage0_12[467], stage0_12[468], stage0_12[469], stage0_12[470], stage0_12[471]},
      {stage0_13[135]},
      {stage0_14[324], stage0_14[325], stage0_14[326], stage0_14[327], stage0_14[328], stage0_14[329]},
      {stage1_16[54],stage1_15[71],stage1_14[99],stage1_13[164],stage1_12[213]}
   );
   gpc615_5 gpc583 (
      {stage0_12[472], stage0_12[473], stage0_12[474], stage0_12[475], stage0_12[476]},
      {stage0_13[136]},
      {stage0_14[330], stage0_14[331], stage0_14[332], stage0_14[333], stage0_14[334], stage0_14[335]},
      {stage1_16[55],stage1_15[72],stage1_14[100],stage1_13[165],stage1_12[214]}
   );
   gpc615_5 gpc584 (
      {stage0_12[477], stage0_12[478], stage0_12[479], stage0_12[480], stage0_12[481]},
      {stage0_13[137]},
      {stage0_14[336], stage0_14[337], stage0_14[338], stage0_14[339], stage0_14[340], stage0_14[341]},
      {stage1_16[56],stage1_15[73],stage1_14[101],stage1_13[166],stage1_12[215]}
   );
   gpc615_5 gpc585 (
      {stage0_12[482], stage0_12[483], stage0_12[484], stage0_12[485], stage0_12[486]},
      {stage0_13[138]},
      {stage0_14[342], stage0_14[343], stage0_14[344], stage0_14[345], stage0_14[346], stage0_14[347]},
      {stage1_16[57],stage1_15[74],stage1_14[102],stage1_13[167],stage1_12[216]}
   );
   gpc615_5 gpc586 (
      {stage0_12[487], stage0_12[488], stage0_12[489], stage0_12[490], stage0_12[491]},
      {stage0_13[139]},
      {stage0_14[348], stage0_14[349], stage0_14[350], stage0_14[351], stage0_14[352], stage0_14[353]},
      {stage1_16[58],stage1_15[75],stage1_14[103],stage1_13[168],stage1_12[217]}
   );
   gpc615_5 gpc587 (
      {stage0_12[492], stage0_12[493], stage0_12[494], stage0_12[495], stage0_12[496]},
      {stage0_13[140]},
      {stage0_14[354], stage0_14[355], stage0_14[356], stage0_14[357], stage0_14[358], stage0_14[359]},
      {stage1_16[59],stage1_15[76],stage1_14[104],stage1_13[169],stage1_12[218]}
   );
   gpc615_5 gpc588 (
      {stage0_12[497], stage0_12[498], stage0_12[499], stage0_12[500], stage0_12[501]},
      {stage0_13[141]},
      {stage0_14[360], stage0_14[361], stage0_14[362], stage0_14[363], stage0_14[364], stage0_14[365]},
      {stage1_16[60],stage1_15[77],stage1_14[105],stage1_13[170],stage1_12[219]}
   );
   gpc615_5 gpc589 (
      {stage0_12[502], stage0_12[503], stage0_12[504], stage0_12[505], stage0_12[506]},
      {stage0_13[142]},
      {stage0_14[366], stage0_14[367], stage0_14[368], stage0_14[369], stage0_14[370], stage0_14[371]},
      {stage1_16[61],stage1_15[78],stage1_14[106],stage1_13[171],stage1_12[220]}
   );
   gpc615_5 gpc590 (
      {stage0_12[507], stage0_12[508], stage0_12[509], stage0_12[510], stage0_12[511]},
      {stage0_13[143]},
      {stage0_14[372], stage0_14[373], stage0_14[374], stage0_14[375], stage0_14[376], stage0_14[377]},
      {stage1_16[62],stage1_15[79],stage1_14[107],stage1_13[172],stage1_12[221]}
   );
   gpc606_5 gpc591 (
      {stage0_13[144], stage0_13[145], stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[63],stage1_15[80],stage1_14[108],stage1_13[173]}
   );
   gpc606_5 gpc592 (
      {stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154], stage0_13[155]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[64],stage1_15[81],stage1_14[109],stage1_13[174]}
   );
   gpc606_5 gpc593 (
      {stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159], stage0_13[160], stage0_13[161]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[65],stage1_15[82],stage1_14[110],stage1_13[175]}
   );
   gpc615_5 gpc594 (
      {stage0_13[162], stage0_13[163], stage0_13[164], stage0_13[165], stage0_13[166]},
      {stage0_14[378]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[66],stage1_15[83],stage1_14[111],stage1_13[176]}
   );
   gpc615_5 gpc595 (
      {stage0_13[167], stage0_13[168], stage0_13[169], stage0_13[170], stage0_13[171]},
      {stage0_14[379]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[67],stage1_15[84],stage1_14[112],stage1_13[177]}
   );
   gpc615_5 gpc596 (
      {stage0_13[172], stage0_13[173], stage0_13[174], stage0_13[175], stage0_13[176]},
      {stage0_14[380]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[68],stage1_15[85],stage1_14[113],stage1_13[178]}
   );
   gpc615_5 gpc597 (
      {stage0_13[177], stage0_13[178], stage0_13[179], stage0_13[180], stage0_13[181]},
      {stage0_14[381]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[69],stage1_15[86],stage1_14[114],stage1_13[179]}
   );
   gpc615_5 gpc598 (
      {stage0_13[182], stage0_13[183], stage0_13[184], stage0_13[185], stage0_13[186]},
      {stage0_14[382]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[70],stage1_15[87],stage1_14[115],stage1_13[180]}
   );
   gpc615_5 gpc599 (
      {stage0_13[187], stage0_13[188], stage0_13[189], stage0_13[190], stage0_13[191]},
      {stage0_14[383]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[71],stage1_15[88],stage1_14[116],stage1_13[181]}
   );
   gpc615_5 gpc600 (
      {stage0_13[192], stage0_13[193], stage0_13[194], stage0_13[195], stage0_13[196]},
      {stage0_14[384]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[72],stage1_15[89],stage1_14[117],stage1_13[182]}
   );
   gpc615_5 gpc601 (
      {stage0_13[197], stage0_13[198], stage0_13[199], stage0_13[200], stage0_13[201]},
      {stage0_14[385]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[73],stage1_15[90],stage1_14[118],stage1_13[183]}
   );
   gpc615_5 gpc602 (
      {stage0_13[202], stage0_13[203], stage0_13[204], stage0_13[205], stage0_13[206]},
      {stage0_14[386]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[74],stage1_15[91],stage1_14[119],stage1_13[184]}
   );
   gpc615_5 gpc603 (
      {stage0_13[207], stage0_13[208], stage0_13[209], stage0_13[210], stage0_13[211]},
      {stage0_14[387]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[75],stage1_15[92],stage1_14[120],stage1_13[185]}
   );
   gpc615_5 gpc604 (
      {stage0_13[212], stage0_13[213], stage0_13[214], stage0_13[215], stage0_13[216]},
      {stage0_14[388]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[76],stage1_15[93],stage1_14[121],stage1_13[186]}
   );
   gpc615_5 gpc605 (
      {stage0_13[217], stage0_13[218], stage0_13[219], stage0_13[220], stage0_13[221]},
      {stage0_14[389]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[77],stage1_15[94],stage1_14[122],stage1_13[187]}
   );
   gpc615_5 gpc606 (
      {stage0_13[222], stage0_13[223], stage0_13[224], stage0_13[225], stage0_13[226]},
      {stage0_14[390]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[78],stage1_15[95],stage1_14[123],stage1_13[188]}
   );
   gpc615_5 gpc607 (
      {stage0_13[227], stage0_13[228], stage0_13[229], stage0_13[230], stage0_13[231]},
      {stage0_14[391]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[79],stage1_15[96],stage1_14[124],stage1_13[189]}
   );
   gpc615_5 gpc608 (
      {stage0_13[232], stage0_13[233], stage0_13[234], stage0_13[235], stage0_13[236]},
      {stage0_14[392]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[80],stage1_15[97],stage1_14[125],stage1_13[190]}
   );
   gpc615_5 gpc609 (
      {stage0_13[237], stage0_13[238], stage0_13[239], stage0_13[240], stage0_13[241]},
      {stage0_14[393]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[81],stage1_15[98],stage1_14[126],stage1_13[191]}
   );
   gpc615_5 gpc610 (
      {stage0_13[242], stage0_13[243], stage0_13[244], stage0_13[245], stage0_13[246]},
      {stage0_14[394]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[82],stage1_15[99],stage1_14[127],stage1_13[192]}
   );
   gpc615_5 gpc611 (
      {stage0_13[247], stage0_13[248], stage0_13[249], stage0_13[250], stage0_13[251]},
      {stage0_14[395]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[83],stage1_15[100],stage1_14[128],stage1_13[193]}
   );
   gpc615_5 gpc612 (
      {stage0_13[252], stage0_13[253], stage0_13[254], stage0_13[255], stage0_13[256]},
      {stage0_14[396]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[84],stage1_15[101],stage1_14[129],stage1_13[194]}
   );
   gpc615_5 gpc613 (
      {stage0_13[257], stage0_13[258], stage0_13[259], stage0_13[260], stage0_13[261]},
      {stage0_14[397]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[85],stage1_15[102],stage1_14[130],stage1_13[195]}
   );
   gpc615_5 gpc614 (
      {stage0_13[262], stage0_13[263], stage0_13[264], stage0_13[265], stage0_13[266]},
      {stage0_14[398]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[86],stage1_15[103],stage1_14[131],stage1_13[196]}
   );
   gpc615_5 gpc615 (
      {stage0_13[267], stage0_13[268], stage0_13[269], stage0_13[270], stage0_13[271]},
      {stage0_14[399]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[87],stage1_15[104],stage1_14[132],stage1_13[197]}
   );
   gpc615_5 gpc616 (
      {stage0_13[272], stage0_13[273], stage0_13[274], stage0_13[275], stage0_13[276]},
      {stage0_14[400]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[88],stage1_15[105],stage1_14[133],stage1_13[198]}
   );
   gpc615_5 gpc617 (
      {stage0_13[277], stage0_13[278], stage0_13[279], stage0_13[280], stage0_13[281]},
      {stage0_14[401]},
      {stage0_15[156], stage0_15[157], stage0_15[158], stage0_15[159], stage0_15[160], stage0_15[161]},
      {stage1_17[26],stage1_16[89],stage1_15[106],stage1_14[134],stage1_13[199]}
   );
   gpc615_5 gpc618 (
      {stage0_13[282], stage0_13[283], stage0_13[284], stage0_13[285], stage0_13[286]},
      {stage0_14[402]},
      {stage0_15[162], stage0_15[163], stage0_15[164], stage0_15[165], stage0_15[166], stage0_15[167]},
      {stage1_17[27],stage1_16[90],stage1_15[107],stage1_14[135],stage1_13[200]}
   );
   gpc615_5 gpc619 (
      {stage0_13[287], stage0_13[288], stage0_13[289], stage0_13[290], stage0_13[291]},
      {stage0_14[403]},
      {stage0_15[168], stage0_15[169], stage0_15[170], stage0_15[171], stage0_15[172], stage0_15[173]},
      {stage1_17[28],stage1_16[91],stage1_15[108],stage1_14[136],stage1_13[201]}
   );
   gpc615_5 gpc620 (
      {stage0_13[292], stage0_13[293], stage0_13[294], stage0_13[295], stage0_13[296]},
      {stage0_14[404]},
      {stage0_15[174], stage0_15[175], stage0_15[176], stage0_15[177], stage0_15[178], stage0_15[179]},
      {stage1_17[29],stage1_16[92],stage1_15[109],stage1_14[137],stage1_13[202]}
   );
   gpc615_5 gpc621 (
      {stage0_13[297], stage0_13[298], stage0_13[299], stage0_13[300], stage0_13[301]},
      {stage0_14[405]},
      {stage0_15[180], stage0_15[181], stage0_15[182], stage0_15[183], stage0_15[184], stage0_15[185]},
      {stage1_17[30],stage1_16[93],stage1_15[110],stage1_14[138],stage1_13[203]}
   );
   gpc615_5 gpc622 (
      {stage0_13[302], stage0_13[303], stage0_13[304], stage0_13[305], stage0_13[306]},
      {stage0_14[406]},
      {stage0_15[186], stage0_15[187], stage0_15[188], stage0_15[189], stage0_15[190], stage0_15[191]},
      {stage1_17[31],stage1_16[94],stage1_15[111],stage1_14[139],stage1_13[204]}
   );
   gpc615_5 gpc623 (
      {stage0_13[307], stage0_13[308], stage0_13[309], stage0_13[310], stage0_13[311]},
      {stage0_14[407]},
      {stage0_15[192], stage0_15[193], stage0_15[194], stage0_15[195], stage0_15[196], stage0_15[197]},
      {stage1_17[32],stage1_16[95],stage1_15[112],stage1_14[140],stage1_13[205]}
   );
   gpc615_5 gpc624 (
      {stage0_13[312], stage0_13[313], stage0_13[314], stage0_13[315], stage0_13[316]},
      {stage0_14[408]},
      {stage0_15[198], stage0_15[199], stage0_15[200], stage0_15[201], stage0_15[202], stage0_15[203]},
      {stage1_17[33],stage1_16[96],stage1_15[113],stage1_14[141],stage1_13[206]}
   );
   gpc615_5 gpc625 (
      {stage0_13[317], stage0_13[318], stage0_13[319], stage0_13[320], stage0_13[321]},
      {stage0_14[409]},
      {stage0_15[204], stage0_15[205], stage0_15[206], stage0_15[207], stage0_15[208], stage0_15[209]},
      {stage1_17[34],stage1_16[97],stage1_15[114],stage1_14[142],stage1_13[207]}
   );
   gpc615_5 gpc626 (
      {stage0_13[322], stage0_13[323], stage0_13[324], stage0_13[325], stage0_13[326]},
      {stage0_14[410]},
      {stage0_15[210], stage0_15[211], stage0_15[212], stage0_15[213], stage0_15[214], stage0_15[215]},
      {stage1_17[35],stage1_16[98],stage1_15[115],stage1_14[143],stage1_13[208]}
   );
   gpc615_5 gpc627 (
      {stage0_13[327], stage0_13[328], stage0_13[329], stage0_13[330], stage0_13[331]},
      {stage0_14[411]},
      {stage0_15[216], stage0_15[217], stage0_15[218], stage0_15[219], stage0_15[220], stage0_15[221]},
      {stage1_17[36],stage1_16[99],stage1_15[116],stage1_14[144],stage1_13[209]}
   );
   gpc615_5 gpc628 (
      {stage0_13[332], stage0_13[333], stage0_13[334], stage0_13[335], stage0_13[336]},
      {stage0_14[412]},
      {stage0_15[222], stage0_15[223], stage0_15[224], stage0_15[225], stage0_15[226], stage0_15[227]},
      {stage1_17[37],stage1_16[100],stage1_15[117],stage1_14[145],stage1_13[210]}
   );
   gpc615_5 gpc629 (
      {stage0_13[337], stage0_13[338], stage0_13[339], stage0_13[340], stage0_13[341]},
      {stage0_14[413]},
      {stage0_15[228], stage0_15[229], stage0_15[230], stage0_15[231], stage0_15[232], stage0_15[233]},
      {stage1_17[38],stage1_16[101],stage1_15[118],stage1_14[146],stage1_13[211]}
   );
   gpc615_5 gpc630 (
      {stage0_13[342], stage0_13[343], stage0_13[344], stage0_13[345], stage0_13[346]},
      {stage0_14[414]},
      {stage0_15[234], stage0_15[235], stage0_15[236], stage0_15[237], stage0_15[238], stage0_15[239]},
      {stage1_17[39],stage1_16[102],stage1_15[119],stage1_14[147],stage1_13[212]}
   );
   gpc615_5 gpc631 (
      {stage0_13[347], stage0_13[348], stage0_13[349], stage0_13[350], stage0_13[351]},
      {stage0_14[415]},
      {stage0_15[240], stage0_15[241], stage0_15[242], stage0_15[243], stage0_15[244], stage0_15[245]},
      {stage1_17[40],stage1_16[103],stage1_15[120],stage1_14[148],stage1_13[213]}
   );
   gpc615_5 gpc632 (
      {stage0_13[352], stage0_13[353], stage0_13[354], stage0_13[355], stage0_13[356]},
      {stage0_14[416]},
      {stage0_15[246], stage0_15[247], stage0_15[248], stage0_15[249], stage0_15[250], stage0_15[251]},
      {stage1_17[41],stage1_16[104],stage1_15[121],stage1_14[149],stage1_13[214]}
   );
   gpc615_5 gpc633 (
      {stage0_13[357], stage0_13[358], stage0_13[359], stage0_13[360], stage0_13[361]},
      {stage0_14[417]},
      {stage0_15[252], stage0_15[253], stage0_15[254], stage0_15[255], stage0_15[256], stage0_15[257]},
      {stage1_17[42],stage1_16[105],stage1_15[122],stage1_14[150],stage1_13[215]}
   );
   gpc615_5 gpc634 (
      {stage0_13[362], stage0_13[363], stage0_13[364], stage0_13[365], stage0_13[366]},
      {stage0_14[418]},
      {stage0_15[258], stage0_15[259], stage0_15[260], stage0_15[261], stage0_15[262], stage0_15[263]},
      {stage1_17[43],stage1_16[106],stage1_15[123],stage1_14[151],stage1_13[216]}
   );
   gpc615_5 gpc635 (
      {stage0_13[367], stage0_13[368], stage0_13[369], stage0_13[370], stage0_13[371]},
      {stage0_14[419]},
      {stage0_15[264], stage0_15[265], stage0_15[266], stage0_15[267], stage0_15[268], stage0_15[269]},
      {stage1_17[44],stage1_16[107],stage1_15[124],stage1_14[152],stage1_13[217]}
   );
   gpc615_5 gpc636 (
      {stage0_13[372], stage0_13[373], stage0_13[374], stage0_13[375], stage0_13[376]},
      {stage0_14[420]},
      {stage0_15[270], stage0_15[271], stage0_15[272], stage0_15[273], stage0_15[274], stage0_15[275]},
      {stage1_17[45],stage1_16[108],stage1_15[125],stage1_14[153],stage1_13[218]}
   );
   gpc615_5 gpc637 (
      {stage0_13[377], stage0_13[378], stage0_13[379], stage0_13[380], stage0_13[381]},
      {stage0_14[421]},
      {stage0_15[276], stage0_15[277], stage0_15[278], stage0_15[279], stage0_15[280], stage0_15[281]},
      {stage1_17[46],stage1_16[109],stage1_15[126],stage1_14[154],stage1_13[219]}
   );
   gpc615_5 gpc638 (
      {stage0_13[382], stage0_13[383], stage0_13[384], stage0_13[385], stage0_13[386]},
      {stage0_14[422]},
      {stage0_15[282], stage0_15[283], stage0_15[284], stage0_15[285], stage0_15[286], stage0_15[287]},
      {stage1_17[47],stage1_16[110],stage1_15[127],stage1_14[155],stage1_13[220]}
   );
   gpc615_5 gpc639 (
      {stage0_13[387], stage0_13[388], stage0_13[389], stage0_13[390], stage0_13[391]},
      {stage0_14[423]},
      {stage0_15[288], stage0_15[289], stage0_15[290], stage0_15[291], stage0_15[292], stage0_15[293]},
      {stage1_17[48],stage1_16[111],stage1_15[128],stage1_14[156],stage1_13[221]}
   );
   gpc615_5 gpc640 (
      {stage0_13[392], stage0_13[393], stage0_13[394], stage0_13[395], stage0_13[396]},
      {stage0_14[424]},
      {stage0_15[294], stage0_15[295], stage0_15[296], stage0_15[297], stage0_15[298], stage0_15[299]},
      {stage1_17[49],stage1_16[112],stage1_15[129],stage1_14[157],stage1_13[222]}
   );
   gpc615_5 gpc641 (
      {stage0_13[397], stage0_13[398], stage0_13[399], stage0_13[400], stage0_13[401]},
      {stage0_14[425]},
      {stage0_15[300], stage0_15[301], stage0_15[302], stage0_15[303], stage0_15[304], stage0_15[305]},
      {stage1_17[50],stage1_16[113],stage1_15[130],stage1_14[158],stage1_13[223]}
   );
   gpc615_5 gpc642 (
      {stage0_13[402], stage0_13[403], stage0_13[404], stage0_13[405], stage0_13[406]},
      {stage0_14[426]},
      {stage0_15[306], stage0_15[307], stage0_15[308], stage0_15[309], stage0_15[310], stage0_15[311]},
      {stage1_17[51],stage1_16[114],stage1_15[131],stage1_14[159],stage1_13[224]}
   );
   gpc615_5 gpc643 (
      {stage0_13[407], stage0_13[408], stage0_13[409], stage0_13[410], stage0_13[411]},
      {stage0_14[427]},
      {stage0_15[312], stage0_15[313], stage0_15[314], stage0_15[315], stage0_15[316], stage0_15[317]},
      {stage1_17[52],stage1_16[115],stage1_15[132],stage1_14[160],stage1_13[225]}
   );
   gpc615_5 gpc644 (
      {stage0_13[412], stage0_13[413], stage0_13[414], stage0_13[415], stage0_13[416]},
      {stage0_14[428]},
      {stage0_15[318], stage0_15[319], stage0_15[320], stage0_15[321], stage0_15[322], stage0_15[323]},
      {stage1_17[53],stage1_16[116],stage1_15[133],stage1_14[161],stage1_13[226]}
   );
   gpc615_5 gpc645 (
      {stage0_13[417], stage0_13[418], stage0_13[419], stage0_13[420], stage0_13[421]},
      {stage0_14[429]},
      {stage0_15[324], stage0_15[325], stage0_15[326], stage0_15[327], stage0_15[328], stage0_15[329]},
      {stage1_17[54],stage1_16[117],stage1_15[134],stage1_14[162],stage1_13[227]}
   );
   gpc615_5 gpc646 (
      {stage0_13[422], stage0_13[423], stage0_13[424], stage0_13[425], stage0_13[426]},
      {stage0_14[430]},
      {stage0_15[330], stage0_15[331], stage0_15[332], stage0_15[333], stage0_15[334], stage0_15[335]},
      {stage1_17[55],stage1_16[118],stage1_15[135],stage1_14[163],stage1_13[228]}
   );
   gpc615_5 gpc647 (
      {stage0_13[427], stage0_13[428], stage0_13[429], stage0_13[430], stage0_13[431]},
      {stage0_14[431]},
      {stage0_15[336], stage0_15[337], stage0_15[338], stage0_15[339], stage0_15[340], stage0_15[341]},
      {stage1_17[56],stage1_16[119],stage1_15[136],stage1_14[164],stage1_13[229]}
   );
   gpc615_5 gpc648 (
      {stage0_13[432], stage0_13[433], stage0_13[434], stage0_13[435], stage0_13[436]},
      {stage0_14[432]},
      {stage0_15[342], stage0_15[343], stage0_15[344], stage0_15[345], stage0_15[346], stage0_15[347]},
      {stage1_17[57],stage1_16[120],stage1_15[137],stage1_14[165],stage1_13[230]}
   );
   gpc615_5 gpc649 (
      {stage0_13[437], stage0_13[438], stage0_13[439], stage0_13[440], stage0_13[441]},
      {stage0_14[433]},
      {stage0_15[348], stage0_15[349], stage0_15[350], stage0_15[351], stage0_15[352], stage0_15[353]},
      {stage1_17[58],stage1_16[121],stage1_15[138],stage1_14[166],stage1_13[231]}
   );
   gpc615_5 gpc650 (
      {stage0_13[442], stage0_13[443], stage0_13[444], stage0_13[445], stage0_13[446]},
      {stage0_14[434]},
      {stage0_15[354], stage0_15[355], stage0_15[356], stage0_15[357], stage0_15[358], stage0_15[359]},
      {stage1_17[59],stage1_16[122],stage1_15[139],stage1_14[167],stage1_13[232]}
   );
   gpc615_5 gpc651 (
      {stage0_13[447], stage0_13[448], stage0_13[449], stage0_13[450], stage0_13[451]},
      {stage0_14[435]},
      {stage0_15[360], stage0_15[361], stage0_15[362], stage0_15[363], stage0_15[364], stage0_15[365]},
      {stage1_17[60],stage1_16[123],stage1_15[140],stage1_14[168],stage1_13[233]}
   );
   gpc615_5 gpc652 (
      {stage0_13[452], stage0_13[453], stage0_13[454], stage0_13[455], stage0_13[456]},
      {stage0_14[436]},
      {stage0_15[366], stage0_15[367], stage0_15[368], stage0_15[369], stage0_15[370], stage0_15[371]},
      {stage1_17[61],stage1_16[124],stage1_15[141],stage1_14[169],stage1_13[234]}
   );
   gpc615_5 gpc653 (
      {stage0_13[457], stage0_13[458], stage0_13[459], stage0_13[460], stage0_13[461]},
      {stage0_14[437]},
      {stage0_15[372], stage0_15[373], stage0_15[374], stage0_15[375], stage0_15[376], stage0_15[377]},
      {stage1_17[62],stage1_16[125],stage1_15[142],stage1_14[170],stage1_13[235]}
   );
   gpc615_5 gpc654 (
      {stage0_13[462], stage0_13[463], stage0_13[464], stage0_13[465], stage0_13[466]},
      {stage0_14[438]},
      {stage0_15[378], stage0_15[379], stage0_15[380], stage0_15[381], stage0_15[382], stage0_15[383]},
      {stage1_17[63],stage1_16[126],stage1_15[143],stage1_14[171],stage1_13[236]}
   );
   gpc1_1 gpc655 (
      {stage0_0[509]},
      {stage1_0[98]}
   );
   gpc1_1 gpc656 (
      {stage0_0[510]},
      {stage1_0[99]}
   );
   gpc1_1 gpc657 (
      {stage0_0[511]},
      {stage1_0[100]}
   );
   gpc1_1 gpc658 (
      {stage0_1[476]},
      {stage1_1[144]}
   );
   gpc1_1 gpc659 (
      {stage0_1[477]},
      {stage1_1[145]}
   );
   gpc1_1 gpc660 (
      {stage0_1[478]},
      {stage1_1[146]}
   );
   gpc1_1 gpc661 (
      {stage0_1[479]},
      {stage1_1[147]}
   );
   gpc1_1 gpc662 (
      {stage0_1[480]},
      {stage1_1[148]}
   );
   gpc1_1 gpc663 (
      {stage0_1[481]},
      {stage1_1[149]}
   );
   gpc1_1 gpc664 (
      {stage0_1[482]},
      {stage1_1[150]}
   );
   gpc1_1 gpc665 (
      {stage0_1[483]},
      {stage1_1[151]}
   );
   gpc1_1 gpc666 (
      {stage0_1[484]},
      {stage1_1[152]}
   );
   gpc1_1 gpc667 (
      {stage0_1[485]},
      {stage1_1[153]}
   );
   gpc1_1 gpc668 (
      {stage0_1[486]},
      {stage1_1[154]}
   );
   gpc1_1 gpc669 (
      {stage0_1[487]},
      {stage1_1[155]}
   );
   gpc1_1 gpc670 (
      {stage0_1[488]},
      {stage1_1[156]}
   );
   gpc1_1 gpc671 (
      {stage0_1[489]},
      {stage1_1[157]}
   );
   gpc1_1 gpc672 (
      {stage0_1[490]},
      {stage1_1[158]}
   );
   gpc1_1 gpc673 (
      {stage0_1[491]},
      {stage1_1[159]}
   );
   gpc1_1 gpc674 (
      {stage0_1[492]},
      {stage1_1[160]}
   );
   gpc1_1 gpc675 (
      {stage0_1[493]},
      {stage1_1[161]}
   );
   gpc1_1 gpc676 (
      {stage0_1[494]},
      {stage1_1[162]}
   );
   gpc1_1 gpc677 (
      {stage0_1[495]},
      {stage1_1[163]}
   );
   gpc1_1 gpc678 (
      {stage0_1[496]},
      {stage1_1[164]}
   );
   gpc1_1 gpc679 (
      {stage0_1[497]},
      {stage1_1[165]}
   );
   gpc1_1 gpc680 (
      {stage0_1[498]},
      {stage1_1[166]}
   );
   gpc1_1 gpc681 (
      {stage0_1[499]},
      {stage1_1[167]}
   );
   gpc1_1 gpc682 (
      {stage0_1[500]},
      {stage1_1[168]}
   );
   gpc1_1 gpc683 (
      {stage0_1[501]},
      {stage1_1[169]}
   );
   gpc1_1 gpc684 (
      {stage0_1[502]},
      {stage1_1[170]}
   );
   gpc1_1 gpc685 (
      {stage0_1[503]},
      {stage1_1[171]}
   );
   gpc1_1 gpc686 (
      {stage0_1[504]},
      {stage1_1[172]}
   );
   gpc1_1 gpc687 (
      {stage0_1[505]},
      {stage1_1[173]}
   );
   gpc1_1 gpc688 (
      {stage0_1[506]},
      {stage1_1[174]}
   );
   gpc1_1 gpc689 (
      {stage0_1[507]},
      {stage1_1[175]}
   );
   gpc1_1 gpc690 (
      {stage0_1[508]},
      {stage1_1[176]}
   );
   gpc1_1 gpc691 (
      {stage0_1[509]},
      {stage1_1[177]}
   );
   gpc1_1 gpc692 (
      {stage0_1[510]},
      {stage1_1[178]}
   );
   gpc1_1 gpc693 (
      {stage0_1[511]},
      {stage1_1[179]}
   );
   gpc1_1 gpc694 (
      {stage0_3[466]},
      {stage1_3[200]}
   );
   gpc1_1 gpc695 (
      {stage0_3[467]},
      {stage1_3[201]}
   );
   gpc1_1 gpc696 (
      {stage0_3[468]},
      {stage1_3[202]}
   );
   gpc1_1 gpc697 (
      {stage0_3[469]},
      {stage1_3[203]}
   );
   gpc1_1 gpc698 (
      {stage0_3[470]},
      {stage1_3[204]}
   );
   gpc1_1 gpc699 (
      {stage0_3[471]},
      {stage1_3[205]}
   );
   gpc1_1 gpc700 (
      {stage0_3[472]},
      {stage1_3[206]}
   );
   gpc1_1 gpc701 (
      {stage0_3[473]},
      {stage1_3[207]}
   );
   gpc1_1 gpc702 (
      {stage0_3[474]},
      {stage1_3[208]}
   );
   gpc1_1 gpc703 (
      {stage0_3[475]},
      {stage1_3[209]}
   );
   gpc1_1 gpc704 (
      {stage0_3[476]},
      {stage1_3[210]}
   );
   gpc1_1 gpc705 (
      {stage0_3[477]},
      {stage1_3[211]}
   );
   gpc1_1 gpc706 (
      {stage0_3[478]},
      {stage1_3[212]}
   );
   gpc1_1 gpc707 (
      {stage0_3[479]},
      {stage1_3[213]}
   );
   gpc1_1 gpc708 (
      {stage0_3[480]},
      {stage1_3[214]}
   );
   gpc1_1 gpc709 (
      {stage0_3[481]},
      {stage1_3[215]}
   );
   gpc1_1 gpc710 (
      {stage0_3[482]},
      {stage1_3[216]}
   );
   gpc1_1 gpc711 (
      {stage0_3[483]},
      {stage1_3[217]}
   );
   gpc1_1 gpc712 (
      {stage0_3[484]},
      {stage1_3[218]}
   );
   gpc1_1 gpc713 (
      {stage0_3[485]},
      {stage1_3[219]}
   );
   gpc1_1 gpc714 (
      {stage0_3[486]},
      {stage1_3[220]}
   );
   gpc1_1 gpc715 (
      {stage0_3[487]},
      {stage1_3[221]}
   );
   gpc1_1 gpc716 (
      {stage0_3[488]},
      {stage1_3[222]}
   );
   gpc1_1 gpc717 (
      {stage0_3[489]},
      {stage1_3[223]}
   );
   gpc1_1 gpc718 (
      {stage0_3[490]},
      {stage1_3[224]}
   );
   gpc1_1 gpc719 (
      {stage0_3[491]},
      {stage1_3[225]}
   );
   gpc1_1 gpc720 (
      {stage0_3[492]},
      {stage1_3[226]}
   );
   gpc1_1 gpc721 (
      {stage0_3[493]},
      {stage1_3[227]}
   );
   gpc1_1 gpc722 (
      {stage0_3[494]},
      {stage1_3[228]}
   );
   gpc1_1 gpc723 (
      {stage0_3[495]},
      {stage1_3[229]}
   );
   gpc1_1 gpc724 (
      {stage0_3[496]},
      {stage1_3[230]}
   );
   gpc1_1 gpc725 (
      {stage0_3[497]},
      {stage1_3[231]}
   );
   gpc1_1 gpc726 (
      {stage0_3[498]},
      {stage1_3[232]}
   );
   gpc1_1 gpc727 (
      {stage0_3[499]},
      {stage1_3[233]}
   );
   gpc1_1 gpc728 (
      {stage0_3[500]},
      {stage1_3[234]}
   );
   gpc1_1 gpc729 (
      {stage0_3[501]},
      {stage1_3[235]}
   );
   gpc1_1 gpc730 (
      {stage0_3[502]},
      {stage1_3[236]}
   );
   gpc1_1 gpc731 (
      {stage0_3[503]},
      {stage1_3[237]}
   );
   gpc1_1 gpc732 (
      {stage0_3[504]},
      {stage1_3[238]}
   );
   gpc1_1 gpc733 (
      {stage0_3[505]},
      {stage1_3[239]}
   );
   gpc1_1 gpc734 (
      {stage0_3[506]},
      {stage1_3[240]}
   );
   gpc1_1 gpc735 (
      {stage0_3[507]},
      {stage1_3[241]}
   );
   gpc1_1 gpc736 (
      {stage0_3[508]},
      {stage1_3[242]}
   );
   gpc1_1 gpc737 (
      {stage0_3[509]},
      {stage1_3[243]}
   );
   gpc1_1 gpc738 (
      {stage0_3[510]},
      {stage1_3[244]}
   );
   gpc1_1 gpc739 (
      {stage0_3[511]},
      {stage1_3[245]}
   );
   gpc1_1 gpc740 (
      {stage0_5[505]},
      {stage1_5[211]}
   );
   gpc1_1 gpc741 (
      {stage0_5[506]},
      {stage1_5[212]}
   );
   gpc1_1 gpc742 (
      {stage0_5[507]},
      {stage1_5[213]}
   );
   gpc1_1 gpc743 (
      {stage0_5[508]},
      {stage1_5[214]}
   );
   gpc1_1 gpc744 (
      {stage0_5[509]},
      {stage1_5[215]}
   );
   gpc1_1 gpc745 (
      {stage0_5[510]},
      {stage1_5[216]}
   );
   gpc1_1 gpc746 (
      {stage0_5[511]},
      {stage1_5[217]}
   );
   gpc1_1 gpc747 (
      {stage0_6[505]},
      {stage1_6[200]}
   );
   gpc1_1 gpc748 (
      {stage0_6[506]},
      {stage1_6[201]}
   );
   gpc1_1 gpc749 (
      {stage0_6[507]},
      {stage1_6[202]}
   );
   gpc1_1 gpc750 (
      {stage0_6[508]},
      {stage1_6[203]}
   );
   gpc1_1 gpc751 (
      {stage0_6[509]},
      {stage1_6[204]}
   );
   gpc1_1 gpc752 (
      {stage0_6[510]},
      {stage1_6[205]}
   );
   gpc1_1 gpc753 (
      {stage0_6[511]},
      {stage1_6[206]}
   );
   gpc1_1 gpc754 (
      {stage0_7[501]},
      {stage1_7[196]}
   );
   gpc1_1 gpc755 (
      {stage0_7[502]},
      {stage1_7[197]}
   );
   gpc1_1 gpc756 (
      {stage0_7[503]},
      {stage1_7[198]}
   );
   gpc1_1 gpc757 (
      {stage0_7[504]},
      {stage1_7[199]}
   );
   gpc1_1 gpc758 (
      {stage0_7[505]},
      {stage1_7[200]}
   );
   gpc1_1 gpc759 (
      {stage0_7[506]},
      {stage1_7[201]}
   );
   gpc1_1 gpc760 (
      {stage0_7[507]},
      {stage1_7[202]}
   );
   gpc1_1 gpc761 (
      {stage0_7[508]},
      {stage1_7[203]}
   );
   gpc1_1 gpc762 (
      {stage0_7[509]},
      {stage1_7[204]}
   );
   gpc1_1 gpc763 (
      {stage0_7[510]},
      {stage1_7[205]}
   );
   gpc1_1 gpc764 (
      {stage0_7[511]},
      {stage1_7[206]}
   );
   gpc1_1 gpc765 (
      {stage0_9[476]},
      {stage1_9[228]}
   );
   gpc1_1 gpc766 (
      {stage0_9[477]},
      {stage1_9[229]}
   );
   gpc1_1 gpc767 (
      {stage0_9[478]},
      {stage1_9[230]}
   );
   gpc1_1 gpc768 (
      {stage0_9[479]},
      {stage1_9[231]}
   );
   gpc1_1 gpc769 (
      {stage0_9[480]},
      {stage1_9[232]}
   );
   gpc1_1 gpc770 (
      {stage0_9[481]},
      {stage1_9[233]}
   );
   gpc1_1 gpc771 (
      {stage0_9[482]},
      {stage1_9[234]}
   );
   gpc1_1 gpc772 (
      {stage0_9[483]},
      {stage1_9[235]}
   );
   gpc1_1 gpc773 (
      {stage0_9[484]},
      {stage1_9[236]}
   );
   gpc1_1 gpc774 (
      {stage0_9[485]},
      {stage1_9[237]}
   );
   gpc1_1 gpc775 (
      {stage0_9[486]},
      {stage1_9[238]}
   );
   gpc1_1 gpc776 (
      {stage0_9[487]},
      {stage1_9[239]}
   );
   gpc1_1 gpc777 (
      {stage0_9[488]},
      {stage1_9[240]}
   );
   gpc1_1 gpc778 (
      {stage0_9[489]},
      {stage1_9[241]}
   );
   gpc1_1 gpc779 (
      {stage0_9[490]},
      {stage1_9[242]}
   );
   gpc1_1 gpc780 (
      {stage0_9[491]},
      {stage1_9[243]}
   );
   gpc1_1 gpc781 (
      {stage0_9[492]},
      {stage1_9[244]}
   );
   gpc1_1 gpc782 (
      {stage0_9[493]},
      {stage1_9[245]}
   );
   gpc1_1 gpc783 (
      {stage0_9[494]},
      {stage1_9[246]}
   );
   gpc1_1 gpc784 (
      {stage0_9[495]},
      {stage1_9[247]}
   );
   gpc1_1 gpc785 (
      {stage0_9[496]},
      {stage1_9[248]}
   );
   gpc1_1 gpc786 (
      {stage0_9[497]},
      {stage1_9[249]}
   );
   gpc1_1 gpc787 (
      {stage0_9[498]},
      {stage1_9[250]}
   );
   gpc1_1 gpc788 (
      {stage0_9[499]},
      {stage1_9[251]}
   );
   gpc1_1 gpc789 (
      {stage0_9[500]},
      {stage1_9[252]}
   );
   gpc1_1 gpc790 (
      {stage0_9[501]},
      {stage1_9[253]}
   );
   gpc1_1 gpc791 (
      {stage0_9[502]},
      {stage1_9[254]}
   );
   gpc1_1 gpc792 (
      {stage0_9[503]},
      {stage1_9[255]}
   );
   gpc1_1 gpc793 (
      {stage0_9[504]},
      {stage1_9[256]}
   );
   gpc1_1 gpc794 (
      {stage0_9[505]},
      {stage1_9[257]}
   );
   gpc1_1 gpc795 (
      {stage0_9[506]},
      {stage1_9[258]}
   );
   gpc1_1 gpc796 (
      {stage0_9[507]},
      {stage1_9[259]}
   );
   gpc1_1 gpc797 (
      {stage0_9[508]},
      {stage1_9[260]}
   );
   gpc1_1 gpc798 (
      {stage0_9[509]},
      {stage1_9[261]}
   );
   gpc1_1 gpc799 (
      {stage0_9[510]},
      {stage1_9[262]}
   );
   gpc1_1 gpc800 (
      {stage0_9[511]},
      {stage1_9[263]}
   );
   gpc1_1 gpc801 (
      {stage0_10[504]},
      {stage1_10[202]}
   );
   gpc1_1 gpc802 (
      {stage0_10[505]},
      {stage1_10[203]}
   );
   gpc1_1 gpc803 (
      {stage0_10[506]},
      {stage1_10[204]}
   );
   gpc1_1 gpc804 (
      {stage0_10[507]},
      {stage1_10[205]}
   );
   gpc1_1 gpc805 (
      {stage0_10[508]},
      {stage1_10[206]}
   );
   gpc1_1 gpc806 (
      {stage0_10[509]},
      {stage1_10[207]}
   );
   gpc1_1 gpc807 (
      {stage0_10[510]},
      {stage1_10[208]}
   );
   gpc1_1 gpc808 (
      {stage0_10[511]},
      {stage1_10[209]}
   );
   gpc1_1 gpc809 (
      {stage0_11[506]},
      {stage1_11[184]}
   );
   gpc1_1 gpc810 (
      {stage0_11[507]},
      {stage1_11[185]}
   );
   gpc1_1 gpc811 (
      {stage0_11[508]},
      {stage1_11[186]}
   );
   gpc1_1 gpc812 (
      {stage0_11[509]},
      {stage1_11[187]}
   );
   gpc1_1 gpc813 (
      {stage0_11[510]},
      {stage1_11[188]}
   );
   gpc1_1 gpc814 (
      {stage0_11[511]},
      {stage1_11[189]}
   );
   gpc1_1 gpc815 (
      {stage0_13[467]},
      {stage1_13[237]}
   );
   gpc1_1 gpc816 (
      {stage0_13[468]},
      {stage1_13[238]}
   );
   gpc1_1 gpc817 (
      {stage0_13[469]},
      {stage1_13[239]}
   );
   gpc1_1 gpc818 (
      {stage0_13[470]},
      {stage1_13[240]}
   );
   gpc1_1 gpc819 (
      {stage0_13[471]},
      {stage1_13[241]}
   );
   gpc1_1 gpc820 (
      {stage0_13[472]},
      {stage1_13[242]}
   );
   gpc1_1 gpc821 (
      {stage0_13[473]},
      {stage1_13[243]}
   );
   gpc1_1 gpc822 (
      {stage0_13[474]},
      {stage1_13[244]}
   );
   gpc1_1 gpc823 (
      {stage0_13[475]},
      {stage1_13[245]}
   );
   gpc1_1 gpc824 (
      {stage0_13[476]},
      {stage1_13[246]}
   );
   gpc1_1 gpc825 (
      {stage0_13[477]},
      {stage1_13[247]}
   );
   gpc1_1 gpc826 (
      {stage0_13[478]},
      {stage1_13[248]}
   );
   gpc1_1 gpc827 (
      {stage0_13[479]},
      {stage1_13[249]}
   );
   gpc1_1 gpc828 (
      {stage0_13[480]},
      {stage1_13[250]}
   );
   gpc1_1 gpc829 (
      {stage0_13[481]},
      {stage1_13[251]}
   );
   gpc1_1 gpc830 (
      {stage0_13[482]},
      {stage1_13[252]}
   );
   gpc1_1 gpc831 (
      {stage0_13[483]},
      {stage1_13[253]}
   );
   gpc1_1 gpc832 (
      {stage0_13[484]},
      {stage1_13[254]}
   );
   gpc1_1 gpc833 (
      {stage0_13[485]},
      {stage1_13[255]}
   );
   gpc1_1 gpc834 (
      {stage0_13[486]},
      {stage1_13[256]}
   );
   gpc1_1 gpc835 (
      {stage0_13[487]},
      {stage1_13[257]}
   );
   gpc1_1 gpc836 (
      {stage0_13[488]},
      {stage1_13[258]}
   );
   gpc1_1 gpc837 (
      {stage0_13[489]},
      {stage1_13[259]}
   );
   gpc1_1 gpc838 (
      {stage0_13[490]},
      {stage1_13[260]}
   );
   gpc1_1 gpc839 (
      {stage0_13[491]},
      {stage1_13[261]}
   );
   gpc1_1 gpc840 (
      {stage0_13[492]},
      {stage1_13[262]}
   );
   gpc1_1 gpc841 (
      {stage0_13[493]},
      {stage1_13[263]}
   );
   gpc1_1 gpc842 (
      {stage0_13[494]},
      {stage1_13[264]}
   );
   gpc1_1 gpc843 (
      {stage0_13[495]},
      {stage1_13[265]}
   );
   gpc1_1 gpc844 (
      {stage0_13[496]},
      {stage1_13[266]}
   );
   gpc1_1 gpc845 (
      {stage0_13[497]},
      {stage1_13[267]}
   );
   gpc1_1 gpc846 (
      {stage0_13[498]},
      {stage1_13[268]}
   );
   gpc1_1 gpc847 (
      {stage0_13[499]},
      {stage1_13[269]}
   );
   gpc1_1 gpc848 (
      {stage0_13[500]},
      {stage1_13[270]}
   );
   gpc1_1 gpc849 (
      {stage0_13[501]},
      {stage1_13[271]}
   );
   gpc1_1 gpc850 (
      {stage0_13[502]},
      {stage1_13[272]}
   );
   gpc1_1 gpc851 (
      {stage0_13[503]},
      {stage1_13[273]}
   );
   gpc1_1 gpc852 (
      {stage0_13[504]},
      {stage1_13[274]}
   );
   gpc1_1 gpc853 (
      {stage0_13[505]},
      {stage1_13[275]}
   );
   gpc1_1 gpc854 (
      {stage0_13[506]},
      {stage1_13[276]}
   );
   gpc1_1 gpc855 (
      {stage0_13[507]},
      {stage1_13[277]}
   );
   gpc1_1 gpc856 (
      {stage0_13[508]},
      {stage1_13[278]}
   );
   gpc1_1 gpc857 (
      {stage0_13[509]},
      {stage1_13[279]}
   );
   gpc1_1 gpc858 (
      {stage0_13[510]},
      {stage1_13[280]}
   );
   gpc1_1 gpc859 (
      {stage0_13[511]},
      {stage1_13[281]}
   );
   gpc1_1 gpc860 (
      {stage0_14[439]},
      {stage1_14[172]}
   );
   gpc1_1 gpc861 (
      {stage0_14[440]},
      {stage1_14[173]}
   );
   gpc1_1 gpc862 (
      {stage0_14[441]},
      {stage1_14[174]}
   );
   gpc1_1 gpc863 (
      {stage0_14[442]},
      {stage1_14[175]}
   );
   gpc1_1 gpc864 (
      {stage0_14[443]},
      {stage1_14[176]}
   );
   gpc1_1 gpc865 (
      {stage0_14[444]},
      {stage1_14[177]}
   );
   gpc1_1 gpc866 (
      {stage0_14[445]},
      {stage1_14[178]}
   );
   gpc1_1 gpc867 (
      {stage0_14[446]},
      {stage1_14[179]}
   );
   gpc1_1 gpc868 (
      {stage0_14[447]},
      {stage1_14[180]}
   );
   gpc1_1 gpc869 (
      {stage0_14[448]},
      {stage1_14[181]}
   );
   gpc1_1 gpc870 (
      {stage0_14[449]},
      {stage1_14[182]}
   );
   gpc1_1 gpc871 (
      {stage0_14[450]},
      {stage1_14[183]}
   );
   gpc1_1 gpc872 (
      {stage0_14[451]},
      {stage1_14[184]}
   );
   gpc1_1 gpc873 (
      {stage0_14[452]},
      {stage1_14[185]}
   );
   gpc1_1 gpc874 (
      {stage0_14[453]},
      {stage1_14[186]}
   );
   gpc1_1 gpc875 (
      {stage0_14[454]},
      {stage1_14[187]}
   );
   gpc1_1 gpc876 (
      {stage0_14[455]},
      {stage1_14[188]}
   );
   gpc1_1 gpc877 (
      {stage0_14[456]},
      {stage1_14[189]}
   );
   gpc1_1 gpc878 (
      {stage0_14[457]},
      {stage1_14[190]}
   );
   gpc1_1 gpc879 (
      {stage0_14[458]},
      {stage1_14[191]}
   );
   gpc1_1 gpc880 (
      {stage0_14[459]},
      {stage1_14[192]}
   );
   gpc1_1 gpc881 (
      {stage0_14[460]},
      {stage1_14[193]}
   );
   gpc1_1 gpc882 (
      {stage0_14[461]},
      {stage1_14[194]}
   );
   gpc1_1 gpc883 (
      {stage0_14[462]},
      {stage1_14[195]}
   );
   gpc1_1 gpc884 (
      {stage0_14[463]},
      {stage1_14[196]}
   );
   gpc1_1 gpc885 (
      {stage0_14[464]},
      {stage1_14[197]}
   );
   gpc1_1 gpc886 (
      {stage0_14[465]},
      {stage1_14[198]}
   );
   gpc1_1 gpc887 (
      {stage0_14[466]},
      {stage1_14[199]}
   );
   gpc1_1 gpc888 (
      {stage0_14[467]},
      {stage1_14[200]}
   );
   gpc1_1 gpc889 (
      {stage0_14[468]},
      {stage1_14[201]}
   );
   gpc1_1 gpc890 (
      {stage0_14[469]},
      {stage1_14[202]}
   );
   gpc1_1 gpc891 (
      {stage0_14[470]},
      {stage1_14[203]}
   );
   gpc1_1 gpc892 (
      {stage0_14[471]},
      {stage1_14[204]}
   );
   gpc1_1 gpc893 (
      {stage0_14[472]},
      {stage1_14[205]}
   );
   gpc1_1 gpc894 (
      {stage0_14[473]},
      {stage1_14[206]}
   );
   gpc1_1 gpc895 (
      {stage0_14[474]},
      {stage1_14[207]}
   );
   gpc1_1 gpc896 (
      {stage0_14[475]},
      {stage1_14[208]}
   );
   gpc1_1 gpc897 (
      {stage0_14[476]},
      {stage1_14[209]}
   );
   gpc1_1 gpc898 (
      {stage0_14[477]},
      {stage1_14[210]}
   );
   gpc1_1 gpc899 (
      {stage0_14[478]},
      {stage1_14[211]}
   );
   gpc1_1 gpc900 (
      {stage0_14[479]},
      {stage1_14[212]}
   );
   gpc1_1 gpc901 (
      {stage0_14[480]},
      {stage1_14[213]}
   );
   gpc1_1 gpc902 (
      {stage0_14[481]},
      {stage1_14[214]}
   );
   gpc1_1 gpc903 (
      {stage0_14[482]},
      {stage1_14[215]}
   );
   gpc1_1 gpc904 (
      {stage0_14[483]},
      {stage1_14[216]}
   );
   gpc1_1 gpc905 (
      {stage0_14[484]},
      {stage1_14[217]}
   );
   gpc1_1 gpc906 (
      {stage0_14[485]},
      {stage1_14[218]}
   );
   gpc1_1 gpc907 (
      {stage0_14[486]},
      {stage1_14[219]}
   );
   gpc1_1 gpc908 (
      {stage0_14[487]},
      {stage1_14[220]}
   );
   gpc1_1 gpc909 (
      {stage0_14[488]},
      {stage1_14[221]}
   );
   gpc1_1 gpc910 (
      {stage0_14[489]},
      {stage1_14[222]}
   );
   gpc1_1 gpc911 (
      {stage0_14[490]},
      {stage1_14[223]}
   );
   gpc1_1 gpc912 (
      {stage0_14[491]},
      {stage1_14[224]}
   );
   gpc1_1 gpc913 (
      {stage0_14[492]},
      {stage1_14[225]}
   );
   gpc1_1 gpc914 (
      {stage0_14[493]},
      {stage1_14[226]}
   );
   gpc1_1 gpc915 (
      {stage0_14[494]},
      {stage1_14[227]}
   );
   gpc1_1 gpc916 (
      {stage0_14[495]},
      {stage1_14[228]}
   );
   gpc1_1 gpc917 (
      {stage0_14[496]},
      {stage1_14[229]}
   );
   gpc1_1 gpc918 (
      {stage0_14[497]},
      {stage1_14[230]}
   );
   gpc1_1 gpc919 (
      {stage0_14[498]},
      {stage1_14[231]}
   );
   gpc1_1 gpc920 (
      {stage0_14[499]},
      {stage1_14[232]}
   );
   gpc1_1 gpc921 (
      {stage0_14[500]},
      {stage1_14[233]}
   );
   gpc1_1 gpc922 (
      {stage0_14[501]},
      {stage1_14[234]}
   );
   gpc1_1 gpc923 (
      {stage0_14[502]},
      {stage1_14[235]}
   );
   gpc1_1 gpc924 (
      {stage0_14[503]},
      {stage1_14[236]}
   );
   gpc1_1 gpc925 (
      {stage0_14[504]},
      {stage1_14[237]}
   );
   gpc1_1 gpc926 (
      {stage0_14[505]},
      {stage1_14[238]}
   );
   gpc1_1 gpc927 (
      {stage0_14[506]},
      {stage1_14[239]}
   );
   gpc1_1 gpc928 (
      {stage0_14[507]},
      {stage1_14[240]}
   );
   gpc1_1 gpc929 (
      {stage0_14[508]},
      {stage1_14[241]}
   );
   gpc1_1 gpc930 (
      {stage0_14[509]},
      {stage1_14[242]}
   );
   gpc1_1 gpc931 (
      {stage0_14[510]},
      {stage1_14[243]}
   );
   gpc1_1 gpc932 (
      {stage0_14[511]},
      {stage1_14[244]}
   );
   gpc1_1 gpc933 (
      {stage0_15[384]},
      {stage1_15[144]}
   );
   gpc1_1 gpc934 (
      {stage0_15[385]},
      {stage1_15[145]}
   );
   gpc1_1 gpc935 (
      {stage0_15[386]},
      {stage1_15[146]}
   );
   gpc1_1 gpc936 (
      {stage0_15[387]},
      {stage1_15[147]}
   );
   gpc1_1 gpc937 (
      {stage0_15[388]},
      {stage1_15[148]}
   );
   gpc1_1 gpc938 (
      {stage0_15[389]},
      {stage1_15[149]}
   );
   gpc1_1 gpc939 (
      {stage0_15[390]},
      {stage1_15[150]}
   );
   gpc1_1 gpc940 (
      {stage0_15[391]},
      {stage1_15[151]}
   );
   gpc1_1 gpc941 (
      {stage0_15[392]},
      {stage1_15[152]}
   );
   gpc1_1 gpc942 (
      {stage0_15[393]},
      {stage1_15[153]}
   );
   gpc1_1 gpc943 (
      {stage0_15[394]},
      {stage1_15[154]}
   );
   gpc1_1 gpc944 (
      {stage0_15[395]},
      {stage1_15[155]}
   );
   gpc1_1 gpc945 (
      {stage0_15[396]},
      {stage1_15[156]}
   );
   gpc1_1 gpc946 (
      {stage0_15[397]},
      {stage1_15[157]}
   );
   gpc1_1 gpc947 (
      {stage0_15[398]},
      {stage1_15[158]}
   );
   gpc1_1 gpc948 (
      {stage0_15[399]},
      {stage1_15[159]}
   );
   gpc1_1 gpc949 (
      {stage0_15[400]},
      {stage1_15[160]}
   );
   gpc1_1 gpc950 (
      {stage0_15[401]},
      {stage1_15[161]}
   );
   gpc1_1 gpc951 (
      {stage0_15[402]},
      {stage1_15[162]}
   );
   gpc1_1 gpc952 (
      {stage0_15[403]},
      {stage1_15[163]}
   );
   gpc1_1 gpc953 (
      {stage0_15[404]},
      {stage1_15[164]}
   );
   gpc1_1 gpc954 (
      {stage0_15[405]},
      {stage1_15[165]}
   );
   gpc1_1 gpc955 (
      {stage0_15[406]},
      {stage1_15[166]}
   );
   gpc1_1 gpc956 (
      {stage0_15[407]},
      {stage1_15[167]}
   );
   gpc1_1 gpc957 (
      {stage0_15[408]},
      {stage1_15[168]}
   );
   gpc1_1 gpc958 (
      {stage0_15[409]},
      {stage1_15[169]}
   );
   gpc1_1 gpc959 (
      {stage0_15[410]},
      {stage1_15[170]}
   );
   gpc1_1 gpc960 (
      {stage0_15[411]},
      {stage1_15[171]}
   );
   gpc1_1 gpc961 (
      {stage0_15[412]},
      {stage1_15[172]}
   );
   gpc1_1 gpc962 (
      {stage0_15[413]},
      {stage1_15[173]}
   );
   gpc1_1 gpc963 (
      {stage0_15[414]},
      {stage1_15[174]}
   );
   gpc1_1 gpc964 (
      {stage0_15[415]},
      {stage1_15[175]}
   );
   gpc1_1 gpc965 (
      {stage0_15[416]},
      {stage1_15[176]}
   );
   gpc1_1 gpc966 (
      {stage0_15[417]},
      {stage1_15[177]}
   );
   gpc1_1 gpc967 (
      {stage0_15[418]},
      {stage1_15[178]}
   );
   gpc1_1 gpc968 (
      {stage0_15[419]},
      {stage1_15[179]}
   );
   gpc1_1 gpc969 (
      {stage0_15[420]},
      {stage1_15[180]}
   );
   gpc1_1 gpc970 (
      {stage0_15[421]},
      {stage1_15[181]}
   );
   gpc1_1 gpc971 (
      {stage0_15[422]},
      {stage1_15[182]}
   );
   gpc1_1 gpc972 (
      {stage0_15[423]},
      {stage1_15[183]}
   );
   gpc1_1 gpc973 (
      {stage0_15[424]},
      {stage1_15[184]}
   );
   gpc1_1 gpc974 (
      {stage0_15[425]},
      {stage1_15[185]}
   );
   gpc1_1 gpc975 (
      {stage0_15[426]},
      {stage1_15[186]}
   );
   gpc1_1 gpc976 (
      {stage0_15[427]},
      {stage1_15[187]}
   );
   gpc1_1 gpc977 (
      {stage0_15[428]},
      {stage1_15[188]}
   );
   gpc1_1 gpc978 (
      {stage0_15[429]},
      {stage1_15[189]}
   );
   gpc1_1 gpc979 (
      {stage0_15[430]},
      {stage1_15[190]}
   );
   gpc1_1 gpc980 (
      {stage0_15[431]},
      {stage1_15[191]}
   );
   gpc1_1 gpc981 (
      {stage0_15[432]},
      {stage1_15[192]}
   );
   gpc1_1 gpc982 (
      {stage0_15[433]},
      {stage1_15[193]}
   );
   gpc1_1 gpc983 (
      {stage0_15[434]},
      {stage1_15[194]}
   );
   gpc1_1 gpc984 (
      {stage0_15[435]},
      {stage1_15[195]}
   );
   gpc1_1 gpc985 (
      {stage0_15[436]},
      {stage1_15[196]}
   );
   gpc1_1 gpc986 (
      {stage0_15[437]},
      {stage1_15[197]}
   );
   gpc1_1 gpc987 (
      {stage0_15[438]},
      {stage1_15[198]}
   );
   gpc1_1 gpc988 (
      {stage0_15[439]},
      {stage1_15[199]}
   );
   gpc1_1 gpc989 (
      {stage0_15[440]},
      {stage1_15[200]}
   );
   gpc1_1 gpc990 (
      {stage0_15[441]},
      {stage1_15[201]}
   );
   gpc1_1 gpc991 (
      {stage0_15[442]},
      {stage1_15[202]}
   );
   gpc1_1 gpc992 (
      {stage0_15[443]},
      {stage1_15[203]}
   );
   gpc1_1 gpc993 (
      {stage0_15[444]},
      {stage1_15[204]}
   );
   gpc1_1 gpc994 (
      {stage0_15[445]},
      {stage1_15[205]}
   );
   gpc1_1 gpc995 (
      {stage0_15[446]},
      {stage1_15[206]}
   );
   gpc1_1 gpc996 (
      {stage0_15[447]},
      {stage1_15[207]}
   );
   gpc1_1 gpc997 (
      {stage0_15[448]},
      {stage1_15[208]}
   );
   gpc1_1 gpc998 (
      {stage0_15[449]},
      {stage1_15[209]}
   );
   gpc1_1 gpc999 (
      {stage0_15[450]},
      {stage1_15[210]}
   );
   gpc1_1 gpc1000 (
      {stage0_15[451]},
      {stage1_15[211]}
   );
   gpc1_1 gpc1001 (
      {stage0_15[452]},
      {stage1_15[212]}
   );
   gpc1_1 gpc1002 (
      {stage0_15[453]},
      {stage1_15[213]}
   );
   gpc1_1 gpc1003 (
      {stage0_15[454]},
      {stage1_15[214]}
   );
   gpc1_1 gpc1004 (
      {stage0_15[455]},
      {stage1_15[215]}
   );
   gpc1_1 gpc1005 (
      {stage0_15[456]},
      {stage1_15[216]}
   );
   gpc1_1 gpc1006 (
      {stage0_15[457]},
      {stage1_15[217]}
   );
   gpc1_1 gpc1007 (
      {stage0_15[458]},
      {stage1_15[218]}
   );
   gpc1_1 gpc1008 (
      {stage0_15[459]},
      {stage1_15[219]}
   );
   gpc1_1 gpc1009 (
      {stage0_15[460]},
      {stage1_15[220]}
   );
   gpc1_1 gpc1010 (
      {stage0_15[461]},
      {stage1_15[221]}
   );
   gpc1_1 gpc1011 (
      {stage0_15[462]},
      {stage1_15[222]}
   );
   gpc1_1 gpc1012 (
      {stage0_15[463]},
      {stage1_15[223]}
   );
   gpc1_1 gpc1013 (
      {stage0_15[464]},
      {stage1_15[224]}
   );
   gpc1_1 gpc1014 (
      {stage0_15[465]},
      {stage1_15[225]}
   );
   gpc1_1 gpc1015 (
      {stage0_15[466]},
      {stage1_15[226]}
   );
   gpc1_1 gpc1016 (
      {stage0_15[467]},
      {stage1_15[227]}
   );
   gpc1_1 gpc1017 (
      {stage0_15[468]},
      {stage1_15[228]}
   );
   gpc1_1 gpc1018 (
      {stage0_15[469]},
      {stage1_15[229]}
   );
   gpc1_1 gpc1019 (
      {stage0_15[470]},
      {stage1_15[230]}
   );
   gpc1_1 gpc1020 (
      {stage0_15[471]},
      {stage1_15[231]}
   );
   gpc1_1 gpc1021 (
      {stage0_15[472]},
      {stage1_15[232]}
   );
   gpc1_1 gpc1022 (
      {stage0_15[473]},
      {stage1_15[233]}
   );
   gpc1_1 gpc1023 (
      {stage0_15[474]},
      {stage1_15[234]}
   );
   gpc1_1 gpc1024 (
      {stage0_15[475]},
      {stage1_15[235]}
   );
   gpc1_1 gpc1025 (
      {stage0_15[476]},
      {stage1_15[236]}
   );
   gpc1_1 gpc1026 (
      {stage0_15[477]},
      {stage1_15[237]}
   );
   gpc1_1 gpc1027 (
      {stage0_15[478]},
      {stage1_15[238]}
   );
   gpc1_1 gpc1028 (
      {stage0_15[479]},
      {stage1_15[239]}
   );
   gpc1_1 gpc1029 (
      {stage0_15[480]},
      {stage1_15[240]}
   );
   gpc1_1 gpc1030 (
      {stage0_15[481]},
      {stage1_15[241]}
   );
   gpc1_1 gpc1031 (
      {stage0_15[482]},
      {stage1_15[242]}
   );
   gpc1_1 gpc1032 (
      {stage0_15[483]},
      {stage1_15[243]}
   );
   gpc1_1 gpc1033 (
      {stage0_15[484]},
      {stage1_15[244]}
   );
   gpc1_1 gpc1034 (
      {stage0_15[485]},
      {stage1_15[245]}
   );
   gpc1_1 gpc1035 (
      {stage0_15[486]},
      {stage1_15[246]}
   );
   gpc1_1 gpc1036 (
      {stage0_15[487]},
      {stage1_15[247]}
   );
   gpc1_1 gpc1037 (
      {stage0_15[488]},
      {stage1_15[248]}
   );
   gpc1_1 gpc1038 (
      {stage0_15[489]},
      {stage1_15[249]}
   );
   gpc1_1 gpc1039 (
      {stage0_15[490]},
      {stage1_15[250]}
   );
   gpc1_1 gpc1040 (
      {stage0_15[491]},
      {stage1_15[251]}
   );
   gpc1_1 gpc1041 (
      {stage0_15[492]},
      {stage1_15[252]}
   );
   gpc1_1 gpc1042 (
      {stage0_15[493]},
      {stage1_15[253]}
   );
   gpc1_1 gpc1043 (
      {stage0_15[494]},
      {stage1_15[254]}
   );
   gpc1_1 gpc1044 (
      {stage0_15[495]},
      {stage1_15[255]}
   );
   gpc1_1 gpc1045 (
      {stage0_15[496]},
      {stage1_15[256]}
   );
   gpc1_1 gpc1046 (
      {stage0_15[497]},
      {stage1_15[257]}
   );
   gpc1_1 gpc1047 (
      {stage0_15[498]},
      {stage1_15[258]}
   );
   gpc1_1 gpc1048 (
      {stage0_15[499]},
      {stage1_15[259]}
   );
   gpc1_1 gpc1049 (
      {stage0_15[500]},
      {stage1_15[260]}
   );
   gpc1_1 gpc1050 (
      {stage0_15[501]},
      {stage1_15[261]}
   );
   gpc1_1 gpc1051 (
      {stage0_15[502]},
      {stage1_15[262]}
   );
   gpc1_1 gpc1052 (
      {stage0_15[503]},
      {stage1_15[263]}
   );
   gpc1_1 gpc1053 (
      {stage0_15[504]},
      {stage1_15[264]}
   );
   gpc1_1 gpc1054 (
      {stage0_15[505]},
      {stage1_15[265]}
   );
   gpc1_1 gpc1055 (
      {stage0_15[506]},
      {stage1_15[266]}
   );
   gpc1_1 gpc1056 (
      {stage0_15[507]},
      {stage1_15[267]}
   );
   gpc1_1 gpc1057 (
      {stage0_15[508]},
      {stage1_15[268]}
   );
   gpc1_1 gpc1058 (
      {stage0_15[509]},
      {stage1_15[269]}
   );
   gpc1_1 gpc1059 (
      {stage0_15[510]},
      {stage1_15[270]}
   );
   gpc1_1 gpc1060 (
      {stage0_15[511]},
      {stage1_15[271]}
   );
   gpc1163_5 gpc1061 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc1163_5 gpc1062 (
      {stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_2[1]},
      {stage1_3[1]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc1163_5 gpc1063 (
      {stage1_0[6], stage1_0[7], stage1_0[8]},
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_2[2]},
      {stage1_3[2]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc1163_5 gpc1064 (
      {stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_2[3]},
      {stage1_3[3]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc1163_5 gpc1065 (
      {stage1_0[12], stage1_0[13], stage1_0[14]},
      {stage1_1[24], stage1_1[25], stage1_1[26], stage1_1[27], stage1_1[28], stage1_1[29]},
      {stage1_2[4]},
      {stage1_3[4]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc1163_5 gpc1066 (
      {stage1_0[15], stage1_0[16], stage1_0[17]},
      {stage1_1[30], stage1_1[31], stage1_1[32], stage1_1[33], stage1_1[34], stage1_1[35]},
      {stage1_2[5]},
      {stage1_3[5]},
      {stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5],stage2_0[5]}
   );
   gpc1163_5 gpc1067 (
      {stage1_0[18], stage1_0[19], stage1_0[20]},
      {stage1_1[36], stage1_1[37], stage1_1[38], stage1_1[39], stage1_1[40], stage1_1[41]},
      {stage1_2[6]},
      {stage1_3[6]},
      {stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6],stage2_0[6]}
   );
   gpc1163_5 gpc1068 (
      {stage1_0[21], stage1_0[22], stage1_0[23]},
      {stage1_1[42], stage1_1[43], stage1_1[44], stage1_1[45], stage1_1[46], stage1_1[47]},
      {stage1_2[7]},
      {stage1_3[7]},
      {stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7],stage2_0[7]}
   );
   gpc1163_5 gpc1069 (
      {stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[48], stage1_1[49], stage1_1[50], stage1_1[51], stage1_1[52], stage1_1[53]},
      {stage1_2[8]},
      {stage1_3[8]},
      {stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8],stage2_0[8]}
   );
   gpc1163_5 gpc1070 (
      {stage1_0[27], stage1_0[28], stage1_0[29]},
      {stage1_1[54], stage1_1[55], stage1_1[56], stage1_1[57], stage1_1[58], stage1_1[59]},
      {stage1_2[9]},
      {stage1_3[9]},
      {stage2_4[9],stage2_3[9],stage2_2[9],stage2_1[9],stage2_0[9]}
   );
   gpc1163_5 gpc1071 (
      {stage1_0[30], stage1_0[31], stage1_0[32]},
      {stage1_1[60], stage1_1[61], stage1_1[62], stage1_1[63], stage1_1[64], stage1_1[65]},
      {stage1_2[10]},
      {stage1_3[10]},
      {stage2_4[10],stage2_3[10],stage2_2[10],stage2_1[10],stage2_0[10]}
   );
   gpc1163_5 gpc1072 (
      {stage1_0[33], stage1_0[34], stage1_0[35]},
      {stage1_1[66], stage1_1[67], stage1_1[68], stage1_1[69], stage1_1[70], stage1_1[71]},
      {stage1_2[11]},
      {stage1_3[11]},
      {stage2_4[11],stage2_3[11],stage2_2[11],stage2_1[11],stage2_0[11]}
   );
   gpc606_5 gpc1073 (
      {stage1_0[36], stage1_0[37], stage1_0[38], stage1_0[39], stage1_0[40], stage1_0[41]},
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage2_4[12],stage2_3[12],stage2_2[12],stage2_1[12],stage2_0[12]}
   );
   gpc606_5 gpc1074 (
      {stage1_0[42], stage1_0[43], stage1_0[44], stage1_0[45], stage1_0[46], stage1_0[47]},
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage2_4[13],stage2_3[13],stage2_2[13],stage2_1[13],stage2_0[13]}
   );
   gpc606_5 gpc1075 (
      {stage1_0[48], stage1_0[49], stage1_0[50], stage1_0[51], stage1_0[52], stage1_0[53]},
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage2_4[14],stage2_3[14],stage2_2[14],stage2_1[14],stage2_0[14]}
   );
   gpc606_5 gpc1076 (
      {stage1_0[54], stage1_0[55], stage1_0[56], stage1_0[57], stage1_0[58], stage1_0[59]},
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34], stage1_2[35]},
      {stage2_4[15],stage2_3[15],stage2_2[15],stage2_1[15],stage2_0[15]}
   );
   gpc606_5 gpc1077 (
      {stage1_0[60], stage1_0[61], stage1_0[62], stage1_0[63], stage1_0[64], stage1_0[65]},
      {stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41]},
      {stage2_4[16],stage2_3[16],stage2_2[16],stage2_1[16],stage2_0[16]}
   );
   gpc606_5 gpc1078 (
      {stage1_0[66], stage1_0[67], stage1_0[68], stage1_0[69], stage1_0[70], stage1_0[71]},
      {stage1_2[42], stage1_2[43], stage1_2[44], stage1_2[45], stage1_2[46], stage1_2[47]},
      {stage2_4[17],stage2_3[17],stage2_2[17],stage2_1[17],stage2_0[17]}
   );
   gpc606_5 gpc1079 (
      {stage1_0[72], stage1_0[73], stage1_0[74], stage1_0[75], stage1_0[76], stage1_0[77]},
      {stage1_2[48], stage1_2[49], stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53]},
      {stage2_4[18],stage2_3[18],stage2_2[18],stage2_1[18],stage2_0[18]}
   );
   gpc606_5 gpc1080 (
      {stage1_0[78], stage1_0[79], stage1_0[80], stage1_0[81], stage1_0[82], stage1_0[83]},
      {stage1_2[54], stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59]},
      {stage2_4[19],stage2_3[19],stage2_2[19],stage2_1[19],stage2_0[19]}
   );
   gpc606_5 gpc1081 (
      {stage1_0[84], stage1_0[85], stage1_0[86], stage1_0[87], stage1_0[88], stage1_0[89]},
      {stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63], stage1_2[64], stage1_2[65]},
      {stage2_4[20],stage2_3[20],stage2_2[20],stage2_1[20],stage2_0[20]}
   );
   gpc606_5 gpc1082 (
      {stage1_0[90], stage1_0[91], stage1_0[92], stage1_0[93], stage1_0[94], stage1_0[95]},
      {stage1_2[66], stage1_2[67], stage1_2[68], stage1_2[69], stage1_2[70], stage1_2[71]},
      {stage2_4[21],stage2_3[21],stage2_2[21],stage2_1[21],stage2_0[21]}
   );
   gpc615_5 gpc1083 (
      {stage1_0[96], stage1_0[97], stage1_0[98], stage1_0[99], stage1_0[100]},
      {stage1_1[72]},
      {stage1_2[72], stage1_2[73], stage1_2[74], stage1_2[75], stage1_2[76], stage1_2[77]},
      {stage2_4[22],stage2_3[22],stage2_2[22],stage2_1[22],stage2_0[22]}
   );
   gpc606_5 gpc1084 (
      {stage1_1[73], stage1_1[74], stage1_1[75], stage1_1[76], stage1_1[77], stage1_1[78]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[0],stage2_4[23],stage2_3[23],stage2_2[23],stage2_1[23]}
   );
   gpc606_5 gpc1085 (
      {stage1_1[79], stage1_1[80], stage1_1[81], stage1_1[82], stage1_1[83], stage1_1[84]},
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage2_5[1],stage2_4[24],stage2_3[24],stage2_2[24],stage2_1[24]}
   );
   gpc606_5 gpc1086 (
      {stage1_1[85], stage1_1[86], stage1_1[87], stage1_1[88], stage1_1[89], stage1_1[90]},
      {stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27], stage1_3[28], stage1_3[29]},
      {stage2_5[2],stage2_4[25],stage2_3[25],stage2_2[25],stage2_1[25]}
   );
   gpc606_5 gpc1087 (
      {stage1_1[91], stage1_1[92], stage1_1[93], stage1_1[94], stage1_1[95], stage1_1[96]},
      {stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35]},
      {stage2_5[3],stage2_4[26],stage2_3[26],stage2_2[26],stage2_1[26]}
   );
   gpc606_5 gpc1088 (
      {stage1_1[97], stage1_1[98], stage1_1[99], stage1_1[100], stage1_1[101], stage1_1[102]},
      {stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40], stage1_3[41]},
      {stage2_5[4],stage2_4[27],stage2_3[27],stage2_2[27],stage2_1[27]}
   );
   gpc606_5 gpc1089 (
      {stage1_1[103], stage1_1[104], stage1_1[105], stage1_1[106], stage1_1[107], stage1_1[108]},
      {stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45], stage1_3[46], stage1_3[47]},
      {stage2_5[5],stage2_4[28],stage2_3[28],stage2_2[28],stage2_1[28]}
   );
   gpc606_5 gpc1090 (
      {stage1_1[109], stage1_1[110], stage1_1[111], stage1_1[112], stage1_1[113], stage1_1[114]},
      {stage1_3[48], stage1_3[49], stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53]},
      {stage2_5[6],stage2_4[29],stage2_3[29],stage2_2[29],stage2_1[29]}
   );
   gpc606_5 gpc1091 (
      {stage1_1[115], stage1_1[116], stage1_1[117], stage1_1[118], stage1_1[119], stage1_1[120]},
      {stage1_3[54], stage1_3[55], stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59]},
      {stage2_5[7],stage2_4[30],stage2_3[30],stage2_2[30],stage2_1[30]}
   );
   gpc606_5 gpc1092 (
      {stage1_1[121], stage1_1[122], stage1_1[123], stage1_1[124], stage1_1[125], stage1_1[126]},
      {stage1_3[60], stage1_3[61], stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65]},
      {stage2_5[8],stage2_4[31],stage2_3[31],stage2_2[31],stage2_1[31]}
   );
   gpc606_5 gpc1093 (
      {stage1_1[127], stage1_1[128], stage1_1[129], stage1_1[130], stage1_1[131], stage1_1[132]},
      {stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70], stage1_3[71]},
      {stage2_5[9],stage2_4[32],stage2_3[32],stage2_2[32],stage2_1[32]}
   );
   gpc606_5 gpc1094 (
      {stage1_1[133], stage1_1[134], stage1_1[135], stage1_1[136], stage1_1[137], stage1_1[138]},
      {stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75], stage1_3[76], stage1_3[77]},
      {stage2_5[10],stage2_4[33],stage2_3[33],stage2_2[33],stage2_1[33]}
   );
   gpc606_5 gpc1095 (
      {stage1_1[139], stage1_1[140], stage1_1[141], stage1_1[142], stage1_1[143], stage1_1[144]},
      {stage1_3[78], stage1_3[79], stage1_3[80], stage1_3[81], stage1_3[82], stage1_3[83]},
      {stage2_5[11],stage2_4[34],stage2_3[34],stage2_2[34],stage2_1[34]}
   );
   gpc606_5 gpc1096 (
      {stage1_1[145], stage1_1[146], stage1_1[147], stage1_1[148], stage1_1[149], stage1_1[150]},
      {stage1_3[84], stage1_3[85], stage1_3[86], stage1_3[87], stage1_3[88], stage1_3[89]},
      {stage2_5[12],stage2_4[35],stage2_3[35],stage2_2[35],stage2_1[35]}
   );
   gpc606_5 gpc1097 (
      {stage1_1[151], stage1_1[152], stage1_1[153], stage1_1[154], stage1_1[155], stage1_1[156]},
      {stage1_3[90], stage1_3[91], stage1_3[92], stage1_3[93], stage1_3[94], stage1_3[95]},
      {stage2_5[13],stage2_4[36],stage2_3[36],stage2_2[36],stage2_1[36]}
   );
   gpc606_5 gpc1098 (
      {stage1_1[157], stage1_1[158], stage1_1[159], stage1_1[160], stage1_1[161], stage1_1[162]},
      {stage1_3[96], stage1_3[97], stage1_3[98], stage1_3[99], stage1_3[100], stage1_3[101]},
      {stage2_5[14],stage2_4[37],stage2_3[37],stage2_2[37],stage2_1[37]}
   );
   gpc606_5 gpc1099 (
      {stage1_1[163], stage1_1[164], stage1_1[165], stage1_1[166], stage1_1[167], stage1_1[168]},
      {stage1_3[102], stage1_3[103], stage1_3[104], stage1_3[105], stage1_3[106], stage1_3[107]},
      {stage2_5[15],stage2_4[38],stage2_3[38],stage2_2[38],stage2_1[38]}
   );
   gpc606_5 gpc1100 (
      {stage1_1[169], stage1_1[170], stage1_1[171], stage1_1[172], stage1_1[173], stage1_1[174]},
      {stage1_3[108], stage1_3[109], stage1_3[110], stage1_3[111], stage1_3[112], stage1_3[113]},
      {stage2_5[16],stage2_4[39],stage2_3[39],stage2_2[39],stage2_1[39]}
   );
   gpc606_5 gpc1101 (
      {stage1_1[175], stage1_1[176], stage1_1[177], stage1_1[178], stage1_1[179], 1'b0},
      {stage1_3[114], stage1_3[115], stage1_3[116], stage1_3[117], stage1_3[118], stage1_3[119]},
      {stage2_5[17],stage2_4[40],stage2_3[40],stage2_2[40],stage2_1[40]}
   );
   gpc615_5 gpc1102 (
      {stage1_2[78], stage1_2[79], stage1_2[80], stage1_2[81], stage1_2[82]},
      {stage1_3[120]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[18],stage2_4[41],stage2_3[41],stage2_2[41]}
   );
   gpc615_5 gpc1103 (
      {stage1_2[83], stage1_2[84], stage1_2[85], stage1_2[86], stage1_2[87]},
      {stage1_3[121]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[19],stage2_4[42],stage2_3[42],stage2_2[42]}
   );
   gpc615_5 gpc1104 (
      {stage1_2[88], stage1_2[89], stage1_2[90], stage1_2[91], stage1_2[92]},
      {stage1_3[122]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[20],stage2_4[43],stage2_3[43],stage2_2[43]}
   );
   gpc615_5 gpc1105 (
      {stage1_2[93], stage1_2[94], stage1_2[95], stage1_2[96], stage1_2[97]},
      {stage1_3[123]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[21],stage2_4[44],stage2_3[44],stage2_2[44]}
   );
   gpc615_5 gpc1106 (
      {stage1_2[98], stage1_2[99], stage1_2[100], stage1_2[101], stage1_2[102]},
      {stage1_3[124]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[22],stage2_4[45],stage2_3[45],stage2_2[45]}
   );
   gpc615_5 gpc1107 (
      {stage1_2[103], stage1_2[104], stage1_2[105], stage1_2[106], stage1_2[107]},
      {stage1_3[125]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[23],stage2_4[46],stage2_3[46],stage2_2[46]}
   );
   gpc615_5 gpc1108 (
      {stage1_2[108], stage1_2[109], stage1_2[110], stage1_2[111], stage1_2[112]},
      {stage1_3[126]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[24],stage2_4[47],stage2_3[47],stage2_2[47]}
   );
   gpc615_5 gpc1109 (
      {stage1_2[113], stage1_2[114], stage1_2[115], stage1_2[116], stage1_2[117]},
      {stage1_3[127]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[25],stage2_4[48],stage2_3[48],stage2_2[48]}
   );
   gpc615_5 gpc1110 (
      {stage1_2[118], stage1_2[119], stage1_2[120], stage1_2[121], stage1_2[122]},
      {stage1_3[128]},
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53]},
      {stage2_6[8],stage2_5[26],stage2_4[49],stage2_3[49],stage2_2[49]}
   );
   gpc615_5 gpc1111 (
      {stage1_2[123], stage1_2[124], stage1_2[125], stage1_2[126], stage1_2[127]},
      {stage1_3[129]},
      {stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57], stage1_4[58], stage1_4[59]},
      {stage2_6[9],stage2_5[27],stage2_4[50],stage2_3[50],stage2_2[50]}
   );
   gpc615_5 gpc1112 (
      {stage1_2[128], stage1_2[129], stage1_2[130], stage1_2[131], stage1_2[132]},
      {stage1_3[130]},
      {stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63], stage1_4[64], stage1_4[65]},
      {stage2_6[10],stage2_5[28],stage2_4[51],stage2_3[51],stage2_2[51]}
   );
   gpc615_5 gpc1113 (
      {stage1_2[133], stage1_2[134], stage1_2[135], stage1_2[136], stage1_2[137]},
      {stage1_3[131]},
      {stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69], stage1_4[70], stage1_4[71]},
      {stage2_6[11],stage2_5[29],stage2_4[52],stage2_3[52],stage2_2[52]}
   );
   gpc615_5 gpc1114 (
      {stage1_2[138], stage1_2[139], stage1_2[140], stage1_2[141], stage1_2[142]},
      {stage1_3[132]},
      {stage1_4[72], stage1_4[73], stage1_4[74], stage1_4[75], stage1_4[76], stage1_4[77]},
      {stage2_6[12],stage2_5[30],stage2_4[53],stage2_3[53],stage2_2[53]}
   );
   gpc615_5 gpc1115 (
      {stage1_2[143], stage1_2[144], stage1_2[145], stage1_2[146], stage1_2[147]},
      {stage1_3[133]},
      {stage1_4[78], stage1_4[79], stage1_4[80], stage1_4[81], stage1_4[82], stage1_4[83]},
      {stage2_6[13],stage2_5[31],stage2_4[54],stage2_3[54],stage2_2[54]}
   );
   gpc615_5 gpc1116 (
      {stage1_2[148], stage1_2[149], stage1_2[150], stage1_2[151], stage1_2[152]},
      {stage1_3[134]},
      {stage1_4[84], stage1_4[85], stage1_4[86], stage1_4[87], stage1_4[88], stage1_4[89]},
      {stage2_6[14],stage2_5[32],stage2_4[55],stage2_3[55],stage2_2[55]}
   );
   gpc615_5 gpc1117 (
      {stage1_2[153], stage1_2[154], stage1_2[155], stage1_2[156], stage1_2[157]},
      {stage1_3[135]},
      {stage1_4[90], stage1_4[91], stage1_4[92], stage1_4[93], stage1_4[94], stage1_4[95]},
      {stage2_6[15],stage2_5[33],stage2_4[56],stage2_3[56],stage2_2[56]}
   );
   gpc615_5 gpc1118 (
      {stage1_2[158], stage1_2[159], stage1_2[160], stage1_2[161], stage1_2[162]},
      {stage1_3[136]},
      {stage1_4[96], stage1_4[97], stage1_4[98], stage1_4[99], stage1_4[100], stage1_4[101]},
      {stage2_6[16],stage2_5[34],stage2_4[57],stage2_3[57],stage2_2[57]}
   );
   gpc615_5 gpc1119 (
      {stage1_2[163], stage1_2[164], stage1_2[165], stage1_2[166], stage1_2[167]},
      {stage1_3[137]},
      {stage1_4[102], stage1_4[103], stage1_4[104], stage1_4[105], stage1_4[106], stage1_4[107]},
      {stage2_6[17],stage2_5[35],stage2_4[58],stage2_3[58],stage2_2[58]}
   );
   gpc615_5 gpc1120 (
      {stage1_2[168], stage1_2[169], stage1_2[170], stage1_2[171], stage1_2[172]},
      {stage1_3[138]},
      {stage1_4[108], stage1_4[109], stage1_4[110], stage1_4[111], stage1_4[112], stage1_4[113]},
      {stage2_6[18],stage2_5[36],stage2_4[59],stage2_3[59],stage2_2[59]}
   );
   gpc615_5 gpc1121 (
      {stage1_3[139], stage1_3[140], stage1_3[141], stage1_3[142], stage1_3[143]},
      {stage1_4[114]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[19],stage2_5[37],stage2_4[60],stage2_3[60]}
   );
   gpc615_5 gpc1122 (
      {stage1_3[144], stage1_3[145], stage1_3[146], stage1_3[147], stage1_3[148]},
      {stage1_4[115]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[20],stage2_5[38],stage2_4[61],stage2_3[61]}
   );
   gpc615_5 gpc1123 (
      {stage1_3[149], stage1_3[150], stage1_3[151], stage1_3[152], stage1_3[153]},
      {stage1_4[116]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[21],stage2_5[39],stage2_4[62],stage2_3[62]}
   );
   gpc615_5 gpc1124 (
      {stage1_3[154], stage1_3[155], stage1_3[156], stage1_3[157], stage1_3[158]},
      {stage1_4[117]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[22],stage2_5[40],stage2_4[63],stage2_3[63]}
   );
   gpc615_5 gpc1125 (
      {stage1_3[159], stage1_3[160], stage1_3[161], stage1_3[162], stage1_3[163]},
      {stage1_4[118]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[23],stage2_5[41],stage2_4[64],stage2_3[64]}
   );
   gpc615_5 gpc1126 (
      {stage1_3[164], stage1_3[165], stage1_3[166], stage1_3[167], stage1_3[168]},
      {stage1_4[119]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[24],stage2_5[42],stage2_4[65],stage2_3[65]}
   );
   gpc615_5 gpc1127 (
      {stage1_3[169], stage1_3[170], stage1_3[171], stage1_3[172], stage1_3[173]},
      {stage1_4[120]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[25],stage2_5[43],stage2_4[66],stage2_3[66]}
   );
   gpc615_5 gpc1128 (
      {stage1_3[174], stage1_3[175], stage1_3[176], stage1_3[177], stage1_3[178]},
      {stage1_4[121]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[26],stage2_5[44],stage2_4[67],stage2_3[67]}
   );
   gpc615_5 gpc1129 (
      {stage1_3[179], stage1_3[180], stage1_3[181], stage1_3[182], stage1_3[183]},
      {stage1_4[122]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[27],stage2_5[45],stage2_4[68],stage2_3[68]}
   );
   gpc615_5 gpc1130 (
      {stage1_3[184], stage1_3[185], stage1_3[186], stage1_3[187], stage1_3[188]},
      {stage1_4[123]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[28],stage2_5[46],stage2_4[69],stage2_3[69]}
   );
   gpc615_5 gpc1131 (
      {stage1_3[189], stage1_3[190], stage1_3[191], stage1_3[192], stage1_3[193]},
      {stage1_4[124]},
      {stage1_5[60], stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65]},
      {stage2_7[10],stage2_6[29],stage2_5[47],stage2_4[70],stage2_3[70]}
   );
   gpc615_5 gpc1132 (
      {stage1_3[194], stage1_3[195], stage1_3[196], stage1_3[197], stage1_3[198]},
      {stage1_4[125]},
      {stage1_5[66], stage1_5[67], stage1_5[68], stage1_5[69], stage1_5[70], stage1_5[71]},
      {stage2_7[11],stage2_6[30],stage2_5[48],stage2_4[71],stage2_3[71]}
   );
   gpc615_5 gpc1133 (
      {stage1_3[199], stage1_3[200], stage1_3[201], stage1_3[202], stage1_3[203]},
      {stage1_4[126]},
      {stage1_5[72], stage1_5[73], stage1_5[74], stage1_5[75], stage1_5[76], stage1_5[77]},
      {stage2_7[12],stage2_6[31],stage2_5[49],stage2_4[72],stage2_3[72]}
   );
   gpc615_5 gpc1134 (
      {stage1_3[204], stage1_3[205], stage1_3[206], stage1_3[207], stage1_3[208]},
      {stage1_4[127]},
      {stage1_5[78], stage1_5[79], stage1_5[80], stage1_5[81], stage1_5[82], stage1_5[83]},
      {stage2_7[13],stage2_6[32],stage2_5[50],stage2_4[73],stage2_3[73]}
   );
   gpc615_5 gpc1135 (
      {stage1_3[209], stage1_3[210], stage1_3[211], stage1_3[212], stage1_3[213]},
      {stage1_4[128]},
      {stage1_5[84], stage1_5[85], stage1_5[86], stage1_5[87], stage1_5[88], stage1_5[89]},
      {stage2_7[14],stage2_6[33],stage2_5[51],stage2_4[74],stage2_3[74]}
   );
   gpc615_5 gpc1136 (
      {stage1_3[214], stage1_3[215], stage1_3[216], stage1_3[217], stage1_3[218]},
      {stage1_4[129]},
      {stage1_5[90], stage1_5[91], stage1_5[92], stage1_5[93], stage1_5[94], stage1_5[95]},
      {stage2_7[15],stage2_6[34],stage2_5[52],stage2_4[75],stage2_3[75]}
   );
   gpc606_5 gpc1137 (
      {stage1_4[130], stage1_4[131], stage1_4[132], stage1_4[133], stage1_4[134], stage1_4[135]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[16],stage2_6[35],stage2_5[53],stage2_4[76]}
   );
   gpc606_5 gpc1138 (
      {stage1_4[136], stage1_4[137], stage1_4[138], stage1_4[139], stage1_4[140], stage1_4[141]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[17],stage2_6[36],stage2_5[54],stage2_4[77]}
   );
   gpc606_5 gpc1139 (
      {stage1_4[142], stage1_4[143], stage1_4[144], stage1_4[145], stage1_4[146], stage1_4[147]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[18],stage2_6[37],stage2_5[55],stage2_4[78]}
   );
   gpc606_5 gpc1140 (
      {stage1_4[148], stage1_4[149], stage1_4[150], stage1_4[151], stage1_4[152], stage1_4[153]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[19],stage2_6[38],stage2_5[56],stage2_4[79]}
   );
   gpc606_5 gpc1141 (
      {stage1_4[154], stage1_4[155], stage1_4[156], stage1_4[157], stage1_4[158], stage1_4[159]},
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage2_8[4],stage2_7[20],stage2_6[39],stage2_5[57],stage2_4[80]}
   );
   gpc606_5 gpc1142 (
      {stage1_4[160], stage1_4[161], stage1_4[162], stage1_4[163], stage1_4[164], stage1_4[165]},
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage2_8[5],stage2_7[21],stage2_6[40],stage2_5[58],stage2_4[81]}
   );
   gpc606_5 gpc1143 (
      {stage1_4[166], stage1_4[167], stage1_4[168], stage1_4[169], stage1_4[170], stage1_4[171]},
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage2_8[6],stage2_7[22],stage2_6[41],stage2_5[59],stage2_4[82]}
   );
   gpc606_5 gpc1144 (
      {stage1_4[172], stage1_4[173], stage1_4[174], stage1_4[175], stage1_4[176], stage1_4[177]},
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage2_8[7],stage2_7[23],stage2_6[42],stage2_5[60],stage2_4[83]}
   );
   gpc606_5 gpc1145 (
      {stage1_4[178], stage1_4[179], stage1_4[180], stage1_4[181], stage1_4[182], stage1_4[183]},
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53]},
      {stage2_8[8],stage2_7[24],stage2_6[43],stage2_5[61],stage2_4[84]}
   );
   gpc606_5 gpc1146 (
      {stage1_4[184], stage1_4[185], stage1_4[186], stage1_4[187], stage1_4[188], stage1_4[189]},
      {stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage2_8[9],stage2_7[25],stage2_6[44],stage2_5[62],stage2_4[85]}
   );
   gpc606_5 gpc1147 (
      {stage1_4[190], stage1_4[191], stage1_4[192], stage1_4[193], stage1_4[194], stage1_4[195]},
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64], stage1_6[65]},
      {stage2_8[10],stage2_7[26],stage2_6[45],stage2_5[63],stage2_4[86]}
   );
   gpc606_5 gpc1148 (
      {stage1_4[196], stage1_4[197], stage1_4[198], stage1_4[199], stage1_4[200], stage1_4[201]},
      {stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69], stage1_6[70], stage1_6[71]},
      {stage2_8[11],stage2_7[27],stage2_6[46],stage2_5[64],stage2_4[87]}
   );
   gpc606_5 gpc1149 (
      {stage1_4[202], stage1_4[203], stage1_4[204], stage1_4[205], stage1_4[206], stage1_4[207]},
      {stage1_6[72], stage1_6[73], stage1_6[74], stage1_6[75], stage1_6[76], stage1_6[77]},
      {stage2_8[12],stage2_7[28],stage2_6[47],stage2_5[65],stage2_4[88]}
   );
   gpc606_5 gpc1150 (
      {stage1_4[208], stage1_4[209], stage1_4[210], stage1_4[211], stage1_4[212], stage1_4[213]},
      {stage1_6[78], stage1_6[79], stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83]},
      {stage2_8[13],stage2_7[29],stage2_6[48],stage2_5[66],stage2_4[89]}
   );
   gpc606_5 gpc1151 (
      {stage1_5[96], stage1_5[97], stage1_5[98], stage1_5[99], stage1_5[100], stage1_5[101]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[14],stage2_7[30],stage2_6[49],stage2_5[67]}
   );
   gpc606_5 gpc1152 (
      {stage1_5[102], stage1_5[103], stage1_5[104], stage1_5[105], stage1_5[106], stage1_5[107]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[15],stage2_7[31],stage2_6[50],stage2_5[68]}
   );
   gpc606_5 gpc1153 (
      {stage1_5[108], stage1_5[109], stage1_5[110], stage1_5[111], stage1_5[112], stage1_5[113]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[16],stage2_7[32],stage2_6[51],stage2_5[69]}
   );
   gpc606_5 gpc1154 (
      {stage1_5[114], stage1_5[115], stage1_5[116], stage1_5[117], stage1_5[118], stage1_5[119]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[17],stage2_7[33],stage2_6[52],stage2_5[70]}
   );
   gpc606_5 gpc1155 (
      {stage1_5[120], stage1_5[121], stage1_5[122], stage1_5[123], stage1_5[124], stage1_5[125]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[18],stage2_7[34],stage2_6[53],stage2_5[71]}
   );
   gpc606_5 gpc1156 (
      {stage1_5[126], stage1_5[127], stage1_5[128], stage1_5[129], stage1_5[130], stage1_5[131]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[19],stage2_7[35],stage2_6[54],stage2_5[72]}
   );
   gpc606_5 gpc1157 (
      {stage1_5[132], stage1_5[133], stage1_5[134], stage1_5[135], stage1_5[136], stage1_5[137]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[20],stage2_7[36],stage2_6[55],stage2_5[73]}
   );
   gpc606_5 gpc1158 (
      {stage1_5[138], stage1_5[139], stage1_5[140], stage1_5[141], stage1_5[142], stage1_5[143]},
      {stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage2_9[7],stage2_8[21],stage2_7[37],stage2_6[56],stage2_5[74]}
   );
   gpc606_5 gpc1159 (
      {stage1_5[144], stage1_5[145], stage1_5[146], stage1_5[147], stage1_5[148], stage1_5[149]},
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52], stage1_7[53]},
      {stage2_9[8],stage2_8[22],stage2_7[38],stage2_6[57],stage2_5[75]}
   );
   gpc606_5 gpc1160 (
      {stage1_5[150], stage1_5[151], stage1_5[152], stage1_5[153], stage1_5[154], stage1_5[155]},
      {stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58], stage1_7[59]},
      {stage2_9[9],stage2_8[23],stage2_7[39],stage2_6[58],stage2_5[76]}
   );
   gpc606_5 gpc1161 (
      {stage1_5[156], stage1_5[157], stage1_5[158], stage1_5[159], stage1_5[160], stage1_5[161]},
      {stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63], stage1_7[64], stage1_7[65]},
      {stage2_9[10],stage2_8[24],stage2_7[40],stage2_6[59],stage2_5[77]}
   );
   gpc606_5 gpc1162 (
      {stage1_5[162], stage1_5[163], stage1_5[164], stage1_5[165], stage1_5[166], stage1_5[167]},
      {stage1_7[66], stage1_7[67], stage1_7[68], stage1_7[69], stage1_7[70], stage1_7[71]},
      {stage2_9[11],stage2_8[25],stage2_7[41],stage2_6[60],stage2_5[78]}
   );
   gpc606_5 gpc1163 (
      {stage1_5[168], stage1_5[169], stage1_5[170], stage1_5[171], stage1_5[172], stage1_5[173]},
      {stage1_7[72], stage1_7[73], stage1_7[74], stage1_7[75], stage1_7[76], stage1_7[77]},
      {stage2_9[12],stage2_8[26],stage2_7[42],stage2_6[61],stage2_5[79]}
   );
   gpc606_5 gpc1164 (
      {stage1_5[174], stage1_5[175], stage1_5[176], stage1_5[177], stage1_5[178], stage1_5[179]},
      {stage1_7[78], stage1_7[79], stage1_7[80], stage1_7[81], stage1_7[82], stage1_7[83]},
      {stage2_9[13],stage2_8[27],stage2_7[43],stage2_6[62],stage2_5[80]}
   );
   gpc606_5 gpc1165 (
      {stage1_5[180], stage1_5[181], stage1_5[182], stage1_5[183], stage1_5[184], stage1_5[185]},
      {stage1_7[84], stage1_7[85], stage1_7[86], stage1_7[87], stage1_7[88], stage1_7[89]},
      {stage2_9[14],stage2_8[28],stage2_7[44],stage2_6[63],stage2_5[81]}
   );
   gpc606_5 gpc1166 (
      {stage1_5[186], stage1_5[187], stage1_5[188], stage1_5[189], stage1_5[190], stage1_5[191]},
      {stage1_7[90], stage1_7[91], stage1_7[92], stage1_7[93], stage1_7[94], stage1_7[95]},
      {stage2_9[15],stage2_8[29],stage2_7[45],stage2_6[64],stage2_5[82]}
   );
   gpc606_5 gpc1167 (
      {stage1_5[192], stage1_5[193], stage1_5[194], stage1_5[195], stage1_5[196], stage1_5[197]},
      {stage1_7[96], stage1_7[97], stage1_7[98], stage1_7[99], stage1_7[100], stage1_7[101]},
      {stage2_9[16],stage2_8[30],stage2_7[46],stage2_6[65],stage2_5[83]}
   );
   gpc606_5 gpc1168 (
      {stage1_5[198], stage1_5[199], stage1_5[200], stage1_5[201], stage1_5[202], stage1_5[203]},
      {stage1_7[102], stage1_7[103], stage1_7[104], stage1_7[105], stage1_7[106], stage1_7[107]},
      {stage2_9[17],stage2_8[31],stage2_7[47],stage2_6[66],stage2_5[84]}
   );
   gpc606_5 gpc1169 (
      {stage1_5[204], stage1_5[205], stage1_5[206], stage1_5[207], stage1_5[208], stage1_5[209]},
      {stage1_7[108], stage1_7[109], stage1_7[110], stage1_7[111], stage1_7[112], stage1_7[113]},
      {stage2_9[18],stage2_8[32],stage2_7[48],stage2_6[67],stage2_5[85]}
   );
   gpc606_5 gpc1170 (
      {stage1_6[84], stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], stage1_6[89]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[19],stage2_8[33],stage2_7[49],stage2_6[68]}
   );
   gpc606_5 gpc1171 (
      {stage1_6[90], stage1_6[91], stage1_6[92], stage1_6[93], stage1_6[94], stage1_6[95]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[20],stage2_8[34],stage2_7[50],stage2_6[69]}
   );
   gpc606_5 gpc1172 (
      {stage1_6[96], stage1_6[97], stage1_6[98], stage1_6[99], stage1_6[100], stage1_6[101]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[21],stage2_8[35],stage2_7[51],stage2_6[70]}
   );
   gpc606_5 gpc1173 (
      {stage1_6[102], stage1_6[103], stage1_6[104], stage1_6[105], stage1_6[106], stage1_6[107]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[22],stage2_8[36],stage2_7[52],stage2_6[71]}
   );
   gpc606_5 gpc1174 (
      {stage1_6[108], stage1_6[109], stage1_6[110], stage1_6[111], stage1_6[112], stage1_6[113]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[23],stage2_8[37],stage2_7[53],stage2_6[72]}
   );
   gpc606_5 gpc1175 (
      {stage1_6[114], stage1_6[115], stage1_6[116], stage1_6[117], stage1_6[118], stage1_6[119]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[24],stage2_8[38],stage2_7[54],stage2_6[73]}
   );
   gpc606_5 gpc1176 (
      {stage1_6[120], stage1_6[121], stage1_6[122], stage1_6[123], stage1_6[124], stage1_6[125]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[25],stage2_8[39],stage2_7[55],stage2_6[74]}
   );
   gpc606_5 gpc1177 (
      {stage1_6[126], stage1_6[127], stage1_6[128], stage1_6[129], stage1_6[130], stage1_6[131]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[26],stage2_8[40],stage2_7[56],stage2_6[75]}
   );
   gpc606_5 gpc1178 (
      {stage1_6[132], stage1_6[133], stage1_6[134], stage1_6[135], stage1_6[136], stage1_6[137]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[27],stage2_8[41],stage2_7[57],stage2_6[76]}
   );
   gpc606_5 gpc1179 (
      {stage1_6[138], stage1_6[139], stage1_6[140], stage1_6[141], stage1_6[142], stage1_6[143]},
      {stage1_8[54], stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59]},
      {stage2_10[9],stage2_9[28],stage2_8[42],stage2_7[58],stage2_6[77]}
   );
   gpc606_5 gpc1180 (
      {stage1_6[144], stage1_6[145], stage1_6[146], stage1_6[147], stage1_6[148], stage1_6[149]},
      {stage1_8[60], stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65]},
      {stage2_10[10],stage2_9[29],stage2_8[43],stage2_7[59],stage2_6[78]}
   );
   gpc606_5 gpc1181 (
      {stage1_6[150], stage1_6[151], stage1_6[152], stage1_6[153], stage1_6[154], stage1_6[155]},
      {stage1_8[66], stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71]},
      {stage2_10[11],stage2_9[30],stage2_8[44],stage2_7[60],stage2_6[79]}
   );
   gpc606_5 gpc1182 (
      {stage1_6[156], stage1_6[157], stage1_6[158], stage1_6[159], stage1_6[160], stage1_6[161]},
      {stage1_8[72], stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77]},
      {stage2_10[12],stage2_9[31],stage2_8[45],stage2_7[61],stage2_6[80]}
   );
   gpc606_5 gpc1183 (
      {stage1_6[162], stage1_6[163], stage1_6[164], stage1_6[165], stage1_6[166], stage1_6[167]},
      {stage1_8[78], stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83]},
      {stage2_10[13],stage2_9[32],stage2_8[46],stage2_7[62],stage2_6[81]}
   );
   gpc606_5 gpc1184 (
      {stage1_6[168], stage1_6[169], stage1_6[170], stage1_6[171], stage1_6[172], stage1_6[173]},
      {stage1_8[84], stage1_8[85], stage1_8[86], stage1_8[87], stage1_8[88], stage1_8[89]},
      {stage2_10[14],stage2_9[33],stage2_8[47],stage2_7[63],stage2_6[82]}
   );
   gpc615_5 gpc1185 (
      {stage1_6[174], stage1_6[175], stage1_6[176], stage1_6[177], stage1_6[178]},
      {stage1_7[114]},
      {stage1_8[90], stage1_8[91], stage1_8[92], stage1_8[93], stage1_8[94], stage1_8[95]},
      {stage2_10[15],stage2_9[34],stage2_8[48],stage2_7[64],stage2_6[83]}
   );
   gpc615_5 gpc1186 (
      {stage1_6[179], stage1_6[180], stage1_6[181], stage1_6[182], stage1_6[183]},
      {stage1_7[115]},
      {stage1_8[96], stage1_8[97], stage1_8[98], stage1_8[99], stage1_8[100], stage1_8[101]},
      {stage2_10[16],stage2_9[35],stage2_8[49],stage2_7[65],stage2_6[84]}
   );
   gpc615_5 gpc1187 (
      {stage1_6[184], stage1_6[185], stage1_6[186], stage1_6[187], stage1_6[188]},
      {stage1_7[116]},
      {stage1_8[102], stage1_8[103], stage1_8[104], stage1_8[105], stage1_8[106], stage1_8[107]},
      {stage2_10[17],stage2_9[36],stage2_8[50],stage2_7[66],stage2_6[85]}
   );
   gpc615_5 gpc1188 (
      {stage1_7[117], stage1_7[118], stage1_7[119], stage1_7[120], stage1_7[121]},
      {stage1_8[108]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[18],stage2_9[37],stage2_8[51],stage2_7[67]}
   );
   gpc615_5 gpc1189 (
      {stage1_7[122], stage1_7[123], stage1_7[124], stage1_7[125], stage1_7[126]},
      {stage1_8[109]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[19],stage2_9[38],stage2_8[52],stage2_7[68]}
   );
   gpc615_5 gpc1190 (
      {stage1_7[127], stage1_7[128], stage1_7[129], stage1_7[130], stage1_7[131]},
      {stage1_8[110]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[20],stage2_9[39],stage2_8[53],stage2_7[69]}
   );
   gpc615_5 gpc1191 (
      {stage1_7[132], stage1_7[133], stage1_7[134], stage1_7[135], stage1_7[136]},
      {stage1_8[111]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[21],stage2_9[40],stage2_8[54],stage2_7[70]}
   );
   gpc615_5 gpc1192 (
      {stage1_7[137], stage1_7[138], stage1_7[139], stage1_7[140], stage1_7[141]},
      {stage1_8[112]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[22],stage2_9[41],stage2_8[55],stage2_7[71]}
   );
   gpc615_5 gpc1193 (
      {stage1_7[142], stage1_7[143], stage1_7[144], stage1_7[145], stage1_7[146]},
      {stage1_8[113]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[23],stage2_9[42],stage2_8[56],stage2_7[72]}
   );
   gpc615_5 gpc1194 (
      {stage1_7[147], stage1_7[148], stage1_7[149], stage1_7[150], stage1_7[151]},
      {stage1_8[114]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[24],stage2_9[43],stage2_8[57],stage2_7[73]}
   );
   gpc615_5 gpc1195 (
      {stage1_7[152], stage1_7[153], stage1_7[154], stage1_7[155], stage1_7[156]},
      {stage1_8[115]},
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage2_11[7],stage2_10[25],stage2_9[44],stage2_8[58],stage2_7[74]}
   );
   gpc615_5 gpc1196 (
      {stage1_7[157], stage1_7[158], stage1_7[159], stage1_7[160], stage1_7[161]},
      {stage1_8[116]},
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage2_11[8],stage2_10[26],stage2_9[45],stage2_8[59],stage2_7[75]}
   );
   gpc615_5 gpc1197 (
      {stage1_7[162], stage1_7[163], stage1_7[164], stage1_7[165], stage1_7[166]},
      {stage1_8[117]},
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage2_11[9],stage2_10[27],stage2_9[46],stage2_8[60],stage2_7[76]}
   );
   gpc615_5 gpc1198 (
      {stage1_7[167], stage1_7[168], stage1_7[169], stage1_7[170], stage1_7[171]},
      {stage1_8[118]},
      {stage1_9[60], stage1_9[61], stage1_9[62], stage1_9[63], stage1_9[64], stage1_9[65]},
      {stage2_11[10],stage2_10[28],stage2_9[47],stage2_8[61],stage2_7[77]}
   );
   gpc615_5 gpc1199 (
      {stage1_7[172], stage1_7[173], stage1_7[174], stage1_7[175], stage1_7[176]},
      {stage1_8[119]},
      {stage1_9[66], stage1_9[67], stage1_9[68], stage1_9[69], stage1_9[70], stage1_9[71]},
      {stage2_11[11],stage2_10[29],stage2_9[48],stage2_8[62],stage2_7[78]}
   );
   gpc615_5 gpc1200 (
      {stage1_7[177], stage1_7[178], stage1_7[179], stage1_7[180], stage1_7[181]},
      {stage1_8[120]},
      {stage1_9[72], stage1_9[73], stage1_9[74], stage1_9[75], stage1_9[76], stage1_9[77]},
      {stage2_11[12],stage2_10[30],stage2_9[49],stage2_8[63],stage2_7[79]}
   );
   gpc615_5 gpc1201 (
      {stage1_7[182], stage1_7[183], stage1_7[184], stage1_7[185], stage1_7[186]},
      {stage1_8[121]},
      {stage1_9[78], stage1_9[79], stage1_9[80], stage1_9[81], stage1_9[82], stage1_9[83]},
      {stage2_11[13],stage2_10[31],stage2_9[50],stage2_8[64],stage2_7[80]}
   );
   gpc615_5 gpc1202 (
      {stage1_7[187], stage1_7[188], stage1_7[189], stage1_7[190], stage1_7[191]},
      {stage1_8[122]},
      {stage1_9[84], stage1_9[85], stage1_9[86], stage1_9[87], stage1_9[88], stage1_9[89]},
      {stage2_11[14],stage2_10[32],stage2_9[51],stage2_8[65],stage2_7[81]}
   );
   gpc615_5 gpc1203 (
      {stage1_7[192], stage1_7[193], stage1_7[194], stage1_7[195], stage1_7[196]},
      {stage1_8[123]},
      {stage1_9[90], stage1_9[91], stage1_9[92], stage1_9[93], stage1_9[94], stage1_9[95]},
      {stage2_11[15],stage2_10[33],stage2_9[52],stage2_8[66],stage2_7[82]}
   );
   gpc615_5 gpc1204 (
      {stage1_7[197], stage1_7[198], stage1_7[199], stage1_7[200], stage1_7[201]},
      {stage1_8[124]},
      {stage1_9[96], stage1_9[97], stage1_9[98], stage1_9[99], stage1_9[100], stage1_9[101]},
      {stage2_11[16],stage2_10[34],stage2_9[53],stage2_8[67],stage2_7[83]}
   );
   gpc615_5 gpc1205 (
      {stage1_7[202], stage1_7[203], stage1_7[204], stage1_7[205], stage1_7[206]},
      {stage1_8[125]},
      {stage1_9[102], stage1_9[103], stage1_9[104], stage1_9[105], stage1_9[106], stage1_9[107]},
      {stage2_11[17],stage2_10[35],stage2_9[54],stage2_8[68],stage2_7[84]}
   );
   gpc606_5 gpc1206 (
      {stage1_8[126], stage1_8[127], stage1_8[128], stage1_8[129], stage1_8[130], stage1_8[131]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[18],stage2_10[36],stage2_9[55],stage2_8[69]}
   );
   gpc606_5 gpc1207 (
      {stage1_8[132], stage1_8[133], stage1_8[134], stage1_8[135], stage1_8[136], stage1_8[137]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[19],stage2_10[37],stage2_9[56],stage2_8[70]}
   );
   gpc615_5 gpc1208 (
      {stage1_8[138], stage1_8[139], stage1_8[140], stage1_8[141], stage1_8[142]},
      {stage1_9[108]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[20],stage2_10[38],stage2_9[57],stage2_8[71]}
   );
   gpc615_5 gpc1209 (
      {stage1_8[143], stage1_8[144], stage1_8[145], stage1_8[146], stage1_8[147]},
      {stage1_9[109]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[21],stage2_10[39],stage2_9[58],stage2_8[72]}
   );
   gpc615_5 gpc1210 (
      {stage1_8[148], stage1_8[149], stage1_8[150], stage1_8[151], stage1_8[152]},
      {stage1_9[110]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[22],stage2_10[40],stage2_9[59],stage2_8[73]}
   );
   gpc615_5 gpc1211 (
      {stage1_8[153], stage1_8[154], stage1_8[155], stage1_8[156], stage1_8[157]},
      {stage1_9[111]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[23],stage2_10[41],stage2_9[60],stage2_8[74]}
   );
   gpc615_5 gpc1212 (
      {stage1_8[158], stage1_8[159], stage1_8[160], stage1_8[161], stage1_8[162]},
      {stage1_9[112]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[24],stage2_10[42],stage2_9[61],stage2_8[75]}
   );
   gpc615_5 gpc1213 (
      {stage1_8[163], stage1_8[164], stage1_8[165], stage1_8[166], stage1_8[167]},
      {stage1_9[113]},
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage2_12[7],stage2_11[25],stage2_10[43],stage2_9[62],stage2_8[76]}
   );
   gpc615_5 gpc1214 (
      {stage1_8[168], stage1_8[169], stage1_8[170], stage1_8[171], stage1_8[172]},
      {stage1_9[114]},
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage2_12[8],stage2_11[26],stage2_10[44],stage2_9[63],stage2_8[77]}
   );
   gpc615_5 gpc1215 (
      {stage1_8[173], stage1_8[174], stage1_8[175], stage1_8[176], stage1_8[177]},
      {stage1_9[115]},
      {stage1_10[54], stage1_10[55], stage1_10[56], stage1_10[57], stage1_10[58], stage1_10[59]},
      {stage2_12[9],stage2_11[27],stage2_10[45],stage2_9[64],stage2_8[78]}
   );
   gpc615_5 gpc1216 (
      {stage1_8[178], stage1_8[179], stage1_8[180], stage1_8[181], stage1_8[182]},
      {stage1_9[116]},
      {stage1_10[60], stage1_10[61], stage1_10[62], stage1_10[63], stage1_10[64], stage1_10[65]},
      {stage2_12[10],stage2_11[28],stage2_10[46],stage2_9[65],stage2_8[79]}
   );
   gpc615_5 gpc1217 (
      {stage1_8[183], stage1_8[184], stage1_8[185], stage1_8[186], stage1_8[187]},
      {stage1_9[117]},
      {stage1_10[66], stage1_10[67], stage1_10[68], stage1_10[69], stage1_10[70], stage1_10[71]},
      {stage2_12[11],stage2_11[29],stage2_10[47],stage2_9[66],stage2_8[80]}
   );
   gpc615_5 gpc1218 (
      {stage1_8[188], stage1_8[189], stage1_8[190], stage1_8[191], stage1_8[192]},
      {stage1_9[118]},
      {stage1_10[72], stage1_10[73], stage1_10[74], stage1_10[75], stage1_10[76], stage1_10[77]},
      {stage2_12[12],stage2_11[30],stage2_10[48],stage2_9[67],stage2_8[81]}
   );
   gpc615_5 gpc1219 (
      {stage1_8[193], stage1_8[194], stage1_8[195], stage1_8[196], stage1_8[197]},
      {stage1_9[119]},
      {stage1_10[78], stage1_10[79], stage1_10[80], stage1_10[81], stage1_10[82], stage1_10[83]},
      {stage2_12[13],stage2_11[31],stage2_10[49],stage2_9[68],stage2_8[82]}
   );
   gpc615_5 gpc1220 (
      {stage1_8[198], stage1_8[199], stage1_8[200], stage1_8[201], stage1_8[202]},
      {stage1_9[120]},
      {stage1_10[84], stage1_10[85], stage1_10[86], stage1_10[87], stage1_10[88], stage1_10[89]},
      {stage2_12[14],stage2_11[32],stage2_10[50],stage2_9[69],stage2_8[83]}
   );
   gpc615_5 gpc1221 (
      {stage1_8[203], stage1_8[204], stage1_8[205], stage1_8[206], stage1_8[207]},
      {stage1_9[121]},
      {stage1_10[90], stage1_10[91], stage1_10[92], stage1_10[93], stage1_10[94], stage1_10[95]},
      {stage2_12[15],stage2_11[33],stage2_10[51],stage2_9[70],stage2_8[84]}
   );
   gpc615_5 gpc1222 (
      {stage1_8[208], stage1_8[209], stage1_8[210], stage1_8[211], stage1_8[212]},
      {stage1_9[122]},
      {stage1_10[96], stage1_10[97], stage1_10[98], stage1_10[99], stage1_10[100], stage1_10[101]},
      {stage2_12[16],stage2_11[34],stage2_10[52],stage2_9[71],stage2_8[85]}
   );
   gpc615_5 gpc1223 (
      {stage1_8[213], stage1_8[214], stage1_8[215], stage1_8[216], stage1_8[217]},
      {stage1_9[123]},
      {stage1_10[102], stage1_10[103], stage1_10[104], stage1_10[105], stage1_10[106], stage1_10[107]},
      {stage2_12[17],stage2_11[35],stage2_10[53],stage2_9[72],stage2_8[86]}
   );
   gpc606_5 gpc1224 (
      {stage1_9[124], stage1_9[125], stage1_9[126], stage1_9[127], stage1_9[128], stage1_9[129]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[18],stage2_11[36],stage2_10[54],stage2_9[73]}
   );
   gpc606_5 gpc1225 (
      {stage1_9[130], stage1_9[131], stage1_9[132], stage1_9[133], stage1_9[134], stage1_9[135]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[19],stage2_11[37],stage2_10[55],stage2_9[74]}
   );
   gpc606_5 gpc1226 (
      {stage1_9[136], stage1_9[137], stage1_9[138], stage1_9[139], stage1_9[140], stage1_9[141]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[20],stage2_11[38],stage2_10[56],stage2_9[75]}
   );
   gpc606_5 gpc1227 (
      {stage1_9[142], stage1_9[143], stage1_9[144], stage1_9[145], stage1_9[146], stage1_9[147]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[21],stage2_11[39],stage2_10[57],stage2_9[76]}
   );
   gpc606_5 gpc1228 (
      {stage1_9[148], stage1_9[149], stage1_9[150], stage1_9[151], stage1_9[152], stage1_9[153]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[22],stage2_11[40],stage2_10[58],stage2_9[77]}
   );
   gpc606_5 gpc1229 (
      {stage1_9[154], stage1_9[155], stage1_9[156], stage1_9[157], stage1_9[158], stage1_9[159]},
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35]},
      {stage2_13[5],stage2_12[23],stage2_11[41],stage2_10[59],stage2_9[78]}
   );
   gpc606_5 gpc1230 (
      {stage1_9[160], stage1_9[161], stage1_9[162], stage1_9[163], stage1_9[164], stage1_9[165]},
      {stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41]},
      {stage2_13[6],stage2_12[24],stage2_11[42],stage2_10[60],stage2_9[79]}
   );
   gpc606_5 gpc1231 (
      {stage1_9[166], stage1_9[167], stage1_9[168], stage1_9[169], stage1_9[170], stage1_9[171]},
      {stage1_11[42], stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47]},
      {stage2_13[7],stage2_12[25],stage2_11[43],stage2_10[61],stage2_9[80]}
   );
   gpc606_5 gpc1232 (
      {stage1_9[172], stage1_9[173], stage1_9[174], stage1_9[175], stage1_9[176], stage1_9[177]},
      {stage1_11[48], stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage2_13[8],stage2_12[26],stage2_11[44],stage2_10[62],stage2_9[81]}
   );
   gpc606_5 gpc1233 (
      {stage1_9[178], stage1_9[179], stage1_9[180], stage1_9[181], stage1_9[182], stage1_9[183]},
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58], stage1_11[59]},
      {stage2_13[9],stage2_12[27],stage2_11[45],stage2_10[63],stage2_9[82]}
   );
   gpc606_5 gpc1234 (
      {stage1_9[184], stage1_9[185], stage1_9[186], stage1_9[187], stage1_9[188], stage1_9[189]},
      {stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63], stage1_11[64], stage1_11[65]},
      {stage2_13[10],stage2_12[28],stage2_11[46],stage2_10[64],stage2_9[83]}
   );
   gpc606_5 gpc1235 (
      {stage1_9[190], stage1_9[191], stage1_9[192], stage1_9[193], stage1_9[194], stage1_9[195]},
      {stage1_11[66], stage1_11[67], stage1_11[68], stage1_11[69], stage1_11[70], stage1_11[71]},
      {stage2_13[11],stage2_12[29],stage2_11[47],stage2_10[65],stage2_9[84]}
   );
   gpc606_5 gpc1236 (
      {stage1_9[196], stage1_9[197], stage1_9[198], stage1_9[199], stage1_9[200], stage1_9[201]},
      {stage1_11[72], stage1_11[73], stage1_11[74], stage1_11[75], stage1_11[76], stage1_11[77]},
      {stage2_13[12],stage2_12[30],stage2_11[48],stage2_10[66],stage2_9[85]}
   );
   gpc606_5 gpc1237 (
      {stage1_9[202], stage1_9[203], stage1_9[204], stage1_9[205], stage1_9[206], stage1_9[207]},
      {stage1_11[78], stage1_11[79], stage1_11[80], stage1_11[81], stage1_11[82], stage1_11[83]},
      {stage2_13[13],stage2_12[31],stage2_11[49],stage2_10[67],stage2_9[86]}
   );
   gpc606_5 gpc1238 (
      {stage1_9[208], stage1_9[209], stage1_9[210], stage1_9[211], stage1_9[212], stage1_9[213]},
      {stage1_11[84], stage1_11[85], stage1_11[86], stage1_11[87], stage1_11[88], stage1_11[89]},
      {stage2_13[14],stage2_12[32],stage2_11[50],stage2_10[68],stage2_9[87]}
   );
   gpc606_5 gpc1239 (
      {stage1_10[108], stage1_10[109], stage1_10[110], stage1_10[111], stage1_10[112], stage1_10[113]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[15],stage2_12[33],stage2_11[51],stage2_10[69]}
   );
   gpc606_5 gpc1240 (
      {stage1_10[114], stage1_10[115], stage1_10[116], stage1_10[117], stage1_10[118], stage1_10[119]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[16],stage2_12[34],stage2_11[52],stage2_10[70]}
   );
   gpc606_5 gpc1241 (
      {stage1_10[120], stage1_10[121], stage1_10[122], stage1_10[123], stage1_10[124], stage1_10[125]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[17],stage2_12[35],stage2_11[53],stage2_10[71]}
   );
   gpc606_5 gpc1242 (
      {stage1_10[126], stage1_10[127], stage1_10[128], stage1_10[129], stage1_10[130], stage1_10[131]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[18],stage2_12[36],stage2_11[54],stage2_10[72]}
   );
   gpc606_5 gpc1243 (
      {stage1_10[132], stage1_10[133], stage1_10[134], stage1_10[135], stage1_10[136], stage1_10[137]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[19],stage2_12[37],stage2_11[55],stage2_10[73]}
   );
   gpc606_5 gpc1244 (
      {stage1_10[138], stage1_10[139], stage1_10[140], stage1_10[141], stage1_10[142], stage1_10[143]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[20],stage2_12[38],stage2_11[56],stage2_10[74]}
   );
   gpc606_5 gpc1245 (
      {stage1_10[144], stage1_10[145], stage1_10[146], stage1_10[147], stage1_10[148], stage1_10[149]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[21],stage2_12[39],stage2_11[57],stage2_10[75]}
   );
   gpc606_5 gpc1246 (
      {stage1_10[150], stage1_10[151], stage1_10[152], stage1_10[153], stage1_10[154], stage1_10[155]},
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage2_14[7],stage2_13[22],stage2_12[40],stage2_11[58],stage2_10[76]}
   );
   gpc606_5 gpc1247 (
      {stage1_10[156], stage1_10[157], stage1_10[158], stage1_10[159], stage1_10[160], stage1_10[161]},
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage2_14[8],stage2_13[23],stage2_12[41],stage2_11[59],stage2_10[77]}
   );
   gpc606_5 gpc1248 (
      {stage1_10[162], stage1_10[163], stage1_10[164], stage1_10[165], stage1_10[166], stage1_10[167]},
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage2_14[9],stage2_13[24],stage2_12[42],stage2_11[60],stage2_10[78]}
   );
   gpc606_5 gpc1249 (
      {stage1_10[168], stage1_10[169], stage1_10[170], stage1_10[171], stage1_10[172], stage1_10[173]},
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage2_14[10],stage2_13[25],stage2_12[43],stage2_11[61],stage2_10[79]}
   );
   gpc606_5 gpc1250 (
      {stage1_10[174], stage1_10[175], stage1_10[176], stage1_10[177], stage1_10[178], stage1_10[179]},
      {stage1_12[66], stage1_12[67], stage1_12[68], stage1_12[69], stage1_12[70], stage1_12[71]},
      {stage2_14[11],stage2_13[26],stage2_12[44],stage2_11[62],stage2_10[80]}
   );
   gpc606_5 gpc1251 (
      {stage1_10[180], stage1_10[181], stage1_10[182], stage1_10[183], stage1_10[184], stage1_10[185]},
      {stage1_12[72], stage1_12[73], stage1_12[74], stage1_12[75], stage1_12[76], stage1_12[77]},
      {stage2_14[12],stage2_13[27],stage2_12[45],stage2_11[63],stage2_10[81]}
   );
   gpc606_5 gpc1252 (
      {stage1_10[186], stage1_10[187], stage1_10[188], stage1_10[189], stage1_10[190], stage1_10[191]},
      {stage1_12[78], stage1_12[79], stage1_12[80], stage1_12[81], stage1_12[82], stage1_12[83]},
      {stage2_14[13],stage2_13[28],stage2_12[46],stage2_11[64],stage2_10[82]}
   );
   gpc606_5 gpc1253 (
      {stage1_10[192], stage1_10[193], stage1_10[194], stage1_10[195], stage1_10[196], stage1_10[197]},
      {stage1_12[84], stage1_12[85], stage1_12[86], stage1_12[87], stage1_12[88], stage1_12[89]},
      {stage2_14[14],stage2_13[29],stage2_12[47],stage2_11[65],stage2_10[83]}
   );
   gpc606_5 gpc1254 (
      {stage1_10[198], stage1_10[199], stage1_10[200], stage1_10[201], stage1_10[202], stage1_10[203]},
      {stage1_12[90], stage1_12[91], stage1_12[92], stage1_12[93], stage1_12[94], stage1_12[95]},
      {stage2_14[15],stage2_13[30],stage2_12[48],stage2_11[66],stage2_10[84]}
   );
   gpc606_5 gpc1255 (
      {stage1_10[204], stage1_10[205], stage1_10[206], stage1_10[207], stage1_10[208], stage1_10[209]},
      {stage1_12[96], stage1_12[97], stage1_12[98], stage1_12[99], stage1_12[100], stage1_12[101]},
      {stage2_14[16],stage2_13[31],stage2_12[49],stage2_11[67],stage2_10[85]}
   );
   gpc615_5 gpc1256 (
      {stage1_11[90], stage1_11[91], stage1_11[92], stage1_11[93], stage1_11[94]},
      {stage1_12[102]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[17],stage2_13[32],stage2_12[50],stage2_11[68]}
   );
   gpc615_5 gpc1257 (
      {stage1_11[95], stage1_11[96], stage1_11[97], stage1_11[98], stage1_11[99]},
      {stage1_12[103]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[18],stage2_13[33],stage2_12[51],stage2_11[69]}
   );
   gpc615_5 gpc1258 (
      {stage1_11[100], stage1_11[101], stage1_11[102], stage1_11[103], stage1_11[104]},
      {stage1_12[104]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[19],stage2_13[34],stage2_12[52],stage2_11[70]}
   );
   gpc615_5 gpc1259 (
      {stage1_11[105], stage1_11[106], stage1_11[107], stage1_11[108], stage1_11[109]},
      {stage1_12[105]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[20],stage2_13[35],stage2_12[53],stage2_11[71]}
   );
   gpc615_5 gpc1260 (
      {stage1_11[110], stage1_11[111], stage1_11[112], stage1_11[113], stage1_11[114]},
      {stage1_12[106]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[21],stage2_13[36],stage2_12[54],stage2_11[72]}
   );
   gpc615_5 gpc1261 (
      {stage1_11[115], stage1_11[116], stage1_11[117], stage1_11[118], stage1_11[119]},
      {stage1_12[107]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[22],stage2_13[37],stage2_12[55],stage2_11[73]}
   );
   gpc606_5 gpc1262 (
      {stage1_12[108], stage1_12[109], stage1_12[110], stage1_12[111], stage1_12[112], stage1_12[113]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[6],stage2_14[23],stage2_13[38],stage2_12[56]}
   );
   gpc606_5 gpc1263 (
      {stage1_12[114], stage1_12[115], stage1_12[116], stage1_12[117], stage1_12[118], stage1_12[119]},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[7],stage2_14[24],stage2_13[39],stage2_12[57]}
   );
   gpc606_5 gpc1264 (
      {stage1_12[120], stage1_12[121], stage1_12[122], stage1_12[123], stage1_12[124], stage1_12[125]},
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage2_16[2],stage2_15[8],stage2_14[25],stage2_13[40],stage2_12[58]}
   );
   gpc606_5 gpc1265 (
      {stage1_12[126], stage1_12[127], stage1_12[128], stage1_12[129], stage1_12[130], stage1_12[131]},
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23]},
      {stage2_16[3],stage2_15[9],stage2_14[26],stage2_13[41],stage2_12[59]}
   );
   gpc606_5 gpc1266 (
      {stage1_12[132], stage1_12[133], stage1_12[134], stage1_12[135], stage1_12[136], stage1_12[137]},
      {stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29]},
      {stage2_16[4],stage2_15[10],stage2_14[27],stage2_13[42],stage2_12[60]}
   );
   gpc606_5 gpc1267 (
      {stage1_12[138], stage1_12[139], stage1_12[140], stage1_12[141], stage1_12[142], stage1_12[143]},
      {stage1_14[30], stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35]},
      {stage2_16[5],stage2_15[11],stage2_14[28],stage2_13[43],stage2_12[61]}
   );
   gpc606_5 gpc1268 (
      {stage1_12[144], stage1_12[145], stage1_12[146], stage1_12[147], stage1_12[148], stage1_12[149]},
      {stage1_14[36], stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage2_16[6],stage2_15[12],stage2_14[29],stage2_13[44],stage2_12[62]}
   );
   gpc606_5 gpc1269 (
      {stage1_12[150], stage1_12[151], stage1_12[152], stage1_12[153], stage1_12[154], stage1_12[155]},
      {stage1_14[42], stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage2_16[7],stage2_15[13],stage2_14[30],stage2_13[45],stage2_12[63]}
   );
   gpc606_5 gpc1270 (
      {stage1_12[156], stage1_12[157], stage1_12[158], stage1_12[159], stage1_12[160], stage1_12[161]},
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53]},
      {stage2_16[8],stage2_15[14],stage2_14[31],stage2_13[46],stage2_12[64]}
   );
   gpc606_5 gpc1271 (
      {stage1_12[162], stage1_12[163], stage1_12[164], stage1_12[165], stage1_12[166], stage1_12[167]},
      {stage1_14[54], stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59]},
      {stage2_16[9],stage2_15[15],stage2_14[32],stage2_13[47],stage2_12[65]}
   );
   gpc606_5 gpc1272 (
      {stage1_12[168], stage1_12[169], stage1_12[170], stage1_12[171], stage1_12[172], stage1_12[173]},
      {stage1_14[60], stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65]},
      {stage2_16[10],stage2_15[16],stage2_14[33],stage2_13[48],stage2_12[66]}
   );
   gpc606_5 gpc1273 (
      {stage1_12[174], stage1_12[175], stage1_12[176], stage1_12[177], stage1_12[178], stage1_12[179]},
      {stage1_14[66], stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71]},
      {stage2_16[11],stage2_15[17],stage2_14[34],stage2_13[49],stage2_12[67]}
   );
   gpc606_5 gpc1274 (
      {stage1_12[180], stage1_12[181], stage1_12[182], stage1_12[183], stage1_12[184], stage1_12[185]},
      {stage1_14[72], stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76], stage1_14[77]},
      {stage2_16[12],stage2_15[18],stage2_14[35],stage2_13[50],stage2_12[68]}
   );
   gpc606_5 gpc1275 (
      {stage1_12[186], stage1_12[187], stage1_12[188], stage1_12[189], stage1_12[190], stage1_12[191]},
      {stage1_14[78], stage1_14[79], stage1_14[80], stage1_14[81], stage1_14[82], stage1_14[83]},
      {stage2_16[13],stage2_15[19],stage2_14[36],stage2_13[51],stage2_12[69]}
   );
   gpc606_5 gpc1276 (
      {stage1_12[192], stage1_12[193], stage1_12[194], stage1_12[195], stage1_12[196], stage1_12[197]},
      {stage1_14[84], stage1_14[85], stage1_14[86], stage1_14[87], stage1_14[88], stage1_14[89]},
      {stage2_16[14],stage2_15[20],stage2_14[37],stage2_13[52],stage2_12[70]}
   );
   gpc606_5 gpc1277 (
      {stage1_12[198], stage1_12[199], stage1_12[200], stage1_12[201], stage1_12[202], stage1_12[203]},
      {stage1_14[90], stage1_14[91], stage1_14[92], stage1_14[93], stage1_14[94], stage1_14[95]},
      {stage2_16[15],stage2_15[21],stage2_14[38],stage2_13[53],stage2_12[71]}
   );
   gpc606_5 gpc1278 (
      {stage1_12[204], stage1_12[205], stage1_12[206], stage1_12[207], stage1_12[208], stage1_12[209]},
      {stage1_14[96], stage1_14[97], stage1_14[98], stage1_14[99], stage1_14[100], stage1_14[101]},
      {stage2_16[16],stage2_15[22],stage2_14[39],stage2_13[54],stage2_12[72]}
   );
   gpc606_5 gpc1279 (
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[17],stage2_15[23],stage2_14[40],stage2_13[55]}
   );
   gpc606_5 gpc1280 (
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[18],stage2_15[24],stage2_14[41],stage2_13[56]}
   );
   gpc606_5 gpc1281 (
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[19],stage2_15[25],stage2_14[42],stage2_13[57]}
   );
   gpc606_5 gpc1282 (
      {stage1_13[54], stage1_13[55], stage1_13[56], stage1_13[57], stage1_13[58], stage1_13[59]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[20],stage2_15[26],stage2_14[43],stage2_13[58]}
   );
   gpc606_5 gpc1283 (
      {stage1_13[60], stage1_13[61], stage1_13[62], stage1_13[63], stage1_13[64], stage1_13[65]},
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage2_17[4],stage2_16[21],stage2_15[27],stage2_14[44],stage2_13[59]}
   );
   gpc606_5 gpc1284 (
      {stage1_13[66], stage1_13[67], stage1_13[68], stage1_13[69], stage1_13[70], stage1_13[71]},
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage2_17[5],stage2_16[22],stage2_15[28],stage2_14[45],stage2_13[60]}
   );
   gpc606_5 gpc1285 (
      {stage1_13[72], stage1_13[73], stage1_13[74], stage1_13[75], stage1_13[76], stage1_13[77]},
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage2_17[6],stage2_16[23],stage2_15[29],stage2_14[46],stage2_13[61]}
   );
   gpc606_5 gpc1286 (
      {stage1_13[78], stage1_13[79], stage1_13[80], stage1_13[81], stage1_13[82], stage1_13[83]},
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46], stage1_15[47]},
      {stage2_17[7],stage2_16[24],stage2_15[30],stage2_14[47],stage2_13[62]}
   );
   gpc606_5 gpc1287 (
      {stage1_13[84], stage1_13[85], stage1_13[86], stage1_13[87], stage1_13[88], stage1_13[89]},
      {stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51], stage1_15[52], stage1_15[53]},
      {stage2_17[8],stage2_16[25],stage2_15[31],stage2_14[48],stage2_13[63]}
   );
   gpc606_5 gpc1288 (
      {stage1_13[90], stage1_13[91], stage1_13[92], stage1_13[93], stage1_13[94], stage1_13[95]},
      {stage1_15[54], stage1_15[55], stage1_15[56], stage1_15[57], stage1_15[58], stage1_15[59]},
      {stage2_17[9],stage2_16[26],stage2_15[32],stage2_14[49],stage2_13[64]}
   );
   gpc606_5 gpc1289 (
      {stage1_13[96], stage1_13[97], stage1_13[98], stage1_13[99], stage1_13[100], stage1_13[101]},
      {stage1_15[60], stage1_15[61], stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65]},
      {stage2_17[10],stage2_16[27],stage2_15[33],stage2_14[50],stage2_13[65]}
   );
   gpc606_5 gpc1290 (
      {stage1_13[102], stage1_13[103], stage1_13[104], stage1_13[105], stage1_13[106], stage1_13[107]},
      {stage1_15[66], stage1_15[67], stage1_15[68], stage1_15[69], stage1_15[70], stage1_15[71]},
      {stage2_17[11],stage2_16[28],stage2_15[34],stage2_14[51],stage2_13[66]}
   );
   gpc606_5 gpc1291 (
      {stage1_13[108], stage1_13[109], stage1_13[110], stage1_13[111], stage1_13[112], stage1_13[113]},
      {stage1_15[72], stage1_15[73], stage1_15[74], stage1_15[75], stage1_15[76], stage1_15[77]},
      {stage2_17[12],stage2_16[29],stage2_15[35],stage2_14[52],stage2_13[67]}
   );
   gpc606_5 gpc1292 (
      {stage1_13[114], stage1_13[115], stage1_13[116], stage1_13[117], stage1_13[118], stage1_13[119]},
      {stage1_15[78], stage1_15[79], stage1_15[80], stage1_15[81], stage1_15[82], stage1_15[83]},
      {stage2_17[13],stage2_16[30],stage2_15[36],stage2_14[53],stage2_13[68]}
   );
   gpc606_5 gpc1293 (
      {stage1_13[120], stage1_13[121], stage1_13[122], stage1_13[123], stage1_13[124], stage1_13[125]},
      {stage1_15[84], stage1_15[85], stage1_15[86], stage1_15[87], stage1_15[88], stage1_15[89]},
      {stage2_17[14],stage2_16[31],stage2_15[37],stage2_14[54],stage2_13[69]}
   );
   gpc606_5 gpc1294 (
      {stage1_13[126], stage1_13[127], stage1_13[128], stage1_13[129], stage1_13[130], stage1_13[131]},
      {stage1_15[90], stage1_15[91], stage1_15[92], stage1_15[93], stage1_15[94], stage1_15[95]},
      {stage2_17[15],stage2_16[32],stage2_15[38],stage2_14[55],stage2_13[70]}
   );
   gpc615_5 gpc1295 (
      {stage1_13[132], stage1_13[133], stage1_13[134], stage1_13[135], stage1_13[136]},
      {stage1_14[102]},
      {stage1_15[96], stage1_15[97], stage1_15[98], stage1_15[99], stage1_15[100], stage1_15[101]},
      {stage2_17[16],stage2_16[33],stage2_15[39],stage2_14[56],stage2_13[71]}
   );
   gpc615_5 gpc1296 (
      {stage1_13[137], stage1_13[138], stage1_13[139], stage1_13[140], stage1_13[141]},
      {stage1_14[103]},
      {stage1_15[102], stage1_15[103], stage1_15[104], stage1_15[105], stage1_15[106], stage1_15[107]},
      {stage2_17[17],stage2_16[34],stage2_15[40],stage2_14[57],stage2_13[72]}
   );
   gpc615_5 gpc1297 (
      {stage1_13[142], stage1_13[143], stage1_13[144], stage1_13[145], stage1_13[146]},
      {stage1_14[104]},
      {stage1_15[108], stage1_15[109], stage1_15[110], stage1_15[111], stage1_15[112], stage1_15[113]},
      {stage2_17[18],stage2_16[35],stage2_15[41],stage2_14[58],stage2_13[73]}
   );
   gpc615_5 gpc1298 (
      {stage1_13[147], stage1_13[148], stage1_13[149], stage1_13[150], stage1_13[151]},
      {stage1_14[105]},
      {stage1_15[114], stage1_15[115], stage1_15[116], stage1_15[117], stage1_15[118], stage1_15[119]},
      {stage2_17[19],stage2_16[36],stage2_15[42],stage2_14[59],stage2_13[74]}
   );
   gpc615_5 gpc1299 (
      {stage1_13[152], stage1_13[153], stage1_13[154], stage1_13[155], stage1_13[156]},
      {stage1_14[106]},
      {stage1_15[120], stage1_15[121], stage1_15[122], stage1_15[123], stage1_15[124], stage1_15[125]},
      {stage2_17[20],stage2_16[37],stage2_15[43],stage2_14[60],stage2_13[75]}
   );
   gpc615_5 gpc1300 (
      {stage1_13[157], stage1_13[158], stage1_13[159], stage1_13[160], stage1_13[161]},
      {stage1_14[107]},
      {stage1_15[126], stage1_15[127], stage1_15[128], stage1_15[129], stage1_15[130], stage1_15[131]},
      {stage2_17[21],stage2_16[38],stage2_15[44],stage2_14[61],stage2_13[76]}
   );
   gpc615_5 gpc1301 (
      {stage1_13[162], stage1_13[163], stage1_13[164], stage1_13[165], stage1_13[166]},
      {stage1_14[108]},
      {stage1_15[132], stage1_15[133], stage1_15[134], stage1_15[135], stage1_15[136], stage1_15[137]},
      {stage2_17[22],stage2_16[39],stage2_15[45],stage2_14[62],stage2_13[77]}
   );
   gpc615_5 gpc1302 (
      {stage1_13[167], stage1_13[168], stage1_13[169], stage1_13[170], stage1_13[171]},
      {stage1_14[109]},
      {stage1_15[138], stage1_15[139], stage1_15[140], stage1_15[141], stage1_15[142], stage1_15[143]},
      {stage2_17[23],stage2_16[40],stage2_15[46],stage2_14[63],stage2_13[78]}
   );
   gpc615_5 gpc1303 (
      {stage1_13[172], stage1_13[173], stage1_13[174], stage1_13[175], stage1_13[176]},
      {stage1_14[110]},
      {stage1_15[144], stage1_15[145], stage1_15[146], stage1_15[147], stage1_15[148], stage1_15[149]},
      {stage2_17[24],stage2_16[41],stage2_15[47],stage2_14[64],stage2_13[79]}
   );
   gpc615_5 gpc1304 (
      {stage1_13[177], stage1_13[178], stage1_13[179], stage1_13[180], stage1_13[181]},
      {stage1_14[111]},
      {stage1_15[150], stage1_15[151], stage1_15[152], stage1_15[153], stage1_15[154], stage1_15[155]},
      {stage2_17[25],stage2_16[42],stage2_15[48],stage2_14[65],stage2_13[80]}
   );
   gpc615_5 gpc1305 (
      {stage1_13[182], stage1_13[183], stage1_13[184], stage1_13[185], stage1_13[186]},
      {stage1_14[112]},
      {stage1_15[156], stage1_15[157], stage1_15[158], stage1_15[159], stage1_15[160], stage1_15[161]},
      {stage2_17[26],stage2_16[43],stage2_15[49],stage2_14[66],stage2_13[81]}
   );
   gpc615_5 gpc1306 (
      {stage1_13[187], stage1_13[188], stage1_13[189], stage1_13[190], stage1_13[191]},
      {stage1_14[113]},
      {stage1_15[162], stage1_15[163], stage1_15[164], stage1_15[165], stage1_15[166], stage1_15[167]},
      {stage2_17[27],stage2_16[44],stage2_15[50],stage2_14[67],stage2_13[82]}
   );
   gpc615_5 gpc1307 (
      {stage1_13[192], stage1_13[193], stage1_13[194], stage1_13[195], stage1_13[196]},
      {stage1_14[114]},
      {stage1_15[168], stage1_15[169], stage1_15[170], stage1_15[171], stage1_15[172], stage1_15[173]},
      {stage2_17[28],stage2_16[45],stage2_15[51],stage2_14[68],stage2_13[83]}
   );
   gpc615_5 gpc1308 (
      {stage1_13[197], stage1_13[198], stage1_13[199], stage1_13[200], stage1_13[201]},
      {stage1_14[115]},
      {stage1_15[174], stage1_15[175], stage1_15[176], stage1_15[177], stage1_15[178], stage1_15[179]},
      {stage2_17[29],stage2_16[46],stage2_15[52],stage2_14[69],stage2_13[84]}
   );
   gpc615_5 gpc1309 (
      {stage1_13[202], stage1_13[203], stage1_13[204], stage1_13[205], stage1_13[206]},
      {stage1_14[116]},
      {stage1_15[180], stage1_15[181], stage1_15[182], stage1_15[183], stage1_15[184], stage1_15[185]},
      {stage2_17[30],stage2_16[47],stage2_15[53],stage2_14[70],stage2_13[85]}
   );
   gpc615_5 gpc1310 (
      {stage1_13[207], stage1_13[208], stage1_13[209], stage1_13[210], stage1_13[211]},
      {stage1_14[117]},
      {stage1_15[186], stage1_15[187], stage1_15[188], stage1_15[189], stage1_15[190], stage1_15[191]},
      {stage2_17[31],stage2_16[48],stage2_15[54],stage2_14[71],stage2_13[86]}
   );
   gpc615_5 gpc1311 (
      {stage1_13[212], stage1_13[213], stage1_13[214], stage1_13[215], stage1_13[216]},
      {stage1_14[118]},
      {stage1_15[192], stage1_15[193], stage1_15[194], stage1_15[195], stage1_15[196], stage1_15[197]},
      {stage2_17[32],stage2_16[49],stage2_15[55],stage2_14[72],stage2_13[87]}
   );
   gpc615_5 gpc1312 (
      {stage1_13[217], stage1_13[218], stage1_13[219], stage1_13[220], stage1_13[221]},
      {stage1_14[119]},
      {stage1_15[198], stage1_15[199], stage1_15[200], stage1_15[201], stage1_15[202], stage1_15[203]},
      {stage2_17[33],stage2_16[50],stage2_15[56],stage2_14[73],stage2_13[88]}
   );
   gpc615_5 gpc1313 (
      {stage1_13[222], stage1_13[223], stage1_13[224], stage1_13[225], stage1_13[226]},
      {stage1_14[120]},
      {stage1_15[204], stage1_15[205], stage1_15[206], stage1_15[207], stage1_15[208], stage1_15[209]},
      {stage2_17[34],stage2_16[51],stage2_15[57],stage2_14[74],stage2_13[89]}
   );
   gpc615_5 gpc1314 (
      {stage1_13[227], stage1_13[228], stage1_13[229], stage1_13[230], stage1_13[231]},
      {stage1_14[121]},
      {stage1_15[210], stage1_15[211], stage1_15[212], stage1_15[213], stage1_15[214], stage1_15[215]},
      {stage2_17[35],stage2_16[52],stage2_15[58],stage2_14[75],stage2_13[90]}
   );
   gpc606_5 gpc1315 (
      {stage1_14[122], stage1_14[123], stage1_14[124], stage1_14[125], stage1_14[126], stage1_14[127]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[36],stage2_16[53],stage2_15[59],stage2_14[76]}
   );
   gpc606_5 gpc1316 (
      {stage1_14[128], stage1_14[129], stage1_14[130], stage1_14[131], stage1_14[132], stage1_14[133]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[37],stage2_16[54],stage2_15[60],stage2_14[77]}
   );
   gpc606_5 gpc1317 (
      {stage1_14[134], stage1_14[135], stage1_14[136], stage1_14[137], stage1_14[138], stage1_14[139]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[38],stage2_16[55],stage2_15[61],stage2_14[78]}
   );
   gpc606_5 gpc1318 (
      {stage1_14[140], stage1_14[141], stage1_14[142], stage1_14[143], stage1_14[144], stage1_14[145]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[39],stage2_16[56],stage2_15[62],stage2_14[79]}
   );
   gpc606_5 gpc1319 (
      {stage1_14[146], stage1_14[147], stage1_14[148], stage1_14[149], stage1_14[150], stage1_14[151]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[40],stage2_16[57],stage2_15[63],stage2_14[80]}
   );
   gpc606_5 gpc1320 (
      {stage1_14[152], stage1_14[153], stage1_14[154], stage1_14[155], stage1_14[156], stage1_14[157]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[41],stage2_16[58],stage2_15[64],stage2_14[81]}
   );
   gpc606_5 gpc1321 (
      {stage1_14[158], stage1_14[159], stage1_14[160], stage1_14[161], stage1_14[162], stage1_14[163]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[42],stage2_16[59],stage2_15[65],stage2_14[82]}
   );
   gpc606_5 gpc1322 (
      {stage1_14[164], stage1_14[165], stage1_14[166], stage1_14[167], stage1_14[168], stage1_14[169]},
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage2_18[7],stage2_17[43],stage2_16[60],stage2_15[66],stage2_14[83]}
   );
   gpc606_5 gpc1323 (
      {stage1_14[170], stage1_14[171], stage1_14[172], stage1_14[173], stage1_14[174], stage1_14[175]},
      {stage1_16[48], stage1_16[49], stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53]},
      {stage2_18[8],stage2_17[44],stage2_16[61],stage2_15[67],stage2_14[84]}
   );
   gpc606_5 gpc1324 (
      {stage1_14[176], stage1_14[177], stage1_14[178], stage1_14[179], stage1_14[180], stage1_14[181]},
      {stage1_16[54], stage1_16[55], stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59]},
      {stage2_18[9],stage2_17[45],stage2_16[62],stage2_15[68],stage2_14[85]}
   );
   gpc606_5 gpc1325 (
      {stage1_14[182], stage1_14[183], stage1_14[184], stage1_14[185], stage1_14[186], stage1_14[187]},
      {stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63], stage1_16[64], stage1_16[65]},
      {stage2_18[10],stage2_17[46],stage2_16[63],stage2_15[69],stage2_14[86]}
   );
   gpc606_5 gpc1326 (
      {stage1_14[188], stage1_14[189], stage1_14[190], stage1_14[191], stage1_14[192], stage1_14[193]},
      {stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69], stage1_16[70], stage1_16[71]},
      {stage2_18[11],stage2_17[47],stage2_16[64],stage2_15[70],stage2_14[87]}
   );
   gpc606_5 gpc1327 (
      {stage1_14[194], stage1_14[195], stage1_14[196], stage1_14[197], stage1_14[198], stage1_14[199]},
      {stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75], stage1_16[76], stage1_16[77]},
      {stage2_18[12],stage2_17[48],stage2_16[65],stage2_15[71],stage2_14[88]}
   );
   gpc606_5 gpc1328 (
      {stage1_14[200], stage1_14[201], stage1_14[202], stage1_14[203], stage1_14[204], stage1_14[205]},
      {stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81], stage1_16[82], stage1_16[83]},
      {stage2_18[13],stage2_17[49],stage2_16[66],stage2_15[72],stage2_14[89]}
   );
   gpc615_5 gpc1329 (
      {stage1_14[206], stage1_14[207], stage1_14[208], stage1_14[209], stage1_14[210]},
      {stage1_15[216]},
      {stage1_16[84], stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88], stage1_16[89]},
      {stage2_18[14],stage2_17[50],stage2_16[67],stage2_15[73],stage2_14[90]}
   );
   gpc615_5 gpc1330 (
      {stage1_15[217], stage1_15[218], stage1_15[219], stage1_15[220], stage1_15[221]},
      {stage1_16[90]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[15],stage2_17[51],stage2_16[68],stage2_15[74]}
   );
   gpc615_5 gpc1331 (
      {stage1_15[222], stage1_15[223], stage1_15[224], stage1_15[225], stage1_15[226]},
      {stage1_16[91]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[16],stage2_17[52],stage2_16[69],stage2_15[75]}
   );
   gpc615_5 gpc1332 (
      {stage1_15[227], stage1_15[228], stage1_15[229], stage1_15[230], stage1_15[231]},
      {stage1_16[92]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[17],stage2_17[53],stage2_16[70],stage2_15[76]}
   );
   gpc615_5 gpc1333 (
      {stage1_15[232], stage1_15[233], stage1_15[234], stage1_15[235], stage1_15[236]},
      {stage1_16[93]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[18],stage2_17[54],stage2_16[71],stage2_15[77]}
   );
   gpc615_5 gpc1334 (
      {stage1_15[237], stage1_15[238], stage1_15[239], stage1_15[240], stage1_15[241]},
      {stage1_16[94]},
      {stage1_17[24], stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29]},
      {stage2_19[4],stage2_18[19],stage2_17[55],stage2_16[72],stage2_15[78]}
   );
   gpc615_5 gpc1335 (
      {stage1_15[242], stage1_15[243], stage1_15[244], stage1_15[245], stage1_15[246]},
      {stage1_16[95]},
      {stage1_17[30], stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35]},
      {stage2_19[5],stage2_18[20],stage2_17[56],stage2_16[73],stage2_15[79]}
   );
   gpc615_5 gpc1336 (
      {stage1_15[247], stage1_15[248], stage1_15[249], stage1_15[250], stage1_15[251]},
      {stage1_16[96]},
      {stage1_17[36], stage1_17[37], stage1_17[38], stage1_17[39], stage1_17[40], stage1_17[41]},
      {stage2_19[6],stage2_18[21],stage2_17[57],stage2_16[74],stage2_15[80]}
   );
   gpc615_5 gpc1337 (
      {stage1_15[252], stage1_15[253], stage1_15[254], stage1_15[255], stage1_15[256]},
      {stage1_16[97]},
      {stage1_17[42], stage1_17[43], stage1_17[44], stage1_17[45], stage1_17[46], stage1_17[47]},
      {stage2_19[7],stage2_18[22],stage2_17[58],stage2_16[75],stage2_15[81]}
   );
   gpc615_5 gpc1338 (
      {stage1_15[257], stage1_15[258], stage1_15[259], stage1_15[260], stage1_15[261]},
      {stage1_16[98]},
      {stage1_17[48], stage1_17[49], stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53]},
      {stage2_19[8],stage2_18[23],stage2_17[59],stage2_16[76],stage2_15[82]}
   );
   gpc615_5 gpc1339 (
      {stage1_15[262], stage1_15[263], stage1_15[264], stage1_15[265], stage1_15[266]},
      {stage1_16[99]},
      {stage1_17[54], stage1_17[55], stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59]},
      {stage2_19[9],stage2_18[24],stage2_17[60],stage2_16[77],stage2_15[83]}
   );
   gpc615_5 gpc1340 (
      {stage1_15[267], stage1_15[268], stage1_15[269], stage1_15[270], stage1_15[271]},
      {stage1_16[100]},
      {stage1_17[60], stage1_17[61], stage1_17[62], stage1_17[63], 1'b0, 1'b0},
      {stage2_19[10],stage2_18[25],stage2_17[61],stage2_16[78],stage2_15[84]}
   );
   gpc1_1 gpc1341 (
      {stage1_3[219]},
      {stage2_3[76]}
   );
   gpc1_1 gpc1342 (
      {stage1_3[220]},
      {stage2_3[77]}
   );
   gpc1_1 gpc1343 (
      {stage1_3[221]},
      {stage2_3[78]}
   );
   gpc1_1 gpc1344 (
      {stage1_3[222]},
      {stage2_3[79]}
   );
   gpc1_1 gpc1345 (
      {stage1_3[223]},
      {stage2_3[80]}
   );
   gpc1_1 gpc1346 (
      {stage1_3[224]},
      {stage2_3[81]}
   );
   gpc1_1 gpc1347 (
      {stage1_3[225]},
      {stage2_3[82]}
   );
   gpc1_1 gpc1348 (
      {stage1_3[226]},
      {stage2_3[83]}
   );
   gpc1_1 gpc1349 (
      {stage1_3[227]},
      {stage2_3[84]}
   );
   gpc1_1 gpc1350 (
      {stage1_3[228]},
      {stage2_3[85]}
   );
   gpc1_1 gpc1351 (
      {stage1_3[229]},
      {stage2_3[86]}
   );
   gpc1_1 gpc1352 (
      {stage1_3[230]},
      {stage2_3[87]}
   );
   gpc1_1 gpc1353 (
      {stage1_3[231]},
      {stage2_3[88]}
   );
   gpc1_1 gpc1354 (
      {stage1_3[232]},
      {stage2_3[89]}
   );
   gpc1_1 gpc1355 (
      {stage1_3[233]},
      {stage2_3[90]}
   );
   gpc1_1 gpc1356 (
      {stage1_3[234]},
      {stage2_3[91]}
   );
   gpc1_1 gpc1357 (
      {stage1_3[235]},
      {stage2_3[92]}
   );
   gpc1_1 gpc1358 (
      {stage1_3[236]},
      {stage2_3[93]}
   );
   gpc1_1 gpc1359 (
      {stage1_3[237]},
      {stage2_3[94]}
   );
   gpc1_1 gpc1360 (
      {stage1_3[238]},
      {stage2_3[95]}
   );
   gpc1_1 gpc1361 (
      {stage1_3[239]},
      {stage2_3[96]}
   );
   gpc1_1 gpc1362 (
      {stage1_3[240]},
      {stage2_3[97]}
   );
   gpc1_1 gpc1363 (
      {stage1_3[241]},
      {stage2_3[98]}
   );
   gpc1_1 gpc1364 (
      {stage1_3[242]},
      {stage2_3[99]}
   );
   gpc1_1 gpc1365 (
      {stage1_3[243]},
      {stage2_3[100]}
   );
   gpc1_1 gpc1366 (
      {stage1_3[244]},
      {stage2_3[101]}
   );
   gpc1_1 gpc1367 (
      {stage1_3[245]},
      {stage2_3[102]}
   );
   gpc1_1 gpc1368 (
      {stage1_4[214]},
      {stage2_4[90]}
   );
   gpc1_1 gpc1369 (
      {stage1_4[215]},
      {stage2_4[91]}
   );
   gpc1_1 gpc1370 (
      {stage1_4[216]},
      {stage2_4[92]}
   );
   gpc1_1 gpc1371 (
      {stage1_4[217]},
      {stage2_4[93]}
   );
   gpc1_1 gpc1372 (
      {stage1_4[218]},
      {stage2_4[94]}
   );
   gpc1_1 gpc1373 (
      {stage1_4[219]},
      {stage2_4[95]}
   );
   gpc1_1 gpc1374 (
      {stage1_4[220]},
      {stage2_4[96]}
   );
   gpc1_1 gpc1375 (
      {stage1_4[221]},
      {stage2_4[97]}
   );
   gpc1_1 gpc1376 (
      {stage1_4[222]},
      {stage2_4[98]}
   );
   gpc1_1 gpc1377 (
      {stage1_4[223]},
      {stage2_4[99]}
   );
   gpc1_1 gpc1378 (
      {stage1_4[224]},
      {stage2_4[100]}
   );
   gpc1_1 gpc1379 (
      {stage1_4[225]},
      {stage2_4[101]}
   );
   gpc1_1 gpc1380 (
      {stage1_4[226]},
      {stage2_4[102]}
   );
   gpc1_1 gpc1381 (
      {stage1_4[227]},
      {stage2_4[103]}
   );
   gpc1_1 gpc1382 (
      {stage1_4[228]},
      {stage2_4[104]}
   );
   gpc1_1 gpc1383 (
      {stage1_4[229]},
      {stage2_4[105]}
   );
   gpc1_1 gpc1384 (
      {stage1_4[230]},
      {stage2_4[106]}
   );
   gpc1_1 gpc1385 (
      {stage1_4[231]},
      {stage2_4[107]}
   );
   gpc1_1 gpc1386 (
      {stage1_4[232]},
      {stage2_4[108]}
   );
   gpc1_1 gpc1387 (
      {stage1_4[233]},
      {stage2_4[109]}
   );
   gpc1_1 gpc1388 (
      {stage1_4[234]},
      {stage2_4[110]}
   );
   gpc1_1 gpc1389 (
      {stage1_4[235]},
      {stage2_4[111]}
   );
   gpc1_1 gpc1390 (
      {stage1_4[236]},
      {stage2_4[112]}
   );
   gpc1_1 gpc1391 (
      {stage1_4[237]},
      {stage2_4[113]}
   );
   gpc1_1 gpc1392 (
      {stage1_4[238]},
      {stage2_4[114]}
   );
   gpc1_1 gpc1393 (
      {stage1_4[239]},
      {stage2_4[115]}
   );
   gpc1_1 gpc1394 (
      {stage1_4[240]},
      {stage2_4[116]}
   );
   gpc1_1 gpc1395 (
      {stage1_5[210]},
      {stage2_5[86]}
   );
   gpc1_1 gpc1396 (
      {stage1_5[211]},
      {stage2_5[87]}
   );
   gpc1_1 gpc1397 (
      {stage1_5[212]},
      {stage2_5[88]}
   );
   gpc1_1 gpc1398 (
      {stage1_5[213]},
      {stage2_5[89]}
   );
   gpc1_1 gpc1399 (
      {stage1_5[214]},
      {stage2_5[90]}
   );
   gpc1_1 gpc1400 (
      {stage1_5[215]},
      {stage2_5[91]}
   );
   gpc1_1 gpc1401 (
      {stage1_5[216]},
      {stage2_5[92]}
   );
   gpc1_1 gpc1402 (
      {stage1_5[217]},
      {stage2_5[93]}
   );
   gpc1_1 gpc1403 (
      {stage1_6[189]},
      {stage2_6[86]}
   );
   gpc1_1 gpc1404 (
      {stage1_6[190]},
      {stage2_6[87]}
   );
   gpc1_1 gpc1405 (
      {stage1_6[191]},
      {stage2_6[88]}
   );
   gpc1_1 gpc1406 (
      {stage1_6[192]},
      {stage2_6[89]}
   );
   gpc1_1 gpc1407 (
      {stage1_6[193]},
      {stage2_6[90]}
   );
   gpc1_1 gpc1408 (
      {stage1_6[194]},
      {stage2_6[91]}
   );
   gpc1_1 gpc1409 (
      {stage1_6[195]},
      {stage2_6[92]}
   );
   gpc1_1 gpc1410 (
      {stage1_6[196]},
      {stage2_6[93]}
   );
   gpc1_1 gpc1411 (
      {stage1_6[197]},
      {stage2_6[94]}
   );
   gpc1_1 gpc1412 (
      {stage1_6[198]},
      {stage2_6[95]}
   );
   gpc1_1 gpc1413 (
      {stage1_6[199]},
      {stage2_6[96]}
   );
   gpc1_1 gpc1414 (
      {stage1_6[200]},
      {stage2_6[97]}
   );
   gpc1_1 gpc1415 (
      {stage1_6[201]},
      {stage2_6[98]}
   );
   gpc1_1 gpc1416 (
      {stage1_6[202]},
      {stage2_6[99]}
   );
   gpc1_1 gpc1417 (
      {stage1_6[203]},
      {stage2_6[100]}
   );
   gpc1_1 gpc1418 (
      {stage1_6[204]},
      {stage2_6[101]}
   );
   gpc1_1 gpc1419 (
      {stage1_6[205]},
      {stage2_6[102]}
   );
   gpc1_1 gpc1420 (
      {stage1_6[206]},
      {stage2_6[103]}
   );
   gpc1_1 gpc1421 (
      {stage1_9[214]},
      {stage2_9[88]}
   );
   gpc1_1 gpc1422 (
      {stage1_9[215]},
      {stage2_9[89]}
   );
   gpc1_1 gpc1423 (
      {stage1_9[216]},
      {stage2_9[90]}
   );
   gpc1_1 gpc1424 (
      {stage1_9[217]},
      {stage2_9[91]}
   );
   gpc1_1 gpc1425 (
      {stage1_9[218]},
      {stage2_9[92]}
   );
   gpc1_1 gpc1426 (
      {stage1_9[219]},
      {stage2_9[93]}
   );
   gpc1_1 gpc1427 (
      {stage1_9[220]},
      {stage2_9[94]}
   );
   gpc1_1 gpc1428 (
      {stage1_9[221]},
      {stage2_9[95]}
   );
   gpc1_1 gpc1429 (
      {stage1_9[222]},
      {stage2_9[96]}
   );
   gpc1_1 gpc1430 (
      {stage1_9[223]},
      {stage2_9[97]}
   );
   gpc1_1 gpc1431 (
      {stage1_9[224]},
      {stage2_9[98]}
   );
   gpc1_1 gpc1432 (
      {stage1_9[225]},
      {stage2_9[99]}
   );
   gpc1_1 gpc1433 (
      {stage1_9[226]},
      {stage2_9[100]}
   );
   gpc1_1 gpc1434 (
      {stage1_9[227]},
      {stage2_9[101]}
   );
   gpc1_1 gpc1435 (
      {stage1_9[228]},
      {stage2_9[102]}
   );
   gpc1_1 gpc1436 (
      {stage1_9[229]},
      {stage2_9[103]}
   );
   gpc1_1 gpc1437 (
      {stage1_9[230]},
      {stage2_9[104]}
   );
   gpc1_1 gpc1438 (
      {stage1_9[231]},
      {stage2_9[105]}
   );
   gpc1_1 gpc1439 (
      {stage1_9[232]},
      {stage2_9[106]}
   );
   gpc1_1 gpc1440 (
      {stage1_9[233]},
      {stage2_9[107]}
   );
   gpc1_1 gpc1441 (
      {stage1_9[234]},
      {stage2_9[108]}
   );
   gpc1_1 gpc1442 (
      {stage1_9[235]},
      {stage2_9[109]}
   );
   gpc1_1 gpc1443 (
      {stage1_9[236]},
      {stage2_9[110]}
   );
   gpc1_1 gpc1444 (
      {stage1_9[237]},
      {stage2_9[111]}
   );
   gpc1_1 gpc1445 (
      {stage1_9[238]},
      {stage2_9[112]}
   );
   gpc1_1 gpc1446 (
      {stage1_9[239]},
      {stage2_9[113]}
   );
   gpc1_1 gpc1447 (
      {stage1_9[240]},
      {stage2_9[114]}
   );
   gpc1_1 gpc1448 (
      {stage1_9[241]},
      {stage2_9[115]}
   );
   gpc1_1 gpc1449 (
      {stage1_9[242]},
      {stage2_9[116]}
   );
   gpc1_1 gpc1450 (
      {stage1_9[243]},
      {stage2_9[117]}
   );
   gpc1_1 gpc1451 (
      {stage1_9[244]},
      {stage2_9[118]}
   );
   gpc1_1 gpc1452 (
      {stage1_9[245]},
      {stage2_9[119]}
   );
   gpc1_1 gpc1453 (
      {stage1_9[246]},
      {stage2_9[120]}
   );
   gpc1_1 gpc1454 (
      {stage1_9[247]},
      {stage2_9[121]}
   );
   gpc1_1 gpc1455 (
      {stage1_9[248]},
      {stage2_9[122]}
   );
   gpc1_1 gpc1456 (
      {stage1_9[249]},
      {stage2_9[123]}
   );
   gpc1_1 gpc1457 (
      {stage1_9[250]},
      {stage2_9[124]}
   );
   gpc1_1 gpc1458 (
      {stage1_9[251]},
      {stage2_9[125]}
   );
   gpc1_1 gpc1459 (
      {stage1_9[252]},
      {stage2_9[126]}
   );
   gpc1_1 gpc1460 (
      {stage1_9[253]},
      {stage2_9[127]}
   );
   gpc1_1 gpc1461 (
      {stage1_9[254]},
      {stage2_9[128]}
   );
   gpc1_1 gpc1462 (
      {stage1_9[255]},
      {stage2_9[129]}
   );
   gpc1_1 gpc1463 (
      {stage1_9[256]},
      {stage2_9[130]}
   );
   gpc1_1 gpc1464 (
      {stage1_9[257]},
      {stage2_9[131]}
   );
   gpc1_1 gpc1465 (
      {stage1_9[258]},
      {stage2_9[132]}
   );
   gpc1_1 gpc1466 (
      {stage1_9[259]},
      {stage2_9[133]}
   );
   gpc1_1 gpc1467 (
      {stage1_9[260]},
      {stage2_9[134]}
   );
   gpc1_1 gpc1468 (
      {stage1_9[261]},
      {stage2_9[135]}
   );
   gpc1_1 gpc1469 (
      {stage1_9[262]},
      {stage2_9[136]}
   );
   gpc1_1 gpc1470 (
      {stage1_9[263]},
      {stage2_9[137]}
   );
   gpc1_1 gpc1471 (
      {stage1_11[120]},
      {stage2_11[74]}
   );
   gpc1_1 gpc1472 (
      {stage1_11[121]},
      {stage2_11[75]}
   );
   gpc1_1 gpc1473 (
      {stage1_11[122]},
      {stage2_11[76]}
   );
   gpc1_1 gpc1474 (
      {stage1_11[123]},
      {stage2_11[77]}
   );
   gpc1_1 gpc1475 (
      {stage1_11[124]},
      {stage2_11[78]}
   );
   gpc1_1 gpc1476 (
      {stage1_11[125]},
      {stage2_11[79]}
   );
   gpc1_1 gpc1477 (
      {stage1_11[126]},
      {stage2_11[80]}
   );
   gpc1_1 gpc1478 (
      {stage1_11[127]},
      {stage2_11[81]}
   );
   gpc1_1 gpc1479 (
      {stage1_11[128]},
      {stage2_11[82]}
   );
   gpc1_1 gpc1480 (
      {stage1_11[129]},
      {stage2_11[83]}
   );
   gpc1_1 gpc1481 (
      {stage1_11[130]},
      {stage2_11[84]}
   );
   gpc1_1 gpc1482 (
      {stage1_11[131]},
      {stage2_11[85]}
   );
   gpc1_1 gpc1483 (
      {stage1_11[132]},
      {stage2_11[86]}
   );
   gpc1_1 gpc1484 (
      {stage1_11[133]},
      {stage2_11[87]}
   );
   gpc1_1 gpc1485 (
      {stage1_11[134]},
      {stage2_11[88]}
   );
   gpc1_1 gpc1486 (
      {stage1_11[135]},
      {stage2_11[89]}
   );
   gpc1_1 gpc1487 (
      {stage1_11[136]},
      {stage2_11[90]}
   );
   gpc1_1 gpc1488 (
      {stage1_11[137]},
      {stage2_11[91]}
   );
   gpc1_1 gpc1489 (
      {stage1_11[138]},
      {stage2_11[92]}
   );
   gpc1_1 gpc1490 (
      {stage1_11[139]},
      {stage2_11[93]}
   );
   gpc1_1 gpc1491 (
      {stage1_11[140]},
      {stage2_11[94]}
   );
   gpc1_1 gpc1492 (
      {stage1_11[141]},
      {stage2_11[95]}
   );
   gpc1_1 gpc1493 (
      {stage1_11[142]},
      {stage2_11[96]}
   );
   gpc1_1 gpc1494 (
      {stage1_11[143]},
      {stage2_11[97]}
   );
   gpc1_1 gpc1495 (
      {stage1_11[144]},
      {stage2_11[98]}
   );
   gpc1_1 gpc1496 (
      {stage1_11[145]},
      {stage2_11[99]}
   );
   gpc1_1 gpc1497 (
      {stage1_11[146]},
      {stage2_11[100]}
   );
   gpc1_1 gpc1498 (
      {stage1_11[147]},
      {stage2_11[101]}
   );
   gpc1_1 gpc1499 (
      {stage1_11[148]},
      {stage2_11[102]}
   );
   gpc1_1 gpc1500 (
      {stage1_11[149]},
      {stage2_11[103]}
   );
   gpc1_1 gpc1501 (
      {stage1_11[150]},
      {stage2_11[104]}
   );
   gpc1_1 gpc1502 (
      {stage1_11[151]},
      {stage2_11[105]}
   );
   gpc1_1 gpc1503 (
      {stage1_11[152]},
      {stage2_11[106]}
   );
   gpc1_1 gpc1504 (
      {stage1_11[153]},
      {stage2_11[107]}
   );
   gpc1_1 gpc1505 (
      {stage1_11[154]},
      {stage2_11[108]}
   );
   gpc1_1 gpc1506 (
      {stage1_11[155]},
      {stage2_11[109]}
   );
   gpc1_1 gpc1507 (
      {stage1_11[156]},
      {stage2_11[110]}
   );
   gpc1_1 gpc1508 (
      {stage1_11[157]},
      {stage2_11[111]}
   );
   gpc1_1 gpc1509 (
      {stage1_11[158]},
      {stage2_11[112]}
   );
   gpc1_1 gpc1510 (
      {stage1_11[159]},
      {stage2_11[113]}
   );
   gpc1_1 gpc1511 (
      {stage1_11[160]},
      {stage2_11[114]}
   );
   gpc1_1 gpc1512 (
      {stage1_11[161]},
      {stage2_11[115]}
   );
   gpc1_1 gpc1513 (
      {stage1_11[162]},
      {stage2_11[116]}
   );
   gpc1_1 gpc1514 (
      {stage1_11[163]},
      {stage2_11[117]}
   );
   gpc1_1 gpc1515 (
      {stage1_11[164]},
      {stage2_11[118]}
   );
   gpc1_1 gpc1516 (
      {stage1_11[165]},
      {stage2_11[119]}
   );
   gpc1_1 gpc1517 (
      {stage1_11[166]},
      {stage2_11[120]}
   );
   gpc1_1 gpc1518 (
      {stage1_11[167]},
      {stage2_11[121]}
   );
   gpc1_1 gpc1519 (
      {stage1_11[168]},
      {stage2_11[122]}
   );
   gpc1_1 gpc1520 (
      {stage1_11[169]},
      {stage2_11[123]}
   );
   gpc1_1 gpc1521 (
      {stage1_11[170]},
      {stage2_11[124]}
   );
   gpc1_1 gpc1522 (
      {stage1_11[171]},
      {stage2_11[125]}
   );
   gpc1_1 gpc1523 (
      {stage1_11[172]},
      {stage2_11[126]}
   );
   gpc1_1 gpc1524 (
      {stage1_11[173]},
      {stage2_11[127]}
   );
   gpc1_1 gpc1525 (
      {stage1_11[174]},
      {stage2_11[128]}
   );
   gpc1_1 gpc1526 (
      {stage1_11[175]},
      {stage2_11[129]}
   );
   gpc1_1 gpc1527 (
      {stage1_11[176]},
      {stage2_11[130]}
   );
   gpc1_1 gpc1528 (
      {stage1_11[177]},
      {stage2_11[131]}
   );
   gpc1_1 gpc1529 (
      {stage1_11[178]},
      {stage2_11[132]}
   );
   gpc1_1 gpc1530 (
      {stage1_11[179]},
      {stage2_11[133]}
   );
   gpc1_1 gpc1531 (
      {stage1_11[180]},
      {stage2_11[134]}
   );
   gpc1_1 gpc1532 (
      {stage1_11[181]},
      {stage2_11[135]}
   );
   gpc1_1 gpc1533 (
      {stage1_11[182]},
      {stage2_11[136]}
   );
   gpc1_1 gpc1534 (
      {stage1_11[183]},
      {stage2_11[137]}
   );
   gpc1_1 gpc1535 (
      {stage1_11[184]},
      {stage2_11[138]}
   );
   gpc1_1 gpc1536 (
      {stage1_11[185]},
      {stage2_11[139]}
   );
   gpc1_1 gpc1537 (
      {stage1_11[186]},
      {stage2_11[140]}
   );
   gpc1_1 gpc1538 (
      {stage1_11[187]},
      {stage2_11[141]}
   );
   gpc1_1 gpc1539 (
      {stage1_11[188]},
      {stage2_11[142]}
   );
   gpc1_1 gpc1540 (
      {stage1_11[189]},
      {stage2_11[143]}
   );
   gpc1_1 gpc1541 (
      {stage1_12[210]},
      {stage2_12[73]}
   );
   gpc1_1 gpc1542 (
      {stage1_12[211]},
      {stage2_12[74]}
   );
   gpc1_1 gpc1543 (
      {stage1_12[212]},
      {stage2_12[75]}
   );
   gpc1_1 gpc1544 (
      {stage1_12[213]},
      {stage2_12[76]}
   );
   gpc1_1 gpc1545 (
      {stage1_12[214]},
      {stage2_12[77]}
   );
   gpc1_1 gpc1546 (
      {stage1_12[215]},
      {stage2_12[78]}
   );
   gpc1_1 gpc1547 (
      {stage1_12[216]},
      {stage2_12[79]}
   );
   gpc1_1 gpc1548 (
      {stage1_12[217]},
      {stage2_12[80]}
   );
   gpc1_1 gpc1549 (
      {stage1_12[218]},
      {stage2_12[81]}
   );
   gpc1_1 gpc1550 (
      {stage1_12[219]},
      {stage2_12[82]}
   );
   gpc1_1 gpc1551 (
      {stage1_12[220]},
      {stage2_12[83]}
   );
   gpc1_1 gpc1552 (
      {stage1_12[221]},
      {stage2_12[84]}
   );
   gpc1_1 gpc1553 (
      {stage1_13[232]},
      {stage2_13[91]}
   );
   gpc1_1 gpc1554 (
      {stage1_13[233]},
      {stage2_13[92]}
   );
   gpc1_1 gpc1555 (
      {stage1_13[234]},
      {stage2_13[93]}
   );
   gpc1_1 gpc1556 (
      {stage1_13[235]},
      {stage2_13[94]}
   );
   gpc1_1 gpc1557 (
      {stage1_13[236]},
      {stage2_13[95]}
   );
   gpc1_1 gpc1558 (
      {stage1_13[237]},
      {stage2_13[96]}
   );
   gpc1_1 gpc1559 (
      {stage1_13[238]},
      {stage2_13[97]}
   );
   gpc1_1 gpc1560 (
      {stage1_13[239]},
      {stage2_13[98]}
   );
   gpc1_1 gpc1561 (
      {stage1_13[240]},
      {stage2_13[99]}
   );
   gpc1_1 gpc1562 (
      {stage1_13[241]},
      {stage2_13[100]}
   );
   gpc1_1 gpc1563 (
      {stage1_13[242]},
      {stage2_13[101]}
   );
   gpc1_1 gpc1564 (
      {stage1_13[243]},
      {stage2_13[102]}
   );
   gpc1_1 gpc1565 (
      {stage1_13[244]},
      {stage2_13[103]}
   );
   gpc1_1 gpc1566 (
      {stage1_13[245]},
      {stage2_13[104]}
   );
   gpc1_1 gpc1567 (
      {stage1_13[246]},
      {stage2_13[105]}
   );
   gpc1_1 gpc1568 (
      {stage1_13[247]},
      {stage2_13[106]}
   );
   gpc1_1 gpc1569 (
      {stage1_13[248]},
      {stage2_13[107]}
   );
   gpc1_1 gpc1570 (
      {stage1_13[249]},
      {stage2_13[108]}
   );
   gpc1_1 gpc1571 (
      {stage1_13[250]},
      {stage2_13[109]}
   );
   gpc1_1 gpc1572 (
      {stage1_13[251]},
      {stage2_13[110]}
   );
   gpc1_1 gpc1573 (
      {stage1_13[252]},
      {stage2_13[111]}
   );
   gpc1_1 gpc1574 (
      {stage1_13[253]},
      {stage2_13[112]}
   );
   gpc1_1 gpc1575 (
      {stage1_13[254]},
      {stage2_13[113]}
   );
   gpc1_1 gpc1576 (
      {stage1_13[255]},
      {stage2_13[114]}
   );
   gpc1_1 gpc1577 (
      {stage1_13[256]},
      {stage2_13[115]}
   );
   gpc1_1 gpc1578 (
      {stage1_13[257]},
      {stage2_13[116]}
   );
   gpc1_1 gpc1579 (
      {stage1_13[258]},
      {stage2_13[117]}
   );
   gpc1_1 gpc1580 (
      {stage1_13[259]},
      {stage2_13[118]}
   );
   gpc1_1 gpc1581 (
      {stage1_13[260]},
      {stage2_13[119]}
   );
   gpc1_1 gpc1582 (
      {stage1_13[261]},
      {stage2_13[120]}
   );
   gpc1_1 gpc1583 (
      {stage1_13[262]},
      {stage2_13[121]}
   );
   gpc1_1 gpc1584 (
      {stage1_13[263]},
      {stage2_13[122]}
   );
   gpc1_1 gpc1585 (
      {stage1_13[264]},
      {stage2_13[123]}
   );
   gpc1_1 gpc1586 (
      {stage1_13[265]},
      {stage2_13[124]}
   );
   gpc1_1 gpc1587 (
      {stage1_13[266]},
      {stage2_13[125]}
   );
   gpc1_1 gpc1588 (
      {stage1_13[267]},
      {stage2_13[126]}
   );
   gpc1_1 gpc1589 (
      {stage1_13[268]},
      {stage2_13[127]}
   );
   gpc1_1 gpc1590 (
      {stage1_13[269]},
      {stage2_13[128]}
   );
   gpc1_1 gpc1591 (
      {stage1_13[270]},
      {stage2_13[129]}
   );
   gpc1_1 gpc1592 (
      {stage1_13[271]},
      {stage2_13[130]}
   );
   gpc1_1 gpc1593 (
      {stage1_13[272]},
      {stage2_13[131]}
   );
   gpc1_1 gpc1594 (
      {stage1_13[273]},
      {stage2_13[132]}
   );
   gpc1_1 gpc1595 (
      {stage1_13[274]},
      {stage2_13[133]}
   );
   gpc1_1 gpc1596 (
      {stage1_13[275]},
      {stage2_13[134]}
   );
   gpc1_1 gpc1597 (
      {stage1_13[276]},
      {stage2_13[135]}
   );
   gpc1_1 gpc1598 (
      {stage1_13[277]},
      {stage2_13[136]}
   );
   gpc1_1 gpc1599 (
      {stage1_13[278]},
      {stage2_13[137]}
   );
   gpc1_1 gpc1600 (
      {stage1_13[279]},
      {stage2_13[138]}
   );
   gpc1_1 gpc1601 (
      {stage1_13[280]},
      {stage2_13[139]}
   );
   gpc1_1 gpc1602 (
      {stage1_13[281]},
      {stage2_13[140]}
   );
   gpc1_1 gpc1603 (
      {stage1_14[211]},
      {stage2_14[91]}
   );
   gpc1_1 gpc1604 (
      {stage1_14[212]},
      {stage2_14[92]}
   );
   gpc1_1 gpc1605 (
      {stage1_14[213]},
      {stage2_14[93]}
   );
   gpc1_1 gpc1606 (
      {stage1_14[214]},
      {stage2_14[94]}
   );
   gpc1_1 gpc1607 (
      {stage1_14[215]},
      {stage2_14[95]}
   );
   gpc1_1 gpc1608 (
      {stage1_14[216]},
      {stage2_14[96]}
   );
   gpc1_1 gpc1609 (
      {stage1_14[217]},
      {stage2_14[97]}
   );
   gpc1_1 gpc1610 (
      {stage1_14[218]},
      {stage2_14[98]}
   );
   gpc1_1 gpc1611 (
      {stage1_14[219]},
      {stage2_14[99]}
   );
   gpc1_1 gpc1612 (
      {stage1_14[220]},
      {stage2_14[100]}
   );
   gpc1_1 gpc1613 (
      {stage1_14[221]},
      {stage2_14[101]}
   );
   gpc1_1 gpc1614 (
      {stage1_14[222]},
      {stage2_14[102]}
   );
   gpc1_1 gpc1615 (
      {stage1_14[223]},
      {stage2_14[103]}
   );
   gpc1_1 gpc1616 (
      {stage1_14[224]},
      {stage2_14[104]}
   );
   gpc1_1 gpc1617 (
      {stage1_14[225]},
      {stage2_14[105]}
   );
   gpc1_1 gpc1618 (
      {stage1_14[226]},
      {stage2_14[106]}
   );
   gpc1_1 gpc1619 (
      {stage1_14[227]},
      {stage2_14[107]}
   );
   gpc1_1 gpc1620 (
      {stage1_14[228]},
      {stage2_14[108]}
   );
   gpc1_1 gpc1621 (
      {stage1_14[229]},
      {stage2_14[109]}
   );
   gpc1_1 gpc1622 (
      {stage1_14[230]},
      {stage2_14[110]}
   );
   gpc1_1 gpc1623 (
      {stage1_14[231]},
      {stage2_14[111]}
   );
   gpc1_1 gpc1624 (
      {stage1_14[232]},
      {stage2_14[112]}
   );
   gpc1_1 gpc1625 (
      {stage1_14[233]},
      {stage2_14[113]}
   );
   gpc1_1 gpc1626 (
      {stage1_14[234]},
      {stage2_14[114]}
   );
   gpc1_1 gpc1627 (
      {stage1_14[235]},
      {stage2_14[115]}
   );
   gpc1_1 gpc1628 (
      {stage1_14[236]},
      {stage2_14[116]}
   );
   gpc1_1 gpc1629 (
      {stage1_14[237]},
      {stage2_14[117]}
   );
   gpc1_1 gpc1630 (
      {stage1_14[238]},
      {stage2_14[118]}
   );
   gpc1_1 gpc1631 (
      {stage1_14[239]},
      {stage2_14[119]}
   );
   gpc1_1 gpc1632 (
      {stage1_14[240]},
      {stage2_14[120]}
   );
   gpc1_1 gpc1633 (
      {stage1_14[241]},
      {stage2_14[121]}
   );
   gpc1_1 gpc1634 (
      {stage1_14[242]},
      {stage2_14[122]}
   );
   gpc1_1 gpc1635 (
      {stage1_14[243]},
      {stage2_14[123]}
   );
   gpc1_1 gpc1636 (
      {stage1_14[244]},
      {stage2_14[124]}
   );
   gpc1_1 gpc1637 (
      {stage1_16[101]},
      {stage2_16[79]}
   );
   gpc1_1 gpc1638 (
      {stage1_16[102]},
      {stage2_16[80]}
   );
   gpc1_1 gpc1639 (
      {stage1_16[103]},
      {stage2_16[81]}
   );
   gpc1_1 gpc1640 (
      {stage1_16[104]},
      {stage2_16[82]}
   );
   gpc1_1 gpc1641 (
      {stage1_16[105]},
      {stage2_16[83]}
   );
   gpc1_1 gpc1642 (
      {stage1_16[106]},
      {stage2_16[84]}
   );
   gpc1_1 gpc1643 (
      {stage1_16[107]},
      {stage2_16[85]}
   );
   gpc1_1 gpc1644 (
      {stage1_16[108]},
      {stage2_16[86]}
   );
   gpc1_1 gpc1645 (
      {stage1_16[109]},
      {stage2_16[87]}
   );
   gpc1_1 gpc1646 (
      {stage1_16[110]},
      {stage2_16[88]}
   );
   gpc1_1 gpc1647 (
      {stage1_16[111]},
      {stage2_16[89]}
   );
   gpc1_1 gpc1648 (
      {stage1_16[112]},
      {stage2_16[90]}
   );
   gpc1_1 gpc1649 (
      {stage1_16[113]},
      {stage2_16[91]}
   );
   gpc1_1 gpc1650 (
      {stage1_16[114]},
      {stage2_16[92]}
   );
   gpc1_1 gpc1651 (
      {stage1_16[115]},
      {stage2_16[93]}
   );
   gpc1_1 gpc1652 (
      {stage1_16[116]},
      {stage2_16[94]}
   );
   gpc1_1 gpc1653 (
      {stage1_16[117]},
      {stage2_16[95]}
   );
   gpc1_1 gpc1654 (
      {stage1_16[118]},
      {stage2_16[96]}
   );
   gpc1_1 gpc1655 (
      {stage1_16[119]},
      {stage2_16[97]}
   );
   gpc1_1 gpc1656 (
      {stage1_16[120]},
      {stage2_16[98]}
   );
   gpc1_1 gpc1657 (
      {stage1_16[121]},
      {stage2_16[99]}
   );
   gpc1_1 gpc1658 (
      {stage1_16[122]},
      {stage2_16[100]}
   );
   gpc1_1 gpc1659 (
      {stage1_16[123]},
      {stage2_16[101]}
   );
   gpc1_1 gpc1660 (
      {stage1_16[124]},
      {stage2_16[102]}
   );
   gpc1_1 gpc1661 (
      {stage1_16[125]},
      {stage2_16[103]}
   );
   gpc1_1 gpc1662 (
      {stage1_16[126]},
      {stage2_16[104]}
   );
   gpc606_5 gpc1663 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc615_5 gpc1664 (
      {stage2_0[6], stage2_0[7], stage2_0[8], stage2_0[9], stage2_0[10]},
      {stage2_1[0]},
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc615_5 gpc1665 (
      {stage2_0[11], stage2_0[12], stage2_0[13], stage2_0[14], stage2_0[15]},
      {stage2_1[1]},
      {stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc615_5 gpc1666 (
      {stage2_0[16], stage2_0[17], stage2_0[18], stage2_0[19], stage2_0[20]},
      {stage2_1[2]},
      {stage2_2[18], stage2_2[19], stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc606_5 gpc1667 (
      {stage2_1[3], stage2_1[4], stage2_1[5], stage2_1[6], stage2_1[7], stage2_1[8]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4]}
   );
   gpc606_5 gpc1668 (
      {stage2_1[9], stage2_1[10], stage2_1[11], stage2_1[12], stage2_1[13], stage2_1[14]},
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage3_5[1],stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5]}
   );
   gpc606_5 gpc1669 (
      {stage2_1[15], stage2_1[16], stage2_1[17], stage2_1[18], stage2_1[19], stage2_1[20]},
      {stage2_3[12], stage2_3[13], stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17]},
      {stage3_5[2],stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6]}
   );
   gpc606_5 gpc1670 (
      {stage2_1[21], stage2_1[22], stage2_1[23], stage2_1[24], stage2_1[25], stage2_1[26]},
      {stage2_3[18], stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23]},
      {stage3_5[3],stage3_4[7],stage3_3[7],stage3_2[7],stage3_1[7]}
   );
   gpc606_5 gpc1671 (
      {stage2_1[27], stage2_1[28], stage2_1[29], stage2_1[30], stage2_1[31], stage2_1[32]},
      {stage2_3[24], stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29]},
      {stage3_5[4],stage3_4[8],stage3_3[8],stage3_2[8],stage3_1[8]}
   );
   gpc606_5 gpc1672 (
      {stage2_1[33], stage2_1[34], stage2_1[35], stage2_1[36], stage2_1[37], stage2_1[38]},
      {stage2_3[30], stage2_3[31], stage2_3[32], stage2_3[33], stage2_3[34], stage2_3[35]},
      {stage3_5[5],stage3_4[9],stage3_3[9],stage3_2[9],stage3_1[9]}
   );
   gpc606_5 gpc1673 (
      {stage2_2[24], stage2_2[25], stage2_2[26], stage2_2[27], stage2_2[28], stage2_2[29]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[6],stage3_4[10],stage3_3[10],stage3_2[10]}
   );
   gpc615_5 gpc1674 (
      {stage2_2[30], stage2_2[31], stage2_2[32], stage2_2[33], stage2_2[34]},
      {stage2_3[36]},
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage3_6[1],stage3_5[7],stage3_4[11],stage3_3[11],stage3_2[11]}
   );
   gpc615_5 gpc1675 (
      {stage2_2[35], stage2_2[36], stage2_2[37], stage2_2[38], stage2_2[39]},
      {stage2_3[37]},
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage3_6[2],stage3_5[8],stage3_4[12],stage3_3[12],stage3_2[12]}
   );
   gpc615_5 gpc1676 (
      {stage2_2[40], stage2_2[41], stage2_2[42], stage2_2[43], stage2_2[44]},
      {stage2_3[38]},
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23]},
      {stage3_6[3],stage3_5[9],stage3_4[13],stage3_3[13],stage3_2[13]}
   );
   gpc615_5 gpc1677 (
      {stage2_2[45], stage2_2[46], stage2_2[47], stage2_2[48], stage2_2[49]},
      {stage2_3[39]},
      {stage2_4[24], stage2_4[25], stage2_4[26], stage2_4[27], stage2_4[28], stage2_4[29]},
      {stage3_6[4],stage3_5[10],stage3_4[14],stage3_3[14],stage3_2[14]}
   );
   gpc615_5 gpc1678 (
      {stage2_2[50], stage2_2[51], stage2_2[52], stage2_2[53], stage2_2[54]},
      {stage2_3[40]},
      {stage2_4[30], stage2_4[31], stage2_4[32], stage2_4[33], stage2_4[34], stage2_4[35]},
      {stage3_6[5],stage3_5[11],stage3_4[15],stage3_3[15],stage3_2[15]}
   );
   gpc615_5 gpc1679 (
      {stage2_2[55], stage2_2[56], stage2_2[57], stage2_2[58], stage2_2[59]},
      {stage2_3[41]},
      {stage2_4[36], stage2_4[37], stage2_4[38], stage2_4[39], stage2_4[40], stage2_4[41]},
      {stage3_6[6],stage3_5[12],stage3_4[16],stage3_3[16],stage3_2[16]}
   );
   gpc606_5 gpc1680 (
      {stage2_3[42], stage2_3[43], stage2_3[44], stage2_3[45], stage2_3[46], stage2_3[47]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[7],stage3_5[13],stage3_4[17],stage3_3[17]}
   );
   gpc615_5 gpc1681 (
      {stage2_3[48], stage2_3[49], stage2_3[50], stage2_3[51], stage2_3[52]},
      {stage2_4[42]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[8],stage3_5[14],stage3_4[18],stage3_3[18]}
   );
   gpc615_5 gpc1682 (
      {stage2_3[53], stage2_3[54], stage2_3[55], stage2_3[56], stage2_3[57]},
      {stage2_4[43]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[9],stage3_5[15],stage3_4[19],stage3_3[19]}
   );
   gpc615_5 gpc1683 (
      {stage2_3[58], stage2_3[59], stage2_3[60], stage2_3[61], stage2_3[62]},
      {stage2_4[44]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[10],stage3_5[16],stage3_4[20],stage3_3[20]}
   );
   gpc615_5 gpc1684 (
      {stage2_3[63], stage2_3[64], stage2_3[65], stage2_3[66], stage2_3[67]},
      {stage2_4[45]},
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage3_7[4],stage3_6[11],stage3_5[17],stage3_4[21],stage3_3[21]}
   );
   gpc615_5 gpc1685 (
      {stage2_3[68], stage2_3[69], stage2_3[70], stage2_3[71], stage2_3[72]},
      {stage2_4[46]},
      {stage2_5[30], stage2_5[31], stage2_5[32], stage2_5[33], stage2_5[34], stage2_5[35]},
      {stage3_7[5],stage3_6[12],stage3_5[18],stage3_4[22],stage3_3[22]}
   );
   gpc615_5 gpc1686 (
      {stage2_3[73], stage2_3[74], stage2_3[75], stage2_3[76], stage2_3[77]},
      {stage2_4[47]},
      {stage2_5[36], stage2_5[37], stage2_5[38], stage2_5[39], stage2_5[40], stage2_5[41]},
      {stage3_7[6],stage3_6[13],stage3_5[19],stage3_4[23],stage3_3[23]}
   );
   gpc615_5 gpc1687 (
      {stage2_3[78], stage2_3[79], stage2_3[80], stage2_3[81], stage2_3[82]},
      {stage2_4[48]},
      {stage2_5[42], stage2_5[43], stage2_5[44], stage2_5[45], stage2_5[46], stage2_5[47]},
      {stage3_7[7],stage3_6[14],stage3_5[20],stage3_4[24],stage3_3[24]}
   );
   gpc615_5 gpc1688 (
      {stage2_3[83], stage2_3[84], stage2_3[85], stage2_3[86], stage2_3[87]},
      {stage2_4[49]},
      {stage2_5[48], stage2_5[49], stage2_5[50], stage2_5[51], stage2_5[52], stage2_5[53]},
      {stage3_7[8],stage3_6[15],stage3_5[21],stage3_4[25],stage3_3[25]}
   );
   gpc615_5 gpc1689 (
      {stage2_3[88], stage2_3[89], stage2_3[90], stage2_3[91], stage2_3[92]},
      {stage2_4[50]},
      {stage2_5[54], stage2_5[55], stage2_5[56], stage2_5[57], stage2_5[58], stage2_5[59]},
      {stage3_7[9],stage3_6[16],stage3_5[22],stage3_4[26],stage3_3[26]}
   );
   gpc615_5 gpc1690 (
      {stage2_3[93], stage2_3[94], stage2_3[95], stage2_3[96], stage2_3[97]},
      {stage2_4[51]},
      {stage2_5[60], stage2_5[61], stage2_5[62], stage2_5[63], stage2_5[64], stage2_5[65]},
      {stage3_7[10],stage3_6[17],stage3_5[23],stage3_4[27],stage3_3[27]}
   );
   gpc615_5 gpc1691 (
      {stage2_3[98], stage2_3[99], stage2_3[100], stage2_3[101], stage2_3[102]},
      {stage2_4[52]},
      {stage2_5[66], stage2_5[67], stage2_5[68], stage2_5[69], stage2_5[70], stage2_5[71]},
      {stage3_7[11],stage3_6[18],stage3_5[24],stage3_4[28],stage3_3[28]}
   );
   gpc606_5 gpc1692 (
      {stage2_4[53], stage2_4[54], stage2_4[55], stage2_4[56], stage2_4[57], stage2_4[58]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[12],stage3_6[19],stage3_5[25],stage3_4[29]}
   );
   gpc606_5 gpc1693 (
      {stage2_4[59], stage2_4[60], stage2_4[61], stage2_4[62], stage2_4[63], stage2_4[64]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[13],stage3_6[20],stage3_5[26],stage3_4[30]}
   );
   gpc606_5 gpc1694 (
      {stage2_4[65], stage2_4[66], stage2_4[67], stage2_4[68], stage2_4[69], stage2_4[70]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[14],stage3_6[21],stage3_5[27],stage3_4[31]}
   );
   gpc606_5 gpc1695 (
      {stage2_4[71], stage2_4[72], stage2_4[73], stage2_4[74], stage2_4[75], stage2_4[76]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[15],stage3_6[22],stage3_5[28],stage3_4[32]}
   );
   gpc606_5 gpc1696 (
      {stage2_4[77], stage2_4[78], stage2_4[79], stage2_4[80], stage2_4[81], stage2_4[82]},
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28], stage2_6[29]},
      {stage3_8[4],stage3_7[16],stage3_6[23],stage3_5[29],stage3_4[33]}
   );
   gpc606_5 gpc1697 (
      {stage2_4[83], stage2_4[84], stage2_4[85], stage2_4[86], stage2_4[87], stage2_4[88]},
      {stage2_6[30], stage2_6[31], stage2_6[32], stage2_6[33], stage2_6[34], stage2_6[35]},
      {stage3_8[5],stage3_7[17],stage3_6[24],stage3_5[30],stage3_4[34]}
   );
   gpc606_5 gpc1698 (
      {stage2_4[89], stage2_4[90], stage2_4[91], stage2_4[92], stage2_4[93], stage2_4[94]},
      {stage2_6[36], stage2_6[37], stage2_6[38], stage2_6[39], stage2_6[40], stage2_6[41]},
      {stage3_8[6],stage3_7[18],stage3_6[25],stage3_5[31],stage3_4[35]}
   );
   gpc606_5 gpc1699 (
      {stage2_4[95], stage2_4[96], stage2_4[97], stage2_4[98], stage2_4[99], stage2_4[100]},
      {stage2_6[42], stage2_6[43], stage2_6[44], stage2_6[45], stage2_6[46], stage2_6[47]},
      {stage3_8[7],stage3_7[19],stage3_6[26],stage3_5[32],stage3_4[36]}
   );
   gpc606_5 gpc1700 (
      {stage2_4[101], stage2_4[102], stage2_4[103], stage2_4[104], stage2_4[105], stage2_4[106]},
      {stage2_6[48], stage2_6[49], stage2_6[50], stage2_6[51], stage2_6[52], stage2_6[53]},
      {stage3_8[8],stage3_7[20],stage3_6[27],stage3_5[33],stage3_4[37]}
   );
   gpc615_5 gpc1701 (
      {stage2_4[107], stage2_4[108], stage2_4[109], stage2_4[110], stage2_4[111]},
      {stage2_5[72]},
      {stage2_6[54], stage2_6[55], stage2_6[56], stage2_6[57], stage2_6[58], stage2_6[59]},
      {stage3_8[9],stage3_7[21],stage3_6[28],stage3_5[34],stage3_4[38]}
   );
   gpc615_5 gpc1702 (
      {stage2_4[112], stage2_4[113], stage2_4[114], stage2_4[115], stage2_4[116]},
      {stage2_5[73]},
      {stage2_6[60], stage2_6[61], stage2_6[62], stage2_6[63], stage2_6[64], stage2_6[65]},
      {stage3_8[10],stage3_7[22],stage3_6[29],stage3_5[35],stage3_4[39]}
   );
   gpc615_5 gpc1703 (
      {stage2_5[74], stage2_5[75], stage2_5[76], stage2_5[77], stage2_5[78]},
      {stage2_6[66]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[11],stage3_7[23],stage3_6[30],stage3_5[36]}
   );
   gpc615_5 gpc1704 (
      {stage2_5[79], stage2_5[80], stage2_5[81], stage2_5[82], stage2_5[83]},
      {stage2_6[67]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[12],stage3_7[24],stage3_6[31],stage3_5[37]}
   );
   gpc606_5 gpc1705 (
      {stage2_6[68], stage2_6[69], stage2_6[70], stage2_6[71], stage2_6[72], stage2_6[73]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[2],stage3_8[13],stage3_7[25],stage3_6[32]}
   );
   gpc606_5 gpc1706 (
      {stage2_6[74], stage2_6[75], stage2_6[76], stage2_6[77], stage2_6[78], stage2_6[79]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[3],stage3_8[14],stage3_7[26],stage3_6[33]}
   );
   gpc606_5 gpc1707 (
      {stage2_6[80], stage2_6[81], stage2_6[82], stage2_6[83], stage2_6[84], stage2_6[85]},
      {stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15], stage2_8[16], stage2_8[17]},
      {stage3_10[2],stage3_9[4],stage3_8[15],stage3_7[27],stage3_6[34]}
   );
   gpc606_5 gpc1708 (
      {stage2_6[86], stage2_6[87], stage2_6[88], stage2_6[89], stage2_6[90], stage2_6[91]},
      {stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21], stage2_8[22], stage2_8[23]},
      {stage3_10[3],stage3_9[5],stage3_8[16],stage3_7[28],stage3_6[35]}
   );
   gpc606_5 gpc1709 (
      {stage2_6[92], stage2_6[93], stage2_6[94], stage2_6[95], stage2_6[96], stage2_6[97]},
      {stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29]},
      {stage3_10[4],stage3_9[6],stage3_8[17],stage3_7[29],stage3_6[36]}
   );
   gpc606_5 gpc1710 (
      {stage2_6[98], stage2_6[99], stage2_6[100], stage2_6[101], stage2_6[102], stage2_6[103]},
      {stage2_8[30], stage2_8[31], stage2_8[32], stage2_8[33], stage2_8[34], stage2_8[35]},
      {stage3_10[5],stage3_9[7],stage3_8[18],stage3_7[30],stage3_6[37]}
   );
   gpc615_5 gpc1711 (
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16]},
      {stage2_8[36]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[6],stage3_9[8],stage3_8[19],stage3_7[31]}
   );
   gpc615_5 gpc1712 (
      {stage2_7[17], stage2_7[18], stage2_7[19], stage2_7[20], stage2_7[21]},
      {stage2_8[37]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[7],stage3_9[9],stage3_8[20],stage3_7[32]}
   );
   gpc615_5 gpc1713 (
      {stage2_7[22], stage2_7[23], stage2_7[24], stage2_7[25], stage2_7[26]},
      {stage2_8[38]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[8],stage3_9[10],stage3_8[21],stage3_7[33]}
   );
   gpc615_5 gpc1714 (
      {stage2_7[27], stage2_7[28], stage2_7[29], stage2_7[30], stage2_7[31]},
      {stage2_8[39]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[9],stage3_9[11],stage3_8[22],stage3_7[34]}
   );
   gpc615_5 gpc1715 (
      {stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36]},
      {stage2_8[40]},
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage3_11[4],stage3_10[10],stage3_9[12],stage3_8[23],stage3_7[35]}
   );
   gpc615_5 gpc1716 (
      {stage2_7[37], stage2_7[38], stage2_7[39], stage2_7[40], stage2_7[41]},
      {stage2_8[41]},
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage3_11[5],stage3_10[11],stage3_9[13],stage3_8[24],stage3_7[36]}
   );
   gpc615_5 gpc1717 (
      {stage2_7[42], stage2_7[43], stage2_7[44], stage2_7[45], stage2_7[46]},
      {stage2_8[42]},
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage3_11[6],stage3_10[12],stage3_9[14],stage3_8[25],stage3_7[37]}
   );
   gpc615_5 gpc1718 (
      {stage2_7[47], stage2_7[48], stage2_7[49], stage2_7[50], stage2_7[51]},
      {stage2_8[43]},
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46], stage2_9[47]},
      {stage3_11[7],stage3_10[13],stage3_9[15],stage3_8[26],stage3_7[38]}
   );
   gpc615_5 gpc1719 (
      {stage2_7[52], stage2_7[53], stage2_7[54], stage2_7[55], stage2_7[56]},
      {stage2_8[44]},
      {stage2_9[48], stage2_9[49], stage2_9[50], stage2_9[51], stage2_9[52], stage2_9[53]},
      {stage3_11[8],stage3_10[14],stage3_9[16],stage3_8[27],stage3_7[39]}
   );
   gpc615_5 gpc1720 (
      {stage2_7[57], stage2_7[58], stage2_7[59], stage2_7[60], stage2_7[61]},
      {stage2_8[45]},
      {stage2_9[54], stage2_9[55], stage2_9[56], stage2_9[57], stage2_9[58], stage2_9[59]},
      {stage3_11[9],stage3_10[15],stage3_9[17],stage3_8[28],stage3_7[40]}
   );
   gpc615_5 gpc1721 (
      {stage2_7[62], stage2_7[63], stage2_7[64], stage2_7[65], stage2_7[66]},
      {stage2_8[46]},
      {stage2_9[60], stage2_9[61], stage2_9[62], stage2_9[63], stage2_9[64], stage2_9[65]},
      {stage3_11[10],stage3_10[16],stage3_9[18],stage3_8[29],stage3_7[41]}
   );
   gpc615_5 gpc1722 (
      {stage2_7[67], stage2_7[68], stage2_7[69], stage2_7[70], stage2_7[71]},
      {stage2_8[47]},
      {stage2_9[66], stage2_9[67], stage2_9[68], stage2_9[69], stage2_9[70], stage2_9[71]},
      {stage3_11[11],stage3_10[17],stage3_9[19],stage3_8[30],stage3_7[42]}
   );
   gpc615_5 gpc1723 (
      {stage2_7[72], stage2_7[73], stage2_7[74], stage2_7[75], stage2_7[76]},
      {stage2_8[48]},
      {stage2_9[72], stage2_9[73], stage2_9[74], stage2_9[75], stage2_9[76], stage2_9[77]},
      {stage3_11[12],stage3_10[18],stage3_9[20],stage3_8[31],stage3_7[43]}
   );
   gpc615_5 gpc1724 (
      {stage2_7[77], stage2_7[78], stage2_7[79], stage2_7[80], stage2_7[81]},
      {stage2_8[49]},
      {stage2_9[78], stage2_9[79], stage2_9[80], stage2_9[81], stage2_9[82], stage2_9[83]},
      {stage3_11[13],stage3_10[19],stage3_9[21],stage3_8[32],stage3_7[44]}
   );
   gpc615_5 gpc1725 (
      {stage2_7[82], stage2_7[83], stage2_7[84], 1'b0, 1'b0},
      {stage2_8[50]},
      {stage2_9[84], stage2_9[85], stage2_9[86], stage2_9[87], stage2_9[88], stage2_9[89]},
      {stage3_11[14],stage3_10[20],stage3_9[22],stage3_8[33],stage3_7[45]}
   );
   gpc606_5 gpc1726 (
      {stage2_8[51], stage2_8[52], stage2_8[53], stage2_8[54], stage2_8[55], stage2_8[56]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[15],stage3_10[21],stage3_9[23],stage3_8[34]}
   );
   gpc615_5 gpc1727 (
      {stage2_8[57], stage2_8[58], stage2_8[59], stage2_8[60], stage2_8[61]},
      {stage2_9[90]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[16],stage3_10[22],stage3_9[24],stage3_8[35]}
   );
   gpc615_5 gpc1728 (
      {stage2_8[62], stage2_8[63], stage2_8[64], stage2_8[65], stage2_8[66]},
      {stage2_9[91]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[17],stage3_10[23],stage3_9[25],stage3_8[36]}
   );
   gpc615_5 gpc1729 (
      {stage2_8[67], stage2_8[68], stage2_8[69], stage2_8[70], stage2_8[71]},
      {stage2_9[92]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[18],stage3_10[24],stage3_9[26],stage3_8[37]}
   );
   gpc615_5 gpc1730 (
      {stage2_8[72], stage2_8[73], stage2_8[74], stage2_8[75], stage2_8[76]},
      {stage2_9[93]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[19],stage3_10[25],stage3_9[27],stage3_8[38]}
   );
   gpc615_5 gpc1731 (
      {stage2_8[77], stage2_8[78], stage2_8[79], stage2_8[80], stage2_8[81]},
      {stage2_9[94]},
      {stage2_10[30], stage2_10[31], stage2_10[32], stage2_10[33], stage2_10[34], stage2_10[35]},
      {stage3_12[5],stage3_11[20],stage3_10[26],stage3_9[28],stage3_8[39]}
   );
   gpc615_5 gpc1732 (
      {stage2_8[82], stage2_8[83], stage2_8[84], stage2_8[85], stage2_8[86]},
      {stage2_9[95]},
      {stage2_10[36], stage2_10[37], stage2_10[38], stage2_10[39], stage2_10[40], stage2_10[41]},
      {stage3_12[6],stage3_11[21],stage3_10[27],stage3_9[29],stage3_8[40]}
   );
   gpc606_5 gpc1733 (
      {stage2_9[96], stage2_9[97], stage2_9[98], stage2_9[99], stage2_9[100], stage2_9[101]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[7],stage3_11[22],stage3_10[28],stage3_9[30]}
   );
   gpc606_5 gpc1734 (
      {stage2_9[102], stage2_9[103], stage2_9[104], stage2_9[105], stage2_9[106], stage2_9[107]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[8],stage3_11[23],stage3_10[29],stage3_9[31]}
   );
   gpc606_5 gpc1735 (
      {stage2_9[108], stage2_9[109], stage2_9[110], stage2_9[111], stage2_9[112], stage2_9[113]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[9],stage3_11[24],stage3_10[30],stage3_9[32]}
   );
   gpc606_5 gpc1736 (
      {stage2_9[114], stage2_9[115], stage2_9[116], stage2_9[117], stage2_9[118], stage2_9[119]},
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage3_13[3],stage3_12[10],stage3_11[25],stage3_10[31],stage3_9[33]}
   );
   gpc615_5 gpc1737 (
      {stage2_10[42], stage2_10[43], stage2_10[44], stage2_10[45], stage2_10[46]},
      {stage2_11[24]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[4],stage3_12[11],stage3_11[26],stage3_10[32]}
   );
   gpc615_5 gpc1738 (
      {stage2_10[47], stage2_10[48], stage2_10[49], stage2_10[50], stage2_10[51]},
      {stage2_11[25]},
      {stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11]},
      {stage3_14[1],stage3_13[5],stage3_12[12],stage3_11[27],stage3_10[33]}
   );
   gpc615_5 gpc1739 (
      {stage2_10[52], stage2_10[53], stage2_10[54], stage2_10[55], stage2_10[56]},
      {stage2_11[26]},
      {stage2_12[12], stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17]},
      {stage3_14[2],stage3_13[6],stage3_12[13],stage3_11[28],stage3_10[34]}
   );
   gpc606_5 gpc1740 (
      {stage2_11[27], stage2_11[28], stage2_11[29], stage2_11[30], stage2_11[31], stage2_11[32]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[3],stage3_13[7],stage3_12[14],stage3_11[29]}
   );
   gpc606_5 gpc1741 (
      {stage2_11[33], stage2_11[34], stage2_11[35], stage2_11[36], stage2_11[37], stage2_11[38]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[4],stage3_13[8],stage3_12[15],stage3_11[30]}
   );
   gpc606_5 gpc1742 (
      {stage2_11[39], stage2_11[40], stage2_11[41], stage2_11[42], stage2_11[43], stage2_11[44]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[5],stage3_13[9],stage3_12[16],stage3_11[31]}
   );
   gpc606_5 gpc1743 (
      {stage2_11[45], stage2_11[46], stage2_11[47], stage2_11[48], stage2_11[49], stage2_11[50]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[6],stage3_13[10],stage3_12[17],stage3_11[32]}
   );
   gpc606_5 gpc1744 (
      {stage2_11[51], stage2_11[52], stage2_11[53], stage2_11[54], stage2_11[55], stage2_11[56]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[7],stage3_13[11],stage3_12[18],stage3_11[33]}
   );
   gpc606_5 gpc1745 (
      {stage2_11[57], stage2_11[58], stage2_11[59], stage2_11[60], stage2_11[61], stage2_11[62]},
      {stage2_13[30], stage2_13[31], stage2_13[32], stage2_13[33], stage2_13[34], stage2_13[35]},
      {stage3_15[5],stage3_14[8],stage3_13[12],stage3_12[19],stage3_11[34]}
   );
   gpc606_5 gpc1746 (
      {stage2_11[63], stage2_11[64], stage2_11[65], stage2_11[66], stage2_11[67], stage2_11[68]},
      {stage2_13[36], stage2_13[37], stage2_13[38], stage2_13[39], stage2_13[40], stage2_13[41]},
      {stage3_15[6],stage3_14[9],stage3_13[13],stage3_12[20],stage3_11[35]}
   );
   gpc606_5 gpc1747 (
      {stage2_11[69], stage2_11[70], stage2_11[71], stage2_11[72], stage2_11[73], stage2_11[74]},
      {stage2_13[42], stage2_13[43], stage2_13[44], stage2_13[45], stage2_13[46], stage2_13[47]},
      {stage3_15[7],stage3_14[10],stage3_13[14],stage3_12[21],stage3_11[36]}
   );
   gpc606_5 gpc1748 (
      {stage2_11[75], stage2_11[76], stage2_11[77], stage2_11[78], stage2_11[79], stage2_11[80]},
      {stage2_13[48], stage2_13[49], stage2_13[50], stage2_13[51], stage2_13[52], stage2_13[53]},
      {stage3_15[8],stage3_14[11],stage3_13[15],stage3_12[22],stage3_11[37]}
   );
   gpc606_5 gpc1749 (
      {stage2_11[81], stage2_11[82], stage2_11[83], stage2_11[84], stage2_11[85], stage2_11[86]},
      {stage2_13[54], stage2_13[55], stage2_13[56], stage2_13[57], stage2_13[58], stage2_13[59]},
      {stage3_15[9],stage3_14[12],stage3_13[16],stage3_12[23],stage3_11[38]}
   );
   gpc606_5 gpc1750 (
      {stage2_11[87], stage2_11[88], stage2_11[89], stage2_11[90], stage2_11[91], stage2_11[92]},
      {stage2_13[60], stage2_13[61], stage2_13[62], stage2_13[63], stage2_13[64], stage2_13[65]},
      {stage3_15[10],stage3_14[13],stage3_13[17],stage3_12[24],stage3_11[39]}
   );
   gpc606_5 gpc1751 (
      {stage2_11[93], stage2_11[94], stage2_11[95], stage2_11[96], stage2_11[97], stage2_11[98]},
      {stage2_13[66], stage2_13[67], stage2_13[68], stage2_13[69], stage2_13[70], stage2_13[71]},
      {stage3_15[11],stage3_14[14],stage3_13[18],stage3_12[25],stage3_11[40]}
   );
   gpc606_5 gpc1752 (
      {stage2_11[99], stage2_11[100], stage2_11[101], stage2_11[102], stage2_11[103], stage2_11[104]},
      {stage2_13[72], stage2_13[73], stage2_13[74], stage2_13[75], stage2_13[76], stage2_13[77]},
      {stage3_15[12],stage3_14[15],stage3_13[19],stage3_12[26],stage3_11[41]}
   );
   gpc606_5 gpc1753 (
      {stage2_11[105], stage2_11[106], stage2_11[107], stage2_11[108], stage2_11[109], stage2_11[110]},
      {stage2_13[78], stage2_13[79], stage2_13[80], stage2_13[81], stage2_13[82], stage2_13[83]},
      {stage3_15[13],stage3_14[16],stage3_13[20],stage3_12[27],stage3_11[42]}
   );
   gpc606_5 gpc1754 (
      {stage2_11[111], stage2_11[112], stage2_11[113], stage2_11[114], stage2_11[115], stage2_11[116]},
      {stage2_13[84], stage2_13[85], stage2_13[86], stage2_13[87], stage2_13[88], stage2_13[89]},
      {stage3_15[14],stage3_14[17],stage3_13[21],stage3_12[28],stage3_11[43]}
   );
   gpc606_5 gpc1755 (
      {stage2_11[117], stage2_11[118], stage2_11[119], stage2_11[120], stage2_11[121], stage2_11[122]},
      {stage2_13[90], stage2_13[91], stage2_13[92], stage2_13[93], stage2_13[94], stage2_13[95]},
      {stage3_15[15],stage3_14[18],stage3_13[22],stage3_12[29],stage3_11[44]}
   );
   gpc606_5 gpc1756 (
      {stage2_11[123], stage2_11[124], stage2_11[125], stage2_11[126], stage2_11[127], stage2_11[128]},
      {stage2_13[96], stage2_13[97], stage2_13[98], stage2_13[99], stage2_13[100], stage2_13[101]},
      {stage3_15[16],stage3_14[19],stage3_13[23],stage3_12[30],stage3_11[45]}
   );
   gpc606_5 gpc1757 (
      {stage2_12[18], stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[17],stage3_14[20],stage3_13[24],stage3_12[31]}
   );
   gpc606_5 gpc1758 (
      {stage2_12[24], stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[18],stage3_14[21],stage3_13[25],stage3_12[32]}
   );
   gpc606_5 gpc1759 (
      {stage2_12[30], stage2_12[31], stage2_12[32], stage2_12[33], stage2_12[34], stage2_12[35]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[19],stage3_14[22],stage3_13[26],stage3_12[33]}
   );
   gpc606_5 gpc1760 (
      {stage2_12[36], stage2_12[37], stage2_12[38], stage2_12[39], stage2_12[40], stage2_12[41]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[20],stage3_14[23],stage3_13[27],stage3_12[34]}
   );
   gpc606_5 gpc1761 (
      {stage2_12[42], stage2_12[43], stage2_12[44], stage2_12[45], stage2_12[46], stage2_12[47]},
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage3_16[4],stage3_15[21],stage3_14[24],stage3_13[28],stage3_12[35]}
   );
   gpc606_5 gpc1762 (
      {stage2_12[48], stage2_12[49], stage2_12[50], stage2_12[51], stage2_12[52], stage2_12[53]},
      {stage2_14[30], stage2_14[31], stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35]},
      {stage3_16[5],stage3_15[22],stage3_14[25],stage3_13[29],stage3_12[36]}
   );
   gpc606_5 gpc1763 (
      {stage2_12[54], stage2_12[55], stage2_12[56], stage2_12[57], stage2_12[58], stage2_12[59]},
      {stage2_14[36], stage2_14[37], stage2_14[38], stage2_14[39], stage2_14[40], stage2_14[41]},
      {stage3_16[6],stage3_15[23],stage3_14[26],stage3_13[30],stage3_12[37]}
   );
   gpc606_5 gpc1764 (
      {stage2_12[60], stage2_12[61], stage2_12[62], stage2_12[63], stage2_12[64], stage2_12[65]},
      {stage2_14[42], stage2_14[43], stage2_14[44], stage2_14[45], stage2_14[46], stage2_14[47]},
      {stage3_16[7],stage3_15[24],stage3_14[27],stage3_13[31],stage3_12[38]}
   );
   gpc606_5 gpc1765 (
      {stage2_12[66], stage2_12[67], stage2_12[68], stage2_12[69], stage2_12[70], stage2_12[71]},
      {stage2_14[48], stage2_14[49], stage2_14[50], stage2_14[51], stage2_14[52], stage2_14[53]},
      {stage3_16[8],stage3_15[25],stage3_14[28],stage3_13[32],stage3_12[39]}
   );
   gpc606_5 gpc1766 (
      {stage2_13[102], stage2_13[103], stage2_13[104], stage2_13[105], stage2_13[106], stage2_13[107]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[9],stage3_15[26],stage3_14[29],stage3_13[33]}
   );
   gpc606_5 gpc1767 (
      {stage2_13[108], stage2_13[109], stage2_13[110], stage2_13[111], stage2_13[112], stage2_13[113]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[10],stage3_15[27],stage3_14[30],stage3_13[34]}
   );
   gpc606_5 gpc1768 (
      {stage2_13[114], stage2_13[115], stage2_13[116], stage2_13[117], stage2_13[118], stage2_13[119]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[11],stage3_15[28],stage3_14[31],stage3_13[35]}
   );
   gpc606_5 gpc1769 (
      {stage2_13[120], stage2_13[121], stage2_13[122], stage2_13[123], stage2_13[124], stage2_13[125]},
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22], stage2_15[23]},
      {stage3_17[3],stage3_16[12],stage3_15[29],stage3_14[32],stage3_13[36]}
   );
   gpc606_5 gpc1770 (
      {stage2_13[126], stage2_13[127], stage2_13[128], stage2_13[129], stage2_13[130], stage2_13[131]},
      {stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27], stage2_15[28], stage2_15[29]},
      {stage3_17[4],stage3_16[13],stage3_15[30],stage3_14[33],stage3_13[37]}
   );
   gpc606_5 gpc1771 (
      {stage2_13[132], stage2_13[133], stage2_13[134], stage2_13[135], stage2_13[136], stage2_13[137]},
      {stage2_15[30], stage2_15[31], stage2_15[32], stage2_15[33], stage2_15[34], stage2_15[35]},
      {stage3_17[5],stage3_16[14],stage3_15[31],stage3_14[34],stage3_13[38]}
   );
   gpc606_5 gpc1772 (
      {stage2_14[54], stage2_14[55], stage2_14[56], stage2_14[57], stage2_14[58], stage2_14[59]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[6],stage3_16[15],stage3_15[32],stage3_14[35]}
   );
   gpc606_5 gpc1773 (
      {stage2_14[60], stage2_14[61], stage2_14[62], stage2_14[63], stage2_14[64], stage2_14[65]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[7],stage3_16[16],stage3_15[33],stage3_14[36]}
   );
   gpc606_5 gpc1774 (
      {stage2_14[66], stage2_14[67], stage2_14[68], stage2_14[69], stage2_14[70], stage2_14[71]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[8],stage3_16[17],stage3_15[34],stage3_14[37]}
   );
   gpc606_5 gpc1775 (
      {stage2_14[72], stage2_14[73], stage2_14[74], stage2_14[75], stage2_14[76], stage2_14[77]},
      {stage2_16[18], stage2_16[19], stage2_16[20], stage2_16[21], stage2_16[22], stage2_16[23]},
      {stage3_18[3],stage3_17[9],stage3_16[18],stage3_15[35],stage3_14[38]}
   );
   gpc606_5 gpc1776 (
      {stage2_14[78], stage2_14[79], stage2_14[80], stage2_14[81], stage2_14[82], stage2_14[83]},
      {stage2_16[24], stage2_16[25], stage2_16[26], stage2_16[27], stage2_16[28], stage2_16[29]},
      {stage3_18[4],stage3_17[10],stage3_16[19],stage3_15[36],stage3_14[39]}
   );
   gpc606_5 gpc1777 (
      {stage2_14[84], stage2_14[85], stage2_14[86], stage2_14[87], stage2_14[88], stage2_14[89]},
      {stage2_16[30], stage2_16[31], stage2_16[32], stage2_16[33], stage2_16[34], stage2_16[35]},
      {stage3_18[5],stage3_17[11],stage3_16[20],stage3_15[37],stage3_14[40]}
   );
   gpc606_5 gpc1778 (
      {stage2_14[90], stage2_14[91], stage2_14[92], stage2_14[93], stage2_14[94], stage2_14[95]},
      {stage2_16[36], stage2_16[37], stage2_16[38], stage2_16[39], stage2_16[40], stage2_16[41]},
      {stage3_18[6],stage3_17[12],stage3_16[21],stage3_15[38],stage3_14[41]}
   );
   gpc606_5 gpc1779 (
      {stage2_14[96], stage2_14[97], stage2_14[98], stage2_14[99], stage2_14[100], stage2_14[101]},
      {stage2_16[42], stage2_16[43], stage2_16[44], stage2_16[45], stage2_16[46], stage2_16[47]},
      {stage3_18[7],stage3_17[13],stage3_16[22],stage3_15[39],stage3_14[42]}
   );
   gpc615_5 gpc1780 (
      {stage2_14[102], stage2_14[103], stage2_14[104], stage2_14[105], stage2_14[106]},
      {stage2_15[36]},
      {stage2_16[48], stage2_16[49], stage2_16[50], stage2_16[51], stage2_16[52], stage2_16[53]},
      {stage3_18[8],stage3_17[14],stage3_16[23],stage3_15[40],stage3_14[43]}
   );
   gpc615_5 gpc1781 (
      {stage2_14[107], stage2_14[108], stage2_14[109], stage2_14[110], stage2_14[111]},
      {stage2_15[37]},
      {stage2_16[54], stage2_16[55], stage2_16[56], stage2_16[57], stage2_16[58], stage2_16[59]},
      {stage3_18[9],stage3_17[15],stage3_16[24],stage3_15[41],stage3_14[44]}
   );
   gpc615_5 gpc1782 (
      {stage2_15[38], stage2_15[39], stage2_15[40], stage2_15[41], stage2_15[42]},
      {stage2_16[60]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[10],stage3_17[16],stage3_16[25],stage3_15[42]}
   );
   gpc615_5 gpc1783 (
      {stage2_15[43], stage2_15[44], stage2_15[45], stage2_15[46], stage2_15[47]},
      {stage2_16[61]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[11],stage3_17[17],stage3_16[26],stage3_15[43]}
   );
   gpc615_5 gpc1784 (
      {stage2_15[48], stage2_15[49], stage2_15[50], stage2_15[51], stage2_15[52]},
      {stage2_16[62]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[12],stage3_17[18],stage3_16[27],stage3_15[44]}
   );
   gpc615_5 gpc1785 (
      {stage2_15[53], stage2_15[54], stage2_15[55], stage2_15[56], stage2_15[57]},
      {stage2_16[63]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[13],stage3_17[19],stage3_16[28],stage3_15[45]}
   );
   gpc615_5 gpc1786 (
      {stage2_15[58], stage2_15[59], stage2_15[60], stage2_15[61], stage2_15[62]},
      {stage2_16[64]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[14],stage3_17[20],stage3_16[29],stage3_15[46]}
   );
   gpc615_5 gpc1787 (
      {stage2_15[63], stage2_15[64], stage2_15[65], stage2_15[66], stage2_15[67]},
      {stage2_16[65]},
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], stage2_17[35]},
      {stage3_19[5],stage3_18[15],stage3_17[21],stage3_16[30],stage3_15[47]}
   );
   gpc615_5 gpc1788 (
      {stage2_15[68], stage2_15[69], stage2_15[70], stage2_15[71], stage2_15[72]},
      {stage2_16[66]},
      {stage2_17[36], stage2_17[37], stage2_17[38], stage2_17[39], stage2_17[40], stage2_17[41]},
      {stage3_19[6],stage3_18[16],stage3_17[22],stage3_16[31],stage3_15[48]}
   );
   gpc615_5 gpc1789 (
      {stage2_15[73], stage2_15[74], stage2_15[75], stage2_15[76], stage2_15[77]},
      {stage2_16[67]},
      {stage2_17[42], stage2_17[43], stage2_17[44], stage2_17[45], stage2_17[46], stage2_17[47]},
      {stage3_19[7],stage3_18[17],stage3_17[23],stage3_16[32],stage3_15[49]}
   );
   gpc606_5 gpc1790 (
      {stage2_16[68], stage2_16[69], stage2_16[70], stage2_16[71], stage2_16[72], stage2_16[73]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[8],stage3_18[18],stage3_17[24],stage3_16[33]}
   );
   gpc606_5 gpc1791 (
      {stage2_16[74], stage2_16[75], stage2_16[76], stage2_16[77], stage2_16[78], stage2_16[79]},
      {stage2_18[6], stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11]},
      {stage3_20[1],stage3_19[9],stage3_18[19],stage3_17[25],stage3_16[34]}
   );
   gpc606_5 gpc1792 (
      {stage2_16[80], stage2_16[81], stage2_16[82], stage2_16[83], stage2_16[84], stage2_16[85]},
      {stage2_18[12], stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17]},
      {stage3_20[2],stage3_19[10],stage3_18[20],stage3_17[26],stage3_16[35]}
   );
   gpc606_5 gpc1793 (
      {stage2_16[86], stage2_16[87], stage2_16[88], stage2_16[89], stage2_16[90], stage2_16[91]},
      {stage2_18[18], stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23]},
      {stage3_20[3],stage3_19[11],stage3_18[21],stage3_17[27],stage3_16[36]}
   );
   gpc606_5 gpc1794 (
      {stage2_17[48], stage2_17[49], stage2_17[50], stage2_17[51], stage2_17[52], stage2_17[53]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[4],stage3_19[12],stage3_18[22],stage3_17[28]}
   );
   gpc606_5 gpc1795 (
      {stage2_17[54], stage2_17[55], stage2_17[56], stage2_17[57], stage2_17[58], stage2_17[59]},
      {stage2_19[6], stage2_19[7], stage2_19[8], stage2_19[9], stage2_19[10], 1'b0},
      {stage3_21[1],stage3_20[5],stage3_19[13],stage3_18[23],stage3_17[29]}
   );
   gpc1_1 gpc1796 (
      {stage2_0[21]},
      {stage3_0[4]}
   );
   gpc1_1 gpc1797 (
      {stage2_0[22]},
      {stage3_0[5]}
   );
   gpc1_1 gpc1798 (
      {stage2_1[39]},
      {stage3_1[10]}
   );
   gpc1_1 gpc1799 (
      {stage2_1[40]},
      {stage3_1[11]}
   );
   gpc1_1 gpc1800 (
      {stage2_5[84]},
      {stage3_5[38]}
   );
   gpc1_1 gpc1801 (
      {stage2_5[85]},
      {stage3_5[39]}
   );
   gpc1_1 gpc1802 (
      {stage2_5[86]},
      {stage3_5[40]}
   );
   gpc1_1 gpc1803 (
      {stage2_5[87]},
      {stage3_5[41]}
   );
   gpc1_1 gpc1804 (
      {stage2_5[88]},
      {stage3_5[42]}
   );
   gpc1_1 gpc1805 (
      {stage2_5[89]},
      {stage3_5[43]}
   );
   gpc1_1 gpc1806 (
      {stage2_5[90]},
      {stage3_5[44]}
   );
   gpc1_1 gpc1807 (
      {stage2_5[91]},
      {stage3_5[45]}
   );
   gpc1_1 gpc1808 (
      {stage2_5[92]},
      {stage3_5[46]}
   );
   gpc1_1 gpc1809 (
      {stage2_5[93]},
      {stage3_5[47]}
   );
   gpc1_1 gpc1810 (
      {stage2_9[120]},
      {stage3_9[34]}
   );
   gpc1_1 gpc1811 (
      {stage2_9[121]},
      {stage3_9[35]}
   );
   gpc1_1 gpc1812 (
      {stage2_9[122]},
      {stage3_9[36]}
   );
   gpc1_1 gpc1813 (
      {stage2_9[123]},
      {stage3_9[37]}
   );
   gpc1_1 gpc1814 (
      {stage2_9[124]},
      {stage3_9[38]}
   );
   gpc1_1 gpc1815 (
      {stage2_9[125]},
      {stage3_9[39]}
   );
   gpc1_1 gpc1816 (
      {stage2_9[126]},
      {stage3_9[40]}
   );
   gpc1_1 gpc1817 (
      {stage2_9[127]},
      {stage3_9[41]}
   );
   gpc1_1 gpc1818 (
      {stage2_9[128]},
      {stage3_9[42]}
   );
   gpc1_1 gpc1819 (
      {stage2_9[129]},
      {stage3_9[43]}
   );
   gpc1_1 gpc1820 (
      {stage2_9[130]},
      {stage3_9[44]}
   );
   gpc1_1 gpc1821 (
      {stage2_9[131]},
      {stage3_9[45]}
   );
   gpc1_1 gpc1822 (
      {stage2_9[132]},
      {stage3_9[46]}
   );
   gpc1_1 gpc1823 (
      {stage2_9[133]},
      {stage3_9[47]}
   );
   gpc1_1 gpc1824 (
      {stage2_9[134]},
      {stage3_9[48]}
   );
   gpc1_1 gpc1825 (
      {stage2_9[135]},
      {stage3_9[49]}
   );
   gpc1_1 gpc1826 (
      {stage2_9[136]},
      {stage3_9[50]}
   );
   gpc1_1 gpc1827 (
      {stage2_9[137]},
      {stage3_9[51]}
   );
   gpc1_1 gpc1828 (
      {stage2_10[57]},
      {stage3_10[35]}
   );
   gpc1_1 gpc1829 (
      {stage2_10[58]},
      {stage3_10[36]}
   );
   gpc1_1 gpc1830 (
      {stage2_10[59]},
      {stage3_10[37]}
   );
   gpc1_1 gpc1831 (
      {stage2_10[60]},
      {stage3_10[38]}
   );
   gpc1_1 gpc1832 (
      {stage2_10[61]},
      {stage3_10[39]}
   );
   gpc1_1 gpc1833 (
      {stage2_10[62]},
      {stage3_10[40]}
   );
   gpc1_1 gpc1834 (
      {stage2_10[63]},
      {stage3_10[41]}
   );
   gpc1_1 gpc1835 (
      {stage2_10[64]},
      {stage3_10[42]}
   );
   gpc1_1 gpc1836 (
      {stage2_10[65]},
      {stage3_10[43]}
   );
   gpc1_1 gpc1837 (
      {stage2_10[66]},
      {stage3_10[44]}
   );
   gpc1_1 gpc1838 (
      {stage2_10[67]},
      {stage3_10[45]}
   );
   gpc1_1 gpc1839 (
      {stage2_10[68]},
      {stage3_10[46]}
   );
   gpc1_1 gpc1840 (
      {stage2_10[69]},
      {stage3_10[47]}
   );
   gpc1_1 gpc1841 (
      {stage2_10[70]},
      {stage3_10[48]}
   );
   gpc1_1 gpc1842 (
      {stage2_10[71]},
      {stage3_10[49]}
   );
   gpc1_1 gpc1843 (
      {stage2_10[72]},
      {stage3_10[50]}
   );
   gpc1_1 gpc1844 (
      {stage2_10[73]},
      {stage3_10[51]}
   );
   gpc1_1 gpc1845 (
      {stage2_10[74]},
      {stage3_10[52]}
   );
   gpc1_1 gpc1846 (
      {stage2_10[75]},
      {stage3_10[53]}
   );
   gpc1_1 gpc1847 (
      {stage2_10[76]},
      {stage3_10[54]}
   );
   gpc1_1 gpc1848 (
      {stage2_10[77]},
      {stage3_10[55]}
   );
   gpc1_1 gpc1849 (
      {stage2_10[78]},
      {stage3_10[56]}
   );
   gpc1_1 gpc1850 (
      {stage2_10[79]},
      {stage3_10[57]}
   );
   gpc1_1 gpc1851 (
      {stage2_10[80]},
      {stage3_10[58]}
   );
   gpc1_1 gpc1852 (
      {stage2_10[81]},
      {stage3_10[59]}
   );
   gpc1_1 gpc1853 (
      {stage2_10[82]},
      {stage3_10[60]}
   );
   gpc1_1 gpc1854 (
      {stage2_10[83]},
      {stage3_10[61]}
   );
   gpc1_1 gpc1855 (
      {stage2_10[84]},
      {stage3_10[62]}
   );
   gpc1_1 gpc1856 (
      {stage2_10[85]},
      {stage3_10[63]}
   );
   gpc1_1 gpc1857 (
      {stage2_11[129]},
      {stage3_11[46]}
   );
   gpc1_1 gpc1858 (
      {stage2_11[130]},
      {stage3_11[47]}
   );
   gpc1_1 gpc1859 (
      {stage2_11[131]},
      {stage3_11[48]}
   );
   gpc1_1 gpc1860 (
      {stage2_11[132]},
      {stage3_11[49]}
   );
   gpc1_1 gpc1861 (
      {stage2_11[133]},
      {stage3_11[50]}
   );
   gpc1_1 gpc1862 (
      {stage2_11[134]},
      {stage3_11[51]}
   );
   gpc1_1 gpc1863 (
      {stage2_11[135]},
      {stage3_11[52]}
   );
   gpc1_1 gpc1864 (
      {stage2_11[136]},
      {stage3_11[53]}
   );
   gpc1_1 gpc1865 (
      {stage2_11[137]},
      {stage3_11[54]}
   );
   gpc1_1 gpc1866 (
      {stage2_11[138]},
      {stage3_11[55]}
   );
   gpc1_1 gpc1867 (
      {stage2_11[139]},
      {stage3_11[56]}
   );
   gpc1_1 gpc1868 (
      {stage2_11[140]},
      {stage3_11[57]}
   );
   gpc1_1 gpc1869 (
      {stage2_11[141]},
      {stage3_11[58]}
   );
   gpc1_1 gpc1870 (
      {stage2_11[142]},
      {stage3_11[59]}
   );
   gpc1_1 gpc1871 (
      {stage2_11[143]},
      {stage3_11[60]}
   );
   gpc1_1 gpc1872 (
      {stage2_12[72]},
      {stage3_12[40]}
   );
   gpc1_1 gpc1873 (
      {stage2_12[73]},
      {stage3_12[41]}
   );
   gpc1_1 gpc1874 (
      {stage2_12[74]},
      {stage3_12[42]}
   );
   gpc1_1 gpc1875 (
      {stage2_12[75]},
      {stage3_12[43]}
   );
   gpc1_1 gpc1876 (
      {stage2_12[76]},
      {stage3_12[44]}
   );
   gpc1_1 gpc1877 (
      {stage2_12[77]},
      {stage3_12[45]}
   );
   gpc1_1 gpc1878 (
      {stage2_12[78]},
      {stage3_12[46]}
   );
   gpc1_1 gpc1879 (
      {stage2_12[79]},
      {stage3_12[47]}
   );
   gpc1_1 gpc1880 (
      {stage2_12[80]},
      {stage3_12[48]}
   );
   gpc1_1 gpc1881 (
      {stage2_12[81]},
      {stage3_12[49]}
   );
   gpc1_1 gpc1882 (
      {stage2_12[82]},
      {stage3_12[50]}
   );
   gpc1_1 gpc1883 (
      {stage2_12[83]},
      {stage3_12[51]}
   );
   gpc1_1 gpc1884 (
      {stage2_12[84]},
      {stage3_12[52]}
   );
   gpc1_1 gpc1885 (
      {stage2_13[138]},
      {stage3_13[39]}
   );
   gpc1_1 gpc1886 (
      {stage2_13[139]},
      {stage3_13[40]}
   );
   gpc1_1 gpc1887 (
      {stage2_13[140]},
      {stage3_13[41]}
   );
   gpc1_1 gpc1888 (
      {stage2_14[112]},
      {stage3_14[45]}
   );
   gpc1_1 gpc1889 (
      {stage2_14[113]},
      {stage3_14[46]}
   );
   gpc1_1 gpc1890 (
      {stage2_14[114]},
      {stage3_14[47]}
   );
   gpc1_1 gpc1891 (
      {stage2_14[115]},
      {stage3_14[48]}
   );
   gpc1_1 gpc1892 (
      {stage2_14[116]},
      {stage3_14[49]}
   );
   gpc1_1 gpc1893 (
      {stage2_14[117]},
      {stage3_14[50]}
   );
   gpc1_1 gpc1894 (
      {stage2_14[118]},
      {stage3_14[51]}
   );
   gpc1_1 gpc1895 (
      {stage2_14[119]},
      {stage3_14[52]}
   );
   gpc1_1 gpc1896 (
      {stage2_14[120]},
      {stage3_14[53]}
   );
   gpc1_1 gpc1897 (
      {stage2_14[121]},
      {stage3_14[54]}
   );
   gpc1_1 gpc1898 (
      {stage2_14[122]},
      {stage3_14[55]}
   );
   gpc1_1 gpc1899 (
      {stage2_14[123]},
      {stage3_14[56]}
   );
   gpc1_1 gpc1900 (
      {stage2_14[124]},
      {stage3_14[57]}
   );
   gpc1_1 gpc1901 (
      {stage2_15[78]},
      {stage3_15[50]}
   );
   gpc1_1 gpc1902 (
      {stage2_15[79]},
      {stage3_15[51]}
   );
   gpc1_1 gpc1903 (
      {stage2_15[80]},
      {stage3_15[52]}
   );
   gpc1_1 gpc1904 (
      {stage2_15[81]},
      {stage3_15[53]}
   );
   gpc1_1 gpc1905 (
      {stage2_15[82]},
      {stage3_15[54]}
   );
   gpc1_1 gpc1906 (
      {stage2_15[83]},
      {stage3_15[55]}
   );
   gpc1_1 gpc1907 (
      {stage2_15[84]},
      {stage3_15[56]}
   );
   gpc1_1 gpc1908 (
      {stage2_16[92]},
      {stage3_16[37]}
   );
   gpc1_1 gpc1909 (
      {stage2_16[93]},
      {stage3_16[38]}
   );
   gpc1_1 gpc1910 (
      {stage2_16[94]},
      {stage3_16[39]}
   );
   gpc1_1 gpc1911 (
      {stage2_16[95]},
      {stage3_16[40]}
   );
   gpc1_1 gpc1912 (
      {stage2_16[96]},
      {stage3_16[41]}
   );
   gpc1_1 gpc1913 (
      {stage2_16[97]},
      {stage3_16[42]}
   );
   gpc1_1 gpc1914 (
      {stage2_16[98]},
      {stage3_16[43]}
   );
   gpc1_1 gpc1915 (
      {stage2_16[99]},
      {stage3_16[44]}
   );
   gpc1_1 gpc1916 (
      {stage2_16[100]},
      {stage3_16[45]}
   );
   gpc1_1 gpc1917 (
      {stage2_16[101]},
      {stage3_16[46]}
   );
   gpc1_1 gpc1918 (
      {stage2_16[102]},
      {stage3_16[47]}
   );
   gpc1_1 gpc1919 (
      {stage2_16[103]},
      {stage3_16[48]}
   );
   gpc1_1 gpc1920 (
      {stage2_16[104]},
      {stage3_16[49]}
   );
   gpc1_1 gpc1921 (
      {stage2_17[60]},
      {stage3_17[30]}
   );
   gpc1_1 gpc1922 (
      {stage2_17[61]},
      {stage3_17[31]}
   );
   gpc1_1 gpc1923 (
      {stage2_18[24]},
      {stage3_18[24]}
   );
   gpc1_1 gpc1924 (
      {stage2_18[25]},
      {stage3_18[25]}
   );
   gpc606_5 gpc1925 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5]},
      {stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0]}
   );
   gpc606_5 gpc1926 (
      {stage3_1[6], stage3_1[7], stage3_1[8], stage3_1[9], stage3_1[10], stage3_1[11]},
      {stage3_3[6], stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc615_5 gpc1927 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4]},
      {stage3_3[12]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[2],stage4_4[2],stage4_3[2],stage4_2[2]}
   );
   gpc615_5 gpc1928 (
      {stage3_2[5], stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9]},
      {stage3_3[13]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[3],stage4_4[3],stage4_3[3],stage4_2[3]}
   );
   gpc615_5 gpc1929 (
      {stage3_3[14], stage3_3[15], stage3_3[16], stage3_3[17], stage3_3[18]},
      {stage3_4[12]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[2],stage4_5[4],stage4_4[4],stage4_3[4]}
   );
   gpc615_5 gpc1930 (
      {stage3_3[19], stage3_3[20], stage3_3[21], stage3_3[22], stage3_3[23]},
      {stage3_4[13]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[3],stage4_5[5],stage4_4[5],stage4_3[5]}
   );
   gpc606_5 gpc1931 (
      {stage3_4[14], stage3_4[15], stage3_4[16], stage3_4[17], stage3_4[18], stage3_4[19]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[2],stage4_6[4],stage4_5[6],stage4_4[6]}
   );
   gpc615_5 gpc1932 (
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16]},
      {stage3_6[6]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage4_9[0],stage4_8[1],stage4_7[3],stage4_6[5],stage4_5[7]}
   );
   gpc615_5 gpc1933 (
      {stage3_5[17], stage3_5[18], stage3_5[19], stage3_5[20], stage3_5[21]},
      {stage3_6[7]},
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage4_9[1],stage4_8[2],stage4_7[4],stage4_6[6],stage4_5[8]}
   );
   gpc615_5 gpc1934 (
      {stage3_5[22], stage3_5[23], stage3_5[24], stage3_5[25], stage3_5[26]},
      {stage3_6[8]},
      {stage3_7[12], stage3_7[13], stage3_7[14], stage3_7[15], stage3_7[16], stage3_7[17]},
      {stage4_9[2],stage4_8[3],stage4_7[5],stage4_6[7],stage4_5[9]}
   );
   gpc615_5 gpc1935 (
      {stage3_5[27], stage3_5[28], stage3_5[29], stage3_5[30], stage3_5[31]},
      {stage3_6[9]},
      {stage3_7[18], stage3_7[19], stage3_7[20], stage3_7[21], stage3_7[22], stage3_7[23]},
      {stage4_9[3],stage4_8[4],stage4_7[6],stage4_6[8],stage4_5[10]}
   );
   gpc615_5 gpc1936 (
      {stage3_5[32], stage3_5[33], stage3_5[34], stage3_5[35], stage3_5[36]},
      {stage3_6[10]},
      {stage3_7[24], stage3_7[25], stage3_7[26], stage3_7[27], stage3_7[28], stage3_7[29]},
      {stage4_9[4],stage4_8[5],stage4_7[7],stage4_6[9],stage4_5[11]}
   );
   gpc615_5 gpc1937 (
      {stage3_5[37], stage3_5[38], stage3_5[39], stage3_5[40], stage3_5[41]},
      {stage3_6[11]},
      {stage3_7[30], stage3_7[31], stage3_7[32], stage3_7[33], stage3_7[34], stage3_7[35]},
      {stage4_9[5],stage4_8[6],stage4_7[8],stage4_6[10],stage4_5[12]}
   );
   gpc615_5 gpc1938 (
      {stage3_5[42], stage3_5[43], stage3_5[44], stage3_5[45], stage3_5[46]},
      {stage3_6[12]},
      {stage3_7[36], stage3_7[37], stage3_7[38], stage3_7[39], stage3_7[40], stage3_7[41]},
      {stage4_9[6],stage4_8[7],stage4_7[9],stage4_6[11],stage4_5[13]}
   );
   gpc606_5 gpc1939 (
      {stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17], stage3_6[18]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[7],stage4_8[8],stage4_7[10],stage4_6[12]}
   );
   gpc606_5 gpc1940 (
      {stage3_6[19], stage3_6[20], stage3_6[21], stage3_6[22], stage3_6[23], stage3_6[24]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[8],stage4_8[9],stage4_7[11],stage4_6[13]}
   );
   gpc606_5 gpc1941 (
      {stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28], stage3_6[29], stage3_6[30]},
      {stage3_8[12], stage3_8[13], stage3_8[14], stage3_8[15], stage3_8[16], stage3_8[17]},
      {stage4_10[2],stage4_9[9],stage4_8[10],stage4_7[12],stage4_6[14]}
   );
   gpc615_5 gpc1942 (
      {stage3_8[18], stage3_8[19], stage3_8[20], stage3_8[21], stage3_8[22]},
      {stage3_9[0]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[0],stage4_10[3],stage4_9[10],stage4_8[11]}
   );
   gpc615_5 gpc1943 (
      {stage3_8[23], stage3_8[24], stage3_8[25], stage3_8[26], stage3_8[27]},
      {stage3_9[1]},
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage4_12[1],stage4_11[1],stage4_10[4],stage4_9[11],stage4_8[12]}
   );
   gpc606_5 gpc1944 (
      {stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5], stage3_9[6], stage3_9[7]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[2],stage4_11[2],stage4_10[5],stage4_9[12]}
   );
   gpc615_5 gpc1945 (
      {stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11], stage3_9[12]},
      {stage3_10[12]},
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage4_13[1],stage4_12[3],stage4_11[3],stage4_10[6],stage4_9[13]}
   );
   gpc615_5 gpc1946 (
      {stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage3_10[13]},
      {stage3_11[12], stage3_11[13], stage3_11[14], stage3_11[15], stage3_11[16], stage3_11[17]},
      {stage4_13[2],stage4_12[4],stage4_11[4],stage4_10[7],stage4_9[14]}
   );
   gpc615_5 gpc1947 (
      {stage3_9[18], stage3_9[19], stage3_9[20], stage3_9[21], stage3_9[22]},
      {stage3_10[14]},
      {stage3_11[18], stage3_11[19], stage3_11[20], stage3_11[21], stage3_11[22], stage3_11[23]},
      {stage4_13[3],stage4_12[5],stage4_11[5],stage4_10[8],stage4_9[15]}
   );
   gpc615_5 gpc1948 (
      {stage3_9[23], stage3_9[24], stage3_9[25], stage3_9[26], stage3_9[27]},
      {stage3_10[15]},
      {stage3_11[24], stage3_11[25], stage3_11[26], stage3_11[27], stage3_11[28], stage3_11[29]},
      {stage4_13[4],stage4_12[6],stage4_11[6],stage4_10[9],stage4_9[16]}
   );
   gpc615_5 gpc1949 (
      {stage3_9[28], stage3_9[29], stage3_9[30], stage3_9[31], stage3_9[32]},
      {stage3_10[16]},
      {stage3_11[30], stage3_11[31], stage3_11[32], stage3_11[33], stage3_11[34], stage3_11[35]},
      {stage4_13[5],stage4_12[7],stage4_11[7],stage4_10[10],stage4_9[17]}
   );
   gpc615_5 gpc1950 (
      {stage3_9[33], stage3_9[34], stage3_9[35], stage3_9[36], stage3_9[37]},
      {stage3_10[17]},
      {stage3_11[36], stage3_11[37], stage3_11[38], stage3_11[39], stage3_11[40], stage3_11[41]},
      {stage4_13[6],stage4_12[8],stage4_11[8],stage4_10[11],stage4_9[18]}
   );
   gpc615_5 gpc1951 (
      {stage3_9[38], stage3_9[39], stage3_9[40], stage3_9[41], stage3_9[42]},
      {stage3_10[18]},
      {stage3_11[42], stage3_11[43], stage3_11[44], stage3_11[45], stage3_11[46], stage3_11[47]},
      {stage4_13[7],stage4_12[9],stage4_11[9],stage4_10[12],stage4_9[19]}
   );
   gpc615_5 gpc1952 (
      {stage3_9[43], stage3_9[44], stage3_9[45], stage3_9[46], stage3_9[47]},
      {stage3_10[19]},
      {stage3_11[48], stage3_11[49], stage3_11[50], stage3_11[51], stage3_11[52], stage3_11[53]},
      {stage4_13[8],stage4_12[10],stage4_11[10],stage4_10[13],stage4_9[20]}
   );
   gpc606_5 gpc1953 (
      {stage3_10[20], stage3_10[21], stage3_10[22], stage3_10[23], stage3_10[24], stage3_10[25]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[9],stage4_12[11],stage4_11[11],stage4_10[14]}
   );
   gpc606_5 gpc1954 (
      {stage3_10[26], stage3_10[27], stage3_10[28], stage3_10[29], stage3_10[30], stage3_10[31]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[10],stage4_12[12],stage4_11[12],stage4_10[15]}
   );
   gpc606_5 gpc1955 (
      {stage3_10[32], stage3_10[33], stage3_10[34], stage3_10[35], stage3_10[36], stage3_10[37]},
      {stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15], stage3_12[16], stage3_12[17]},
      {stage4_14[2],stage4_13[11],stage4_12[13],stage4_11[13],stage4_10[16]}
   );
   gpc606_5 gpc1956 (
      {stage3_10[38], stage3_10[39], stage3_10[40], stage3_10[41], stage3_10[42], stage3_10[43]},
      {stage3_12[18], stage3_12[19], stage3_12[20], stage3_12[21], stage3_12[22], stage3_12[23]},
      {stage4_14[3],stage4_13[12],stage4_12[14],stage4_11[14],stage4_10[17]}
   );
   gpc606_5 gpc1957 (
      {stage3_12[24], stage3_12[25], stage3_12[26], stage3_12[27], stage3_12[28], stage3_12[29]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[0],stage4_14[4],stage4_13[13],stage4_12[15]}
   );
   gpc606_5 gpc1958 (
      {stage3_12[30], stage3_12[31], stage3_12[32], stage3_12[33], stage3_12[34], stage3_12[35]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[1],stage4_14[5],stage4_13[14],stage4_12[16]}
   );
   gpc606_5 gpc1959 (
      {stage3_12[36], stage3_12[37], stage3_12[38], stage3_12[39], stage3_12[40], stage3_12[41]},
      {stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16], stage3_14[17]},
      {stage4_16[2],stage4_15[2],stage4_14[6],stage4_13[15],stage4_12[17]}
   );
   gpc606_5 gpc1960 (
      {stage3_12[42], stage3_12[43], stage3_12[44], stage3_12[45], stage3_12[46], stage3_12[47]},
      {stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21], stage3_14[22], stage3_14[23]},
      {stage4_16[3],stage4_15[3],stage4_14[7],stage4_13[16],stage4_12[18]}
   );
   gpc1163_5 gpc1961 (
      {stage3_13[0], stage3_13[1], stage3_13[2]},
      {stage3_14[24], stage3_14[25], stage3_14[26], stage3_14[27], stage3_14[28], stage3_14[29]},
      {stage3_15[0]},
      {stage3_16[0]},
      {stage4_17[0],stage4_16[4],stage4_15[4],stage4_14[8],stage4_13[17]}
   );
   gpc1163_5 gpc1962 (
      {stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage3_14[30], stage3_14[31], stage3_14[32], stage3_14[33], stage3_14[34], stage3_14[35]},
      {stage3_15[1]},
      {stage3_16[1]},
      {stage4_17[1],stage4_16[5],stage4_15[5],stage4_14[9],stage4_13[18]}
   );
   gpc1163_5 gpc1963 (
      {stage3_13[6], stage3_13[7], stage3_13[8]},
      {stage3_14[36], stage3_14[37], stage3_14[38], stage3_14[39], stage3_14[40], stage3_14[41]},
      {stage3_15[2]},
      {stage3_16[2]},
      {stage4_17[2],stage4_16[6],stage4_15[6],stage4_14[10],stage4_13[19]}
   );
   gpc1163_5 gpc1964 (
      {stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage3_14[42], stage3_14[43], stage3_14[44], stage3_14[45], stage3_14[46], stage3_14[47]},
      {stage3_15[3]},
      {stage3_16[3]},
      {stage4_17[3],stage4_16[7],stage4_15[7],stage4_14[11],stage4_13[20]}
   );
   gpc606_5 gpc1965 (
      {stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15], stage3_13[16], stage3_13[17]},
      {stage3_15[4], stage3_15[5], stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9]},
      {stage4_17[4],stage4_16[8],stage4_15[8],stage4_14[12],stage4_13[21]}
   );
   gpc606_5 gpc1966 (
      {stage3_13[18], stage3_13[19], stage3_13[20], stage3_13[21], stage3_13[22], stage3_13[23]},
      {stage3_15[10], stage3_15[11], stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15]},
      {stage4_17[5],stage4_16[9],stage4_15[9],stage4_14[13],stage4_13[22]}
   );
   gpc606_5 gpc1967 (
      {stage3_13[24], stage3_13[25], stage3_13[26], stage3_13[27], stage3_13[28], stage3_13[29]},
      {stage3_15[16], stage3_15[17], stage3_15[18], stage3_15[19], stage3_15[20], stage3_15[21]},
      {stage4_17[6],stage4_16[10],stage4_15[10],stage4_14[14],stage4_13[23]}
   );
   gpc606_5 gpc1968 (
      {stage3_13[30], stage3_13[31], stage3_13[32], stage3_13[33], stage3_13[34], stage3_13[35]},
      {stage3_15[22], stage3_15[23], stage3_15[24], stage3_15[25], stage3_15[26], stage3_15[27]},
      {stage4_17[7],stage4_16[11],stage4_15[11],stage4_14[15],stage4_13[24]}
   );
   gpc606_5 gpc1969 (
      {stage3_13[36], stage3_13[37], stage3_13[38], stage3_13[39], stage3_13[40], stage3_13[41]},
      {stage3_15[28], stage3_15[29], stage3_15[30], stage3_15[31], stage3_15[32], stage3_15[33]},
      {stage4_17[8],stage4_16[12],stage4_15[12],stage4_14[16],stage4_13[25]}
   );
   gpc615_5 gpc1970 (
      {stage3_14[48], stage3_14[49], stage3_14[50], stage3_14[51], stage3_14[52]},
      {stage3_15[34]},
      {stage3_16[4], stage3_16[5], stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9]},
      {stage4_18[0],stage4_17[9],stage4_16[13],stage4_15[13],stage4_14[17]}
   );
   gpc615_5 gpc1971 (
      {stage3_14[53], stage3_14[54], stage3_14[55], stage3_14[56], stage3_14[57]},
      {stage3_15[35]},
      {stage3_16[10], stage3_16[11], stage3_16[12], stage3_16[13], stage3_16[14], stage3_16[15]},
      {stage4_18[1],stage4_17[10],stage4_16[14],stage4_15[14],stage4_14[18]}
   );
   gpc606_5 gpc1972 (
      {stage3_15[36], stage3_15[37], stage3_15[38], stage3_15[39], stage3_15[40], stage3_15[41]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[2],stage4_17[11],stage4_16[15],stage4_15[15]}
   );
   gpc606_5 gpc1973 (
      {stage3_15[42], stage3_15[43], stage3_15[44], stage3_15[45], stage3_15[46], stage3_15[47]},
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage4_19[1],stage4_18[3],stage4_17[12],stage4_16[16],stage4_15[16]}
   );
   gpc615_5 gpc1974 (
      {stage3_15[48], stage3_15[49], stage3_15[50], stage3_15[51], stage3_15[52]},
      {stage3_16[16]},
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage4_19[2],stage4_18[4],stage4_17[13],stage4_16[17],stage4_15[17]}
   );
   gpc606_5 gpc1975 (
      {stage3_16[17], stage3_16[18], stage3_16[19], stage3_16[20], stage3_16[21], stage3_16[22]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[3],stage4_18[5],stage4_17[14],stage4_16[18]}
   );
   gpc606_5 gpc1976 (
      {stage3_16[23], stage3_16[24], stage3_16[25], stage3_16[26], stage3_16[27], stage3_16[28]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage4_20[1],stage4_19[4],stage4_18[6],stage4_17[15],stage4_16[19]}
   );
   gpc606_5 gpc1977 (
      {stage3_16[29], stage3_16[30], stage3_16[31], stage3_16[32], stage3_16[33], stage3_16[34]},
      {stage3_18[12], stage3_18[13], stage3_18[14], stage3_18[15], stage3_18[16], stage3_18[17]},
      {stage4_20[2],stage4_19[5],stage4_18[7],stage4_17[16],stage4_16[20]}
   );
   gpc606_5 gpc1978 (
      {stage3_16[35], stage3_16[36], stage3_16[37], stage3_16[38], stage3_16[39], stage3_16[40]},
      {stage3_18[18], stage3_18[19], stage3_18[20], stage3_18[21], stage3_18[22], stage3_18[23]},
      {stage4_20[3],stage4_19[6],stage4_18[8],stage4_17[17],stage4_16[21]}
   );
   gpc606_5 gpc1979 (
      {stage3_17[18], stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[4],stage4_19[7],stage4_18[9],stage4_17[18]}
   );
   gpc606_5 gpc1980 (
      {stage3_17[24], stage3_17[25], stage3_17[26], stage3_17[27], stage3_17[28], stage3_17[29]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage4_21[1],stage4_20[5],stage4_19[8],stage4_18[10],stage4_17[19]}
   );
   gpc1_1 gpc1981 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc1982 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc1983 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc1984 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc1985 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc1986 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc1987 (
      {stage3_2[10]},
      {stage4_2[4]}
   );
   gpc1_1 gpc1988 (
      {stage3_2[11]},
      {stage4_2[5]}
   );
   gpc1_1 gpc1989 (
      {stage3_2[12]},
      {stage4_2[6]}
   );
   gpc1_1 gpc1990 (
      {stage3_2[13]},
      {stage4_2[7]}
   );
   gpc1_1 gpc1991 (
      {stage3_2[14]},
      {stage4_2[8]}
   );
   gpc1_1 gpc1992 (
      {stage3_2[15]},
      {stage4_2[9]}
   );
   gpc1_1 gpc1993 (
      {stage3_2[16]},
      {stage4_2[10]}
   );
   gpc1_1 gpc1994 (
      {stage3_3[24]},
      {stage4_3[6]}
   );
   gpc1_1 gpc1995 (
      {stage3_3[25]},
      {stage4_3[7]}
   );
   gpc1_1 gpc1996 (
      {stage3_3[26]},
      {stage4_3[8]}
   );
   gpc1_1 gpc1997 (
      {stage3_3[27]},
      {stage4_3[9]}
   );
   gpc1_1 gpc1998 (
      {stage3_3[28]},
      {stage4_3[10]}
   );
   gpc1_1 gpc1999 (
      {stage3_4[20]},
      {stage4_4[7]}
   );
   gpc1_1 gpc2000 (
      {stage3_4[21]},
      {stage4_4[8]}
   );
   gpc1_1 gpc2001 (
      {stage3_4[22]},
      {stage4_4[9]}
   );
   gpc1_1 gpc2002 (
      {stage3_4[23]},
      {stage4_4[10]}
   );
   gpc1_1 gpc2003 (
      {stage3_4[24]},
      {stage4_4[11]}
   );
   gpc1_1 gpc2004 (
      {stage3_4[25]},
      {stage4_4[12]}
   );
   gpc1_1 gpc2005 (
      {stage3_4[26]},
      {stage4_4[13]}
   );
   gpc1_1 gpc2006 (
      {stage3_4[27]},
      {stage4_4[14]}
   );
   gpc1_1 gpc2007 (
      {stage3_4[28]},
      {stage4_4[15]}
   );
   gpc1_1 gpc2008 (
      {stage3_4[29]},
      {stage4_4[16]}
   );
   gpc1_1 gpc2009 (
      {stage3_4[30]},
      {stage4_4[17]}
   );
   gpc1_1 gpc2010 (
      {stage3_4[31]},
      {stage4_4[18]}
   );
   gpc1_1 gpc2011 (
      {stage3_4[32]},
      {stage4_4[19]}
   );
   gpc1_1 gpc2012 (
      {stage3_4[33]},
      {stage4_4[20]}
   );
   gpc1_1 gpc2013 (
      {stage3_4[34]},
      {stage4_4[21]}
   );
   gpc1_1 gpc2014 (
      {stage3_4[35]},
      {stage4_4[22]}
   );
   gpc1_1 gpc2015 (
      {stage3_4[36]},
      {stage4_4[23]}
   );
   gpc1_1 gpc2016 (
      {stage3_4[37]},
      {stage4_4[24]}
   );
   gpc1_1 gpc2017 (
      {stage3_4[38]},
      {stage4_4[25]}
   );
   gpc1_1 gpc2018 (
      {stage3_4[39]},
      {stage4_4[26]}
   );
   gpc1_1 gpc2019 (
      {stage3_5[47]},
      {stage4_5[14]}
   );
   gpc1_1 gpc2020 (
      {stage3_6[31]},
      {stage4_6[15]}
   );
   gpc1_1 gpc2021 (
      {stage3_6[32]},
      {stage4_6[16]}
   );
   gpc1_1 gpc2022 (
      {stage3_6[33]},
      {stage4_6[17]}
   );
   gpc1_1 gpc2023 (
      {stage3_6[34]},
      {stage4_6[18]}
   );
   gpc1_1 gpc2024 (
      {stage3_6[35]},
      {stage4_6[19]}
   );
   gpc1_1 gpc2025 (
      {stage3_6[36]},
      {stage4_6[20]}
   );
   gpc1_1 gpc2026 (
      {stage3_6[37]},
      {stage4_6[21]}
   );
   gpc1_1 gpc2027 (
      {stage3_7[42]},
      {stage4_7[13]}
   );
   gpc1_1 gpc2028 (
      {stage3_7[43]},
      {stage4_7[14]}
   );
   gpc1_1 gpc2029 (
      {stage3_7[44]},
      {stage4_7[15]}
   );
   gpc1_1 gpc2030 (
      {stage3_7[45]},
      {stage4_7[16]}
   );
   gpc1_1 gpc2031 (
      {stage3_8[28]},
      {stage4_8[13]}
   );
   gpc1_1 gpc2032 (
      {stage3_8[29]},
      {stage4_8[14]}
   );
   gpc1_1 gpc2033 (
      {stage3_8[30]},
      {stage4_8[15]}
   );
   gpc1_1 gpc2034 (
      {stage3_8[31]},
      {stage4_8[16]}
   );
   gpc1_1 gpc2035 (
      {stage3_8[32]},
      {stage4_8[17]}
   );
   gpc1_1 gpc2036 (
      {stage3_8[33]},
      {stage4_8[18]}
   );
   gpc1_1 gpc2037 (
      {stage3_8[34]},
      {stage4_8[19]}
   );
   gpc1_1 gpc2038 (
      {stage3_8[35]},
      {stage4_8[20]}
   );
   gpc1_1 gpc2039 (
      {stage3_8[36]},
      {stage4_8[21]}
   );
   gpc1_1 gpc2040 (
      {stage3_8[37]},
      {stage4_8[22]}
   );
   gpc1_1 gpc2041 (
      {stage3_8[38]},
      {stage4_8[23]}
   );
   gpc1_1 gpc2042 (
      {stage3_8[39]},
      {stage4_8[24]}
   );
   gpc1_1 gpc2043 (
      {stage3_8[40]},
      {stage4_8[25]}
   );
   gpc1_1 gpc2044 (
      {stage3_9[48]},
      {stage4_9[21]}
   );
   gpc1_1 gpc2045 (
      {stage3_9[49]},
      {stage4_9[22]}
   );
   gpc1_1 gpc2046 (
      {stage3_9[50]},
      {stage4_9[23]}
   );
   gpc1_1 gpc2047 (
      {stage3_9[51]},
      {stage4_9[24]}
   );
   gpc1_1 gpc2048 (
      {stage3_10[44]},
      {stage4_10[18]}
   );
   gpc1_1 gpc2049 (
      {stage3_10[45]},
      {stage4_10[19]}
   );
   gpc1_1 gpc2050 (
      {stage3_10[46]},
      {stage4_10[20]}
   );
   gpc1_1 gpc2051 (
      {stage3_10[47]},
      {stage4_10[21]}
   );
   gpc1_1 gpc2052 (
      {stage3_10[48]},
      {stage4_10[22]}
   );
   gpc1_1 gpc2053 (
      {stage3_10[49]},
      {stage4_10[23]}
   );
   gpc1_1 gpc2054 (
      {stage3_10[50]},
      {stage4_10[24]}
   );
   gpc1_1 gpc2055 (
      {stage3_10[51]},
      {stage4_10[25]}
   );
   gpc1_1 gpc2056 (
      {stage3_10[52]},
      {stage4_10[26]}
   );
   gpc1_1 gpc2057 (
      {stage3_10[53]},
      {stage4_10[27]}
   );
   gpc1_1 gpc2058 (
      {stage3_10[54]},
      {stage4_10[28]}
   );
   gpc1_1 gpc2059 (
      {stage3_10[55]},
      {stage4_10[29]}
   );
   gpc1_1 gpc2060 (
      {stage3_10[56]},
      {stage4_10[30]}
   );
   gpc1_1 gpc2061 (
      {stage3_10[57]},
      {stage4_10[31]}
   );
   gpc1_1 gpc2062 (
      {stage3_10[58]},
      {stage4_10[32]}
   );
   gpc1_1 gpc2063 (
      {stage3_10[59]},
      {stage4_10[33]}
   );
   gpc1_1 gpc2064 (
      {stage3_10[60]},
      {stage4_10[34]}
   );
   gpc1_1 gpc2065 (
      {stage3_10[61]},
      {stage4_10[35]}
   );
   gpc1_1 gpc2066 (
      {stage3_10[62]},
      {stage4_10[36]}
   );
   gpc1_1 gpc2067 (
      {stage3_10[63]},
      {stage4_10[37]}
   );
   gpc1_1 gpc2068 (
      {stage3_11[54]},
      {stage4_11[15]}
   );
   gpc1_1 gpc2069 (
      {stage3_11[55]},
      {stage4_11[16]}
   );
   gpc1_1 gpc2070 (
      {stage3_11[56]},
      {stage4_11[17]}
   );
   gpc1_1 gpc2071 (
      {stage3_11[57]},
      {stage4_11[18]}
   );
   gpc1_1 gpc2072 (
      {stage3_11[58]},
      {stage4_11[19]}
   );
   gpc1_1 gpc2073 (
      {stage3_11[59]},
      {stage4_11[20]}
   );
   gpc1_1 gpc2074 (
      {stage3_11[60]},
      {stage4_11[21]}
   );
   gpc1_1 gpc2075 (
      {stage3_12[48]},
      {stage4_12[19]}
   );
   gpc1_1 gpc2076 (
      {stage3_12[49]},
      {stage4_12[20]}
   );
   gpc1_1 gpc2077 (
      {stage3_12[50]},
      {stage4_12[21]}
   );
   gpc1_1 gpc2078 (
      {stage3_12[51]},
      {stage4_12[22]}
   );
   gpc1_1 gpc2079 (
      {stage3_12[52]},
      {stage4_12[23]}
   );
   gpc1_1 gpc2080 (
      {stage3_15[53]},
      {stage4_15[18]}
   );
   gpc1_1 gpc2081 (
      {stage3_15[54]},
      {stage4_15[19]}
   );
   gpc1_1 gpc2082 (
      {stage3_15[55]},
      {stage4_15[20]}
   );
   gpc1_1 gpc2083 (
      {stage3_15[56]},
      {stage4_15[21]}
   );
   gpc1_1 gpc2084 (
      {stage3_16[41]},
      {stage4_16[22]}
   );
   gpc1_1 gpc2085 (
      {stage3_16[42]},
      {stage4_16[23]}
   );
   gpc1_1 gpc2086 (
      {stage3_16[43]},
      {stage4_16[24]}
   );
   gpc1_1 gpc2087 (
      {stage3_16[44]},
      {stage4_16[25]}
   );
   gpc1_1 gpc2088 (
      {stage3_16[45]},
      {stage4_16[26]}
   );
   gpc1_1 gpc2089 (
      {stage3_16[46]},
      {stage4_16[27]}
   );
   gpc1_1 gpc2090 (
      {stage3_16[47]},
      {stage4_16[28]}
   );
   gpc1_1 gpc2091 (
      {stage3_16[48]},
      {stage4_16[29]}
   );
   gpc1_1 gpc2092 (
      {stage3_16[49]},
      {stage4_16[30]}
   );
   gpc1_1 gpc2093 (
      {stage3_17[30]},
      {stage4_17[20]}
   );
   gpc1_1 gpc2094 (
      {stage3_17[31]},
      {stage4_17[21]}
   );
   gpc1_1 gpc2095 (
      {stage3_18[24]},
      {stage4_18[11]}
   );
   gpc1_1 gpc2096 (
      {stage3_18[25]},
      {stage4_18[12]}
   );
   gpc1_1 gpc2097 (
      {stage3_19[12]},
      {stage4_19[9]}
   );
   gpc1_1 gpc2098 (
      {stage3_19[13]},
      {stage4_19[10]}
   );
   gpc1_1 gpc2099 (
      {stage3_20[0]},
      {stage4_20[6]}
   );
   gpc1_1 gpc2100 (
      {stage3_20[1]},
      {stage4_20[7]}
   );
   gpc1_1 gpc2101 (
      {stage3_20[2]},
      {stage4_20[8]}
   );
   gpc1_1 gpc2102 (
      {stage3_20[3]},
      {stage4_20[9]}
   );
   gpc1_1 gpc2103 (
      {stage3_20[4]},
      {stage4_20[10]}
   );
   gpc1_1 gpc2104 (
      {stage3_20[5]},
      {stage4_20[11]}
   );
   gpc1_1 gpc2105 (
      {stage3_21[0]},
      {stage4_21[2]}
   );
   gpc1_1 gpc2106 (
      {stage3_21[1]},
      {stage4_21[3]}
   );
   gpc615_5 gpc2107 (
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4]},
      {stage4_3[0]},
      {stage4_4[0], stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5]},
      {stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[0],stage5_2[0]}
   );
   gpc606_5 gpc2108 (
      {stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5], stage4_3[6]},
      {stage4_5[0], stage4_5[1], stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5]},
      {stage5_7[0],stage5_6[1],stage5_5[1],stage5_4[1],stage5_3[1]}
   );
   gpc1406_5 gpc2109 (
      {stage4_4[6], stage4_4[7], stage4_4[8], stage4_4[9], stage4_4[10], stage4_4[11]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3]},
      {stage4_7[0]},
      {stage5_8[0],stage5_7[1],stage5_6[2],stage5_5[2],stage5_4[2]}
   );
   gpc606_5 gpc2110 (
      {stage4_4[12], stage4_4[13], stage4_4[14], stage4_4[15], stage4_4[16], stage4_4[17]},
      {stage4_6[4], stage4_6[5], stage4_6[6], stage4_6[7], stage4_6[8], stage4_6[9]},
      {stage5_8[1],stage5_7[2],stage5_6[3],stage5_5[3],stage5_4[3]}
   );
   gpc606_5 gpc2111 (
      {stage4_5[6], stage4_5[7], stage4_5[8], stage4_5[9], stage4_5[10], stage4_5[11]},
      {stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5], stage4_7[6]},
      {stage5_9[0],stage5_8[2],stage5_7[3],stage5_6[4],stage5_5[4]}
   );
   gpc615_5 gpc2112 (
      {stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10], stage4_7[11]},
      {stage4_8[0]},
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5]},
      {stage5_11[0],stage5_10[0],stage5_9[1],stage5_8[3],stage5_7[4]}
   );
   gpc615_5 gpc2113 (
      {stage4_7[12], stage4_7[13], stage4_7[14], stage4_7[15], stage4_7[16]},
      {stage4_8[1]},
      {stage4_9[6], stage4_9[7], stage4_9[8], stage4_9[9], stage4_9[10], stage4_9[11]},
      {stage5_11[1],stage5_10[1],stage5_9[2],stage5_8[4],stage5_7[5]}
   );
   gpc1163_5 gpc2114 (
      {stage4_8[2], stage4_8[3], stage4_8[4]},
      {stage4_9[12], stage4_9[13], stage4_9[14], stage4_9[15], stage4_9[16], stage4_9[17]},
      {stage4_10[0]},
      {stage4_11[0]},
      {stage5_12[0],stage5_11[2],stage5_10[2],stage5_9[3],stage5_8[5]}
   );
   gpc1163_5 gpc2115 (
      {stage4_8[5], stage4_8[6], stage4_8[7]},
      {stage4_9[18], stage4_9[19], stage4_9[20], stage4_9[21], stage4_9[22], stage4_9[23]},
      {stage4_10[1]},
      {stage4_11[1]},
      {stage5_12[1],stage5_11[3],stage5_10[3],stage5_9[4],stage5_8[6]}
   );
   gpc606_5 gpc2116 (
      {stage4_8[8], stage4_8[9], stage4_8[10], stage4_8[11], stage4_8[12], stage4_8[13]},
      {stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7]},
      {stage5_12[2],stage5_11[4],stage5_10[4],stage5_9[5],stage5_8[7]}
   );
   gpc606_5 gpc2117 (
      {stage4_8[14], stage4_8[15], stage4_8[16], stage4_8[17], stage4_8[18], stage4_8[19]},
      {stage4_10[8], stage4_10[9], stage4_10[10], stage4_10[11], stage4_10[12], stage4_10[13]},
      {stage5_12[3],stage5_11[5],stage5_10[5],stage5_9[6],stage5_8[8]}
   );
   gpc606_5 gpc2118 (
      {stage4_8[20], stage4_8[21], stage4_8[22], stage4_8[23], stage4_8[24], stage4_8[25]},
      {stage4_10[14], stage4_10[15], stage4_10[16], stage4_10[17], stage4_10[18], stage4_10[19]},
      {stage5_12[4],stage5_11[6],stage5_10[6],stage5_9[7],stage5_8[9]}
   );
   gpc606_5 gpc2119 (
      {stage4_10[20], stage4_10[21], stage4_10[22], stage4_10[23], stage4_10[24], stage4_10[25]},
      {stage4_12[0], stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5]},
      {stage5_14[0],stage5_13[0],stage5_12[5],stage5_11[7],stage5_10[7]}
   );
   gpc606_5 gpc2120 (
      {stage4_10[26], stage4_10[27], stage4_10[28], stage4_10[29], stage4_10[30], stage4_10[31]},
      {stage4_12[6], stage4_12[7], stage4_12[8], stage4_12[9], stage4_12[10], stage4_12[11]},
      {stage5_14[1],stage5_13[1],stage5_12[6],stage5_11[8],stage5_10[8]}
   );
   gpc615_5 gpc2121 (
      {stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5], stage4_11[6]},
      {stage4_12[12]},
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5]},
      {stage5_15[0],stage5_14[2],stage5_13[2],stage5_12[7],stage5_11[9]}
   );
   gpc615_5 gpc2122 (
      {stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11]},
      {stage4_12[13]},
      {stage4_13[6], stage4_13[7], stage4_13[8], stage4_13[9], stage4_13[10], stage4_13[11]},
      {stage5_15[1],stage5_14[3],stage5_13[3],stage5_12[8],stage5_11[10]}
   );
   gpc615_5 gpc2123 (
      {stage4_11[12], stage4_11[13], stage4_11[14], stage4_11[15], stage4_11[16]},
      {stage4_12[14]},
      {stage4_13[12], stage4_13[13], stage4_13[14], stage4_13[15], stage4_13[16], stage4_13[17]},
      {stage5_15[2],stage5_14[4],stage5_13[4],stage5_12[9],stage5_11[11]}
   );
   gpc615_5 gpc2124 (
      {stage4_11[17], stage4_11[18], stage4_11[19], stage4_11[20], stage4_11[21]},
      {stage4_12[15]},
      {stage4_13[18], stage4_13[19], stage4_13[20], stage4_13[21], stage4_13[22], stage4_13[23]},
      {stage5_15[3],stage5_14[5],stage5_13[5],stage5_12[10],stage5_11[12]}
   );
   gpc606_5 gpc2125 (
      {stage4_12[16], stage4_12[17], stage4_12[18], stage4_12[19], stage4_12[20], stage4_12[21]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[4],stage5_14[6],stage5_13[6],stage5_12[11]}
   );
   gpc615_5 gpc2126 (
      {stage4_14[6], stage4_14[7], stage4_14[8], stage4_14[9], stage4_14[10]},
      {stage4_15[0]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[5],stage5_14[7]}
   );
   gpc615_5 gpc2127 (
      {stage4_14[11], stage4_14[12], stage4_14[13], stage4_14[14], stage4_14[15]},
      {stage4_15[1]},
      {stage4_16[6], stage4_16[7], stage4_16[8], stage4_16[9], stage4_16[10], stage4_16[11]},
      {stage5_18[1],stage5_17[1],stage5_16[2],stage5_15[6],stage5_14[8]}
   );
   gpc615_5 gpc2128 (
      {stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5], stage4_15[6]},
      {stage4_16[12]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[2],stage5_17[2],stage5_16[3],stage5_15[7]}
   );
   gpc615_5 gpc2129 (
      {stage4_15[7], stage4_15[8], stage4_15[9], stage4_15[10], stage4_15[11]},
      {stage4_16[13]},
      {stage4_17[6], stage4_17[7], stage4_17[8], stage4_17[9], stage4_17[10], stage4_17[11]},
      {stage5_19[1],stage5_18[3],stage5_17[3],stage5_16[4],stage5_15[8]}
   );
   gpc615_5 gpc2130 (
      {stage4_15[12], stage4_15[13], stage4_15[14], stage4_15[15], stage4_15[16]},
      {stage4_16[14]},
      {stage4_17[12], stage4_17[13], stage4_17[14], stage4_17[15], stage4_17[16], stage4_17[17]},
      {stage5_19[2],stage5_18[4],stage5_17[4],stage5_16[5],stage5_15[9]}
   );
   gpc606_5 gpc2131 (
      {stage4_16[15], stage4_16[16], stage4_16[17], stage4_16[18], stage4_16[19], stage4_16[20]},
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage5_20[0],stage5_19[3],stage5_18[5],stage5_17[5],stage5_16[6]}
   );
   gpc606_5 gpc2132 (
      {stage4_17[18], stage4_17[19], stage4_17[20], stage4_17[21], 1'b0, 1'b0},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[1],stage5_19[4],stage5_18[6],stage5_17[6]}
   );
   gpc606_5 gpc2133 (
      {stage4_18[6], stage4_18[7], stage4_18[8], stage4_18[9], stage4_18[10], stage4_18[11]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[1],stage5_20[2],stage5_19[5],stage5_18[7]}
   );
   gpc1343_5 gpc2134 (
      {stage4_19[6], stage4_19[7], stage4_19[8]},
      {stage4_20[6], stage4_20[7], stage4_20[8], stage4_20[9]},
      {stage4_21[0], stage4_21[1], stage4_21[2]},
      {1'b0},
      {stage5_23[0],stage5_22[1],stage5_21[2],stage5_20[3],stage5_19[6]}
   );
   gpc1_1 gpc2135 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc2136 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc2137 (
      {stage4_0[2]},
      {stage5_0[2]}
   );
   gpc1_1 gpc2138 (
      {stage4_0[3]},
      {stage5_0[3]}
   );
   gpc1_1 gpc2139 (
      {stage4_0[4]},
      {stage5_0[4]}
   );
   gpc1_1 gpc2140 (
      {stage4_0[5]},
      {stage5_0[5]}
   );
   gpc1_1 gpc2141 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc2142 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc2143 (
      {stage4_2[5]},
      {stage5_2[1]}
   );
   gpc1_1 gpc2144 (
      {stage4_2[6]},
      {stage5_2[2]}
   );
   gpc1_1 gpc2145 (
      {stage4_2[7]},
      {stage5_2[3]}
   );
   gpc1_1 gpc2146 (
      {stage4_2[8]},
      {stage5_2[4]}
   );
   gpc1_1 gpc2147 (
      {stage4_2[9]},
      {stage5_2[5]}
   );
   gpc1_1 gpc2148 (
      {stage4_2[10]},
      {stage5_2[6]}
   );
   gpc1_1 gpc2149 (
      {stage4_3[7]},
      {stage5_3[2]}
   );
   gpc1_1 gpc2150 (
      {stage4_3[8]},
      {stage5_3[3]}
   );
   gpc1_1 gpc2151 (
      {stage4_3[9]},
      {stage5_3[4]}
   );
   gpc1_1 gpc2152 (
      {stage4_3[10]},
      {stage5_3[5]}
   );
   gpc1_1 gpc2153 (
      {stage4_4[18]},
      {stage5_4[4]}
   );
   gpc1_1 gpc2154 (
      {stage4_4[19]},
      {stage5_4[5]}
   );
   gpc1_1 gpc2155 (
      {stage4_4[20]},
      {stage5_4[6]}
   );
   gpc1_1 gpc2156 (
      {stage4_4[21]},
      {stage5_4[7]}
   );
   gpc1_1 gpc2157 (
      {stage4_4[22]},
      {stage5_4[8]}
   );
   gpc1_1 gpc2158 (
      {stage4_4[23]},
      {stage5_4[9]}
   );
   gpc1_1 gpc2159 (
      {stage4_4[24]},
      {stage5_4[10]}
   );
   gpc1_1 gpc2160 (
      {stage4_4[25]},
      {stage5_4[11]}
   );
   gpc1_1 gpc2161 (
      {stage4_4[26]},
      {stage5_4[12]}
   );
   gpc1_1 gpc2162 (
      {stage4_5[12]},
      {stage5_5[5]}
   );
   gpc1_1 gpc2163 (
      {stage4_5[13]},
      {stage5_5[6]}
   );
   gpc1_1 gpc2164 (
      {stage4_5[14]},
      {stage5_5[7]}
   );
   gpc1_1 gpc2165 (
      {stage4_6[10]},
      {stage5_6[5]}
   );
   gpc1_1 gpc2166 (
      {stage4_6[11]},
      {stage5_6[6]}
   );
   gpc1_1 gpc2167 (
      {stage4_6[12]},
      {stage5_6[7]}
   );
   gpc1_1 gpc2168 (
      {stage4_6[13]},
      {stage5_6[8]}
   );
   gpc1_1 gpc2169 (
      {stage4_6[14]},
      {stage5_6[9]}
   );
   gpc1_1 gpc2170 (
      {stage4_6[15]},
      {stage5_6[10]}
   );
   gpc1_1 gpc2171 (
      {stage4_6[16]},
      {stage5_6[11]}
   );
   gpc1_1 gpc2172 (
      {stage4_6[17]},
      {stage5_6[12]}
   );
   gpc1_1 gpc2173 (
      {stage4_6[18]},
      {stage5_6[13]}
   );
   gpc1_1 gpc2174 (
      {stage4_6[19]},
      {stage5_6[14]}
   );
   gpc1_1 gpc2175 (
      {stage4_6[20]},
      {stage5_6[15]}
   );
   gpc1_1 gpc2176 (
      {stage4_6[21]},
      {stage5_6[16]}
   );
   gpc1_1 gpc2177 (
      {stage4_9[24]},
      {stage5_9[8]}
   );
   gpc1_1 gpc2178 (
      {stage4_10[32]},
      {stage5_10[9]}
   );
   gpc1_1 gpc2179 (
      {stage4_10[33]},
      {stage5_10[10]}
   );
   gpc1_1 gpc2180 (
      {stage4_10[34]},
      {stage5_10[11]}
   );
   gpc1_1 gpc2181 (
      {stage4_10[35]},
      {stage5_10[12]}
   );
   gpc1_1 gpc2182 (
      {stage4_10[36]},
      {stage5_10[13]}
   );
   gpc1_1 gpc2183 (
      {stage4_10[37]},
      {stage5_10[14]}
   );
   gpc1_1 gpc2184 (
      {stage4_12[22]},
      {stage5_12[12]}
   );
   gpc1_1 gpc2185 (
      {stage4_12[23]},
      {stage5_12[13]}
   );
   gpc1_1 gpc2186 (
      {stage4_13[24]},
      {stage5_13[7]}
   );
   gpc1_1 gpc2187 (
      {stage4_13[25]},
      {stage5_13[8]}
   );
   gpc1_1 gpc2188 (
      {stage4_14[16]},
      {stage5_14[9]}
   );
   gpc1_1 gpc2189 (
      {stage4_14[17]},
      {stage5_14[10]}
   );
   gpc1_1 gpc2190 (
      {stage4_14[18]},
      {stage5_14[11]}
   );
   gpc1_1 gpc2191 (
      {stage4_15[17]},
      {stage5_15[10]}
   );
   gpc1_1 gpc2192 (
      {stage4_15[18]},
      {stage5_15[11]}
   );
   gpc1_1 gpc2193 (
      {stage4_15[19]},
      {stage5_15[12]}
   );
   gpc1_1 gpc2194 (
      {stage4_15[20]},
      {stage5_15[13]}
   );
   gpc1_1 gpc2195 (
      {stage4_15[21]},
      {stage5_15[14]}
   );
   gpc1_1 gpc2196 (
      {stage4_16[21]},
      {stage5_16[7]}
   );
   gpc1_1 gpc2197 (
      {stage4_16[22]},
      {stage5_16[8]}
   );
   gpc1_1 gpc2198 (
      {stage4_16[23]},
      {stage5_16[9]}
   );
   gpc1_1 gpc2199 (
      {stage4_16[24]},
      {stage5_16[10]}
   );
   gpc1_1 gpc2200 (
      {stage4_16[25]},
      {stage5_16[11]}
   );
   gpc1_1 gpc2201 (
      {stage4_16[26]},
      {stage5_16[12]}
   );
   gpc1_1 gpc2202 (
      {stage4_16[27]},
      {stage5_16[13]}
   );
   gpc1_1 gpc2203 (
      {stage4_16[28]},
      {stage5_16[14]}
   );
   gpc1_1 gpc2204 (
      {stage4_16[29]},
      {stage5_16[15]}
   );
   gpc1_1 gpc2205 (
      {stage4_16[30]},
      {stage5_16[16]}
   );
   gpc1_1 gpc2206 (
      {stage4_18[12]},
      {stage5_18[8]}
   );
   gpc1_1 gpc2207 (
      {stage4_19[9]},
      {stage5_19[7]}
   );
   gpc1_1 gpc2208 (
      {stage4_19[10]},
      {stage5_19[8]}
   );
   gpc1_1 gpc2209 (
      {stage4_20[10]},
      {stage5_20[4]}
   );
   gpc1_1 gpc2210 (
      {stage4_20[11]},
      {stage5_20[5]}
   );
   gpc1_1 gpc2211 (
      {stage4_21[3]},
      {stage5_21[3]}
   );
   gpc1163_5 gpc2212 (
      {stage5_2[0], stage5_2[1], stage5_2[2]},
      {stage5_3[0], stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4], stage5_3[5]},
      {stage5_4[0]},
      {stage5_5[0]},
      {stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0]}
   );
   gpc207_4 gpc2213 (
      {stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5], stage5_4[6], stage5_4[7]},
      {stage5_6[0], stage5_6[1]},
      {stage6_7[0],stage6_6[1],stage6_5[1],stage6_4[1]}
   );
   gpc7_3 gpc2214 (
      {stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4], stage5_5[5], stage5_5[6], stage5_5[7]},
      {stage6_7[1],stage6_6[2],stage6_5[2]}
   );
   gpc1325_5 gpc2215 (
      {stage5_6[2], stage5_6[3], stage5_6[4], stage5_6[5], stage5_6[6]},
      {stage5_7[0], stage5_7[1]},
      {stage5_8[0], stage5_8[1], stage5_8[2]},
      {stage5_9[0]},
      {stage6_10[0],stage6_9[0],stage6_8[0],stage6_7[2],stage6_6[3]}
   );
   gpc1325_5 gpc2216 (
      {stage5_6[7], stage5_6[8], stage5_6[9], stage5_6[10], stage5_6[11]},
      {stage5_7[2], stage5_7[3]},
      {stage5_8[3], stage5_8[4], stage5_8[5]},
      {stage5_9[1]},
      {stage6_10[1],stage6_9[1],stage6_8[1],stage6_7[3],stage6_6[4]}
   );
   gpc1325_5 gpc2217 (
      {stage5_6[12], stage5_6[13], stage5_6[14], stage5_6[15], stage5_6[16]},
      {stage5_7[4], stage5_7[5]},
      {stage5_8[6], stage5_8[7], stage5_8[8]},
      {stage5_9[2]},
      {stage6_10[2],stage6_9[2],stage6_8[2],stage6_7[4],stage6_6[5]}
   );
   gpc1163_5 gpc2218 (
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0], stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5]},
      {stage5_12[0]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[0],stage6_12[0],stage6_11[0],stage6_10[3]}
   );
   gpc1163_5 gpc2219 (
      {stage5_10[3], stage5_10[4], stage5_10[5]},
      {stage5_11[6], stage5_11[7], stage5_11[8], stage5_11[9], stage5_11[10], stage5_11[11]},
      {stage5_12[1]},
      {stage5_13[1]},
      {stage6_14[1],stage6_13[1],stage6_12[1],stage6_11[1],stage6_10[4]}
   );
   gpc615_5 gpc2220 (
      {stage5_10[6], stage5_10[7], stage5_10[8], stage5_10[9], stage5_10[10]},
      {stage5_11[12]},
      {stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5], stage5_12[6], stage5_12[7]},
      {stage6_14[2],stage6_13[2],stage6_12[2],stage6_11[2],stage6_10[5]}
   );
   gpc2116_5 gpc2221 (
      {stage5_12[8], stage5_12[9], stage5_12[10], stage5_12[11], stage5_12[12], stage5_12[13]},
      {stage5_13[2]},
      {stage5_14[0]},
      {stage5_15[0], stage5_15[1]},
      {stage6_16[0],stage6_15[0],stage6_14[3],stage6_13[3],stage6_12[3]}
   );
   gpc623_5 gpc2222 (
      {stage5_13[3], stage5_13[4], stage5_13[5]},
      {stage5_14[1], stage5_14[2]},
      {stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5], stage5_15[6], stage5_15[7]},
      {stage6_17[0],stage6_16[1],stage6_15[1],stage6_14[4],stage6_13[4]}
   );
   gpc1423_5 gpc2223 (
      {stage5_14[3], stage5_14[4], stage5_14[5]},
      {stage5_15[8], stage5_15[9]},
      {stage5_16[0], stage5_16[1], stage5_16[2], stage5_16[3]},
      {stage5_17[0]},
      {stage6_18[0],stage6_17[1],stage6_16[2],stage6_15[2],stage6_14[5]}
   );
   gpc615_5 gpc2224 (
      {stage5_14[6], stage5_14[7], stage5_14[8], stage5_14[9], stage5_14[10]},
      {stage5_15[10]},
      {stage5_16[4], stage5_16[5], stage5_16[6], stage5_16[7], stage5_16[8], stage5_16[9]},
      {stage6_18[1],stage6_17[2],stage6_16[3],stage6_15[3],stage6_14[6]}
   );
   gpc606_5 gpc2225 (
      {stage5_16[10], stage5_16[11], stage5_16[12], stage5_16[13], stage5_16[14], stage5_16[15]},
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5]},
      {stage6_20[0],stage6_19[0],stage6_18[2],stage6_17[3],stage6_16[4]}
   );
   gpc606_5 gpc2226 (
      {stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5], stage5_17[6]},
      {stage5_19[0], stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage6_21[0],stage6_20[1],stage6_19[1],stage6_18[3],stage6_17[4]}
   );
   gpc1_1 gpc2227 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc2228 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc2229 (
      {stage5_0[2]},
      {stage6_0[2]}
   );
   gpc1_1 gpc2230 (
      {stage5_0[3]},
      {stage6_0[3]}
   );
   gpc1_1 gpc2231 (
      {stage5_0[4]},
      {stage6_0[4]}
   );
   gpc1_1 gpc2232 (
      {stage5_0[5]},
      {stage6_0[5]}
   );
   gpc1_1 gpc2233 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc2234 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc2235 (
      {stage5_2[3]},
      {stage6_2[1]}
   );
   gpc1_1 gpc2236 (
      {stage5_2[4]},
      {stage6_2[2]}
   );
   gpc1_1 gpc2237 (
      {stage5_2[5]},
      {stage6_2[3]}
   );
   gpc1_1 gpc2238 (
      {stage5_2[6]},
      {stage6_2[4]}
   );
   gpc1_1 gpc2239 (
      {stage5_4[8]},
      {stage6_4[2]}
   );
   gpc1_1 gpc2240 (
      {stage5_4[9]},
      {stage6_4[3]}
   );
   gpc1_1 gpc2241 (
      {stage5_4[10]},
      {stage6_4[4]}
   );
   gpc1_1 gpc2242 (
      {stage5_4[11]},
      {stage6_4[5]}
   );
   gpc1_1 gpc2243 (
      {stage5_4[12]},
      {stage6_4[6]}
   );
   gpc1_1 gpc2244 (
      {stage5_8[9]},
      {stage6_8[3]}
   );
   gpc1_1 gpc2245 (
      {stage5_9[3]},
      {stage6_9[3]}
   );
   gpc1_1 gpc2246 (
      {stage5_9[4]},
      {stage6_9[4]}
   );
   gpc1_1 gpc2247 (
      {stage5_9[5]},
      {stage6_9[5]}
   );
   gpc1_1 gpc2248 (
      {stage5_9[6]},
      {stage6_9[6]}
   );
   gpc1_1 gpc2249 (
      {stage5_9[7]},
      {stage6_9[7]}
   );
   gpc1_1 gpc2250 (
      {stage5_9[8]},
      {stage6_9[8]}
   );
   gpc1_1 gpc2251 (
      {stage5_10[11]},
      {stage6_10[6]}
   );
   gpc1_1 gpc2252 (
      {stage5_10[12]},
      {stage6_10[7]}
   );
   gpc1_1 gpc2253 (
      {stage5_10[13]},
      {stage6_10[8]}
   );
   gpc1_1 gpc2254 (
      {stage5_10[14]},
      {stage6_10[9]}
   );
   gpc1_1 gpc2255 (
      {stage5_13[6]},
      {stage6_13[5]}
   );
   gpc1_1 gpc2256 (
      {stage5_13[7]},
      {stage6_13[6]}
   );
   gpc1_1 gpc2257 (
      {stage5_13[8]},
      {stage6_13[7]}
   );
   gpc1_1 gpc2258 (
      {stage5_14[11]},
      {stage6_14[7]}
   );
   gpc1_1 gpc2259 (
      {stage5_15[11]},
      {stage6_15[4]}
   );
   gpc1_1 gpc2260 (
      {stage5_15[12]},
      {stage6_15[5]}
   );
   gpc1_1 gpc2261 (
      {stage5_15[13]},
      {stage6_15[6]}
   );
   gpc1_1 gpc2262 (
      {stage5_15[14]},
      {stage6_15[7]}
   );
   gpc1_1 gpc2263 (
      {stage5_16[16]},
      {stage6_16[5]}
   );
   gpc1_1 gpc2264 (
      {stage5_18[6]},
      {stage6_18[4]}
   );
   gpc1_1 gpc2265 (
      {stage5_18[7]},
      {stage6_18[5]}
   );
   gpc1_1 gpc2266 (
      {stage5_18[8]},
      {stage6_18[6]}
   );
   gpc1_1 gpc2267 (
      {stage5_19[6]},
      {stage6_19[2]}
   );
   gpc1_1 gpc2268 (
      {stage5_19[7]},
      {stage6_19[3]}
   );
   gpc1_1 gpc2269 (
      {stage5_19[8]},
      {stage6_19[4]}
   );
   gpc1_1 gpc2270 (
      {stage5_20[0]},
      {stage6_20[2]}
   );
   gpc1_1 gpc2271 (
      {stage5_20[1]},
      {stage6_20[3]}
   );
   gpc1_1 gpc2272 (
      {stage5_20[2]},
      {stage6_20[4]}
   );
   gpc1_1 gpc2273 (
      {stage5_20[3]},
      {stage6_20[5]}
   );
   gpc1_1 gpc2274 (
      {stage5_20[4]},
      {stage6_20[6]}
   );
   gpc1_1 gpc2275 (
      {stage5_20[5]},
      {stage6_20[7]}
   );
   gpc1_1 gpc2276 (
      {stage5_21[0]},
      {stage6_21[1]}
   );
   gpc1_1 gpc2277 (
      {stage5_21[1]},
      {stage6_21[2]}
   );
   gpc1_1 gpc2278 (
      {stage5_21[2]},
      {stage6_21[3]}
   );
   gpc1_1 gpc2279 (
      {stage5_21[3]},
      {stage6_21[4]}
   );
   gpc1_1 gpc2280 (
      {stage5_22[0]},
      {stage6_22[0]}
   );
   gpc1_1 gpc2281 (
      {stage5_22[1]},
      {stage6_22[1]}
   );
   gpc1_1 gpc2282 (
      {stage5_23[0]},
      {stage6_23[0]}
   );
   gpc1406_5 gpc2283 (
      {stage6_6[0], stage6_6[1], stage6_6[2], stage6_6[3], stage6_6[4], stage6_6[5]},
      {stage6_8[0], stage6_8[1], stage6_8[2], stage6_8[3]},
      {stage6_9[0]},
      {stage7_10[0],stage7_9[0],stage7_8[0],stage7_7[0],stage7_6[0]}
   );
   gpc117_4 gpc2284 (
      {stage6_9[1], stage6_9[2], stage6_9[3], stage6_9[4], stage6_9[5], stage6_9[6], stage6_9[7]},
      {stage6_10[0]},
      {stage6_11[0]},
      {stage7_12[0],stage7_11[0],stage7_10[1],stage7_9[1]}
   );
   gpc1415_5 gpc2285 (
      {stage6_10[1], stage6_10[2], stage6_10[3], stage6_10[4], stage6_10[5]},
      {stage6_11[1]},
      {stage6_12[0], stage6_12[1], stage6_12[2], stage6_12[3]},
      {stage6_13[0]},
      {stage7_14[0],stage7_13[0],stage7_12[1],stage7_11[1],stage7_10[2]}
   );
   gpc606_5 gpc2286 (
      {stage6_13[1], stage6_13[2], stage6_13[3], stage6_13[4], stage6_13[5], stage6_13[6]},
      {stage6_15[0], stage6_15[1], stage6_15[2], stage6_15[3], stage6_15[4], stage6_15[5]},
      {stage7_17[0],stage7_16[0],stage7_15[0],stage7_14[1],stage7_13[1]}
   );
   gpc606_5 gpc2287 (
      {stage6_14[0], stage6_14[1], stage6_14[2], stage6_14[3], stage6_14[4], stage6_14[5]},
      {stage6_16[0], stage6_16[1], stage6_16[2], stage6_16[3], stage6_16[4], stage6_16[5]},
      {stage7_18[0],stage7_17[1],stage7_16[1],stage7_15[1],stage7_14[2]}
   );
   gpc606_5 gpc2288 (
      {stage6_18[0], stage6_18[1], stage6_18[2], stage6_18[3], stage6_18[4], stage6_18[5]},
      {stage6_20[0], stage6_20[1], stage6_20[2], stage6_20[3], stage6_20[4], stage6_20[5]},
      {stage7_22[0],stage7_21[0],stage7_20[0],stage7_19[0],stage7_18[1]}
   );
   gpc1406_5 gpc2289 (
      {stage6_19[0], stage6_19[1], stage6_19[2], stage6_19[3], stage6_19[4], 1'b0},
      {stage6_21[0], stage6_21[1], stage6_21[2], stage6_21[3]},
      {stage6_22[0]},
      {stage7_23[0],stage7_22[1],stage7_21[1],stage7_20[1],stage7_19[1]}
   );
   gpc1_1 gpc2290 (
      {stage6_0[0]},
      {stage7_0[0]}
   );
   gpc1_1 gpc2291 (
      {stage6_0[1]},
      {stage7_0[1]}
   );
   gpc1_1 gpc2292 (
      {stage6_0[2]},
      {stage7_0[2]}
   );
   gpc1_1 gpc2293 (
      {stage6_0[3]},
      {stage7_0[3]}
   );
   gpc1_1 gpc2294 (
      {stage6_0[4]},
      {stage7_0[4]}
   );
   gpc1_1 gpc2295 (
      {stage6_0[5]},
      {stage7_0[5]}
   );
   gpc1_1 gpc2296 (
      {stage6_1[0]},
      {stage7_1[0]}
   );
   gpc1_1 gpc2297 (
      {stage6_1[1]},
      {stage7_1[1]}
   );
   gpc1_1 gpc2298 (
      {stage6_2[0]},
      {stage7_2[0]}
   );
   gpc1_1 gpc2299 (
      {stage6_2[1]},
      {stage7_2[1]}
   );
   gpc1_1 gpc2300 (
      {stage6_2[2]},
      {stage7_2[2]}
   );
   gpc1_1 gpc2301 (
      {stage6_2[3]},
      {stage7_2[3]}
   );
   gpc1_1 gpc2302 (
      {stage6_2[4]},
      {stage7_2[4]}
   );
   gpc1_1 gpc2303 (
      {stage6_3[0]},
      {stage7_3[0]}
   );
   gpc1_1 gpc2304 (
      {stage6_4[0]},
      {stage7_4[0]}
   );
   gpc1_1 gpc2305 (
      {stage6_4[1]},
      {stage7_4[1]}
   );
   gpc1_1 gpc2306 (
      {stage6_4[2]},
      {stage7_4[2]}
   );
   gpc1_1 gpc2307 (
      {stage6_4[3]},
      {stage7_4[3]}
   );
   gpc1_1 gpc2308 (
      {stage6_4[4]},
      {stage7_4[4]}
   );
   gpc1_1 gpc2309 (
      {stage6_4[5]},
      {stage7_4[5]}
   );
   gpc1_1 gpc2310 (
      {stage6_4[6]},
      {stage7_4[6]}
   );
   gpc1_1 gpc2311 (
      {stage6_5[0]},
      {stage7_5[0]}
   );
   gpc1_1 gpc2312 (
      {stage6_5[1]},
      {stage7_5[1]}
   );
   gpc1_1 gpc2313 (
      {stage6_5[2]},
      {stage7_5[2]}
   );
   gpc1_1 gpc2314 (
      {stage6_7[0]},
      {stage7_7[1]}
   );
   gpc1_1 gpc2315 (
      {stage6_7[1]},
      {stage7_7[2]}
   );
   gpc1_1 gpc2316 (
      {stage6_7[2]},
      {stage7_7[3]}
   );
   gpc1_1 gpc2317 (
      {stage6_7[3]},
      {stage7_7[4]}
   );
   gpc1_1 gpc2318 (
      {stage6_7[4]},
      {stage7_7[5]}
   );
   gpc1_1 gpc2319 (
      {stage6_9[8]},
      {stage7_9[2]}
   );
   gpc1_1 gpc2320 (
      {stage6_10[6]},
      {stage7_10[3]}
   );
   gpc1_1 gpc2321 (
      {stage6_10[7]},
      {stage7_10[4]}
   );
   gpc1_1 gpc2322 (
      {stage6_10[8]},
      {stage7_10[5]}
   );
   gpc1_1 gpc2323 (
      {stage6_10[9]},
      {stage7_10[6]}
   );
   gpc1_1 gpc2324 (
      {stage6_11[2]},
      {stage7_11[2]}
   );
   gpc1_1 gpc2325 (
      {stage6_13[7]},
      {stage7_13[2]}
   );
   gpc1_1 gpc2326 (
      {stage6_14[6]},
      {stage7_14[3]}
   );
   gpc1_1 gpc2327 (
      {stage6_14[7]},
      {stage7_14[4]}
   );
   gpc1_1 gpc2328 (
      {stage6_15[6]},
      {stage7_15[2]}
   );
   gpc1_1 gpc2329 (
      {stage6_15[7]},
      {stage7_15[3]}
   );
   gpc1_1 gpc2330 (
      {stage6_17[0]},
      {stage7_17[2]}
   );
   gpc1_1 gpc2331 (
      {stage6_17[1]},
      {stage7_17[3]}
   );
   gpc1_1 gpc2332 (
      {stage6_17[2]},
      {stage7_17[4]}
   );
   gpc1_1 gpc2333 (
      {stage6_17[3]},
      {stage7_17[5]}
   );
   gpc1_1 gpc2334 (
      {stage6_17[4]},
      {stage7_17[6]}
   );
   gpc1_1 gpc2335 (
      {stage6_18[6]},
      {stage7_18[2]}
   );
   gpc1_1 gpc2336 (
      {stage6_20[6]},
      {stage7_20[2]}
   );
   gpc1_1 gpc2337 (
      {stage6_20[7]},
      {stage7_20[3]}
   );
   gpc1_1 gpc2338 (
      {stage6_21[4]},
      {stage7_21[2]}
   );
   gpc1_1 gpc2339 (
      {stage6_22[1]},
      {stage7_22[2]}
   );
   gpc1_1 gpc2340 (
      {stage6_23[0]},
      {stage7_23[1]}
   );
   gpc615_5 gpc2341 (
      {stage7_0[0], stage7_0[1], stage7_0[2], stage7_0[3], stage7_0[4]},
      {stage7_1[0]},
      {stage7_2[0], stage7_2[1], stage7_2[2], stage7_2[3], stage7_2[4], 1'b0},
      {stage8_4[0],stage8_3[0],stage8_2[0],stage8_1[0],stage8_0[0]}
   );
   gpc7_3 gpc2342 (
      {stage7_4[0], stage7_4[1], stage7_4[2], stage7_4[3], stage7_4[4], stage7_4[5], stage7_4[6]},
      {stage8_6[0],stage8_5[0],stage8_4[1]}
   );
   gpc615_5 gpc2343 (
      {stage7_5[0], stage7_5[1], stage7_5[2], 1'b0, 1'b0},
      {stage7_6[0]},
      {stage7_7[0], stage7_7[1], stage7_7[2], stage7_7[3], stage7_7[4], stage7_7[5]},
      {stage8_9[0],stage8_8[0],stage8_7[0],stage8_6[1],stage8_5[1]}
   );
   gpc23_3 gpc2344 (
      {stage7_9[0], stage7_9[1], stage7_9[2]},
      {stage7_10[0], stage7_10[1]},
      {stage8_11[0],stage8_10[0],stage8_9[1]}
   );
   gpc135_4 gpc2345 (
      {stage7_10[2], stage7_10[3], stage7_10[4], stage7_10[5], stage7_10[6]},
      {stage7_11[0], stage7_11[1], stage7_11[2]},
      {stage7_12[0]},
      {stage8_13[0],stage8_12[0],stage8_11[1],stage8_10[1]}
   );
   gpc1343_5 gpc2346 (
      {stage7_13[0], stage7_13[1], stage7_13[2]},
      {stage7_14[0], stage7_14[1], stage7_14[2], stage7_14[3]},
      {stage7_15[0], stage7_15[1], stage7_15[2]},
      {stage7_16[0]},
      {stage8_17[0],stage8_16[0],stage8_15[0],stage8_14[0],stage8_13[1]}
   );
   gpc7_3 gpc2347 (
      {stage7_17[0], stage7_17[1], stage7_17[2], stage7_17[3], stage7_17[4], stage7_17[5], stage7_17[6]},
      {stage8_19[0],stage8_18[0],stage8_17[1]}
   );
   gpc1325_5 gpc2348 (
      {stage7_18[0], stage7_18[1], stage7_18[2], 1'b0, 1'b0},
      {stage7_19[0], stage7_19[1]},
      {stage7_20[0], stage7_20[1], stage7_20[2]},
      {stage7_21[0]},
      {stage8_22[0],stage8_21[0],stage8_20[0],stage8_19[1],stage8_18[1]}
   );
   gpc1163_5 gpc2349 (
      {stage7_21[1], stage7_21[2], 1'b0},
      {stage7_22[0], stage7_22[1], stage7_22[2], 1'b0, 1'b0, 1'b0},
      {stage7_23[0]},
      {1'b0},
      {stage8_24[0],stage8_23[0],stage8_22[1],stage8_21[1]}
   );
   gpc1_1 gpc2350 (
      {stage7_0[5]},
      {stage8_0[1]}
   );
   gpc1_1 gpc2351 (
      {stage7_1[1]},
      {stage8_1[1]}
   );
   gpc1_1 gpc2352 (
      {stage7_3[0]},
      {stage8_3[1]}
   );
   gpc1_1 gpc2353 (
      {stage7_8[0]},
      {stage8_8[1]}
   );
   gpc1_1 gpc2354 (
      {stage7_12[1]},
      {stage8_12[1]}
   );
   gpc1_1 gpc2355 (
      {stage7_14[4]},
      {stage8_14[1]}
   );
   gpc1_1 gpc2356 (
      {stage7_15[3]},
      {stage8_15[1]}
   );
   gpc1_1 gpc2357 (
      {stage7_16[1]},
      {stage8_16[1]}
   );
   gpc1_1 gpc2358 (
      {stage7_20[3]},
      {stage8_20[1]}
   );
   gpc1_1 gpc2359 (
      {stage7_23[1]},
      {stage8_23[1]}
   );
endmodule

module testbench();
    reg [511:0] src0;
    reg [511:0] src1;
    reg [511:0] src2;
    reg [511:0] src3;
    reg [511:0] src4;
    reg [511:0] src5;
    reg [511:0] src6;
    reg [511:0] src7;
    reg [511:0] src8;
    reg [511:0] src9;
    reg [511:0] src10;
    reg [511:0] src11;
    reg [511:0] src12;
    reg [511:0] src13;
    reg [511:0] src14;
    reg [511:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [24:0] srcsum;
    wire [24:0] dstsum;
    wire test;
    compressor_CLA512_16 compressor_CLA512_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161] + src0[162] + src0[163] + src0[164] + src0[165] + src0[166] + src0[167] + src0[168] + src0[169] + src0[170] + src0[171] + src0[172] + src0[173] + src0[174] + src0[175] + src0[176] + src0[177] + src0[178] + src0[179] + src0[180] + src0[181] + src0[182] + src0[183] + src0[184] + src0[185] + src0[186] + src0[187] + src0[188] + src0[189] + src0[190] + src0[191] + src0[192] + src0[193] + src0[194] + src0[195] + src0[196] + src0[197] + src0[198] + src0[199] + src0[200] + src0[201] + src0[202] + src0[203] + src0[204] + src0[205] + src0[206] + src0[207] + src0[208] + src0[209] + src0[210] + src0[211] + src0[212] + src0[213] + src0[214] + src0[215] + src0[216] + src0[217] + src0[218] + src0[219] + src0[220] + src0[221] + src0[222] + src0[223] + src0[224] + src0[225] + src0[226] + src0[227] + src0[228] + src0[229] + src0[230] + src0[231] + src0[232] + src0[233] + src0[234] + src0[235] + src0[236] + src0[237] + src0[238] + src0[239] + src0[240] + src0[241] + src0[242] + src0[243] + src0[244] + src0[245] + src0[246] + src0[247] + src0[248] + src0[249] + src0[250] + src0[251] + src0[252] + src0[253] + src0[254] + src0[255] + src0[256] + src0[257] + src0[258] + src0[259] + src0[260] + src0[261] + src0[262] + src0[263] + src0[264] + src0[265] + src0[266] + src0[267] + src0[268] + src0[269] + src0[270] + src0[271] + src0[272] + src0[273] + src0[274] + src0[275] + src0[276] + src0[277] + src0[278] + src0[279] + src0[280] + src0[281] + src0[282] + src0[283] + src0[284] + src0[285] + src0[286] + src0[287] + src0[288] + src0[289] + src0[290] + src0[291] + src0[292] + src0[293] + src0[294] + src0[295] + src0[296] + src0[297] + src0[298] + src0[299] + src0[300] + src0[301] + src0[302] + src0[303] + src0[304] + src0[305] + src0[306] + src0[307] + src0[308] + src0[309] + src0[310] + src0[311] + src0[312] + src0[313] + src0[314] + src0[315] + src0[316] + src0[317] + src0[318] + src0[319] + src0[320] + src0[321] + src0[322] + src0[323] + src0[324] + src0[325] + src0[326] + src0[327] + src0[328] + src0[329] + src0[330] + src0[331] + src0[332] + src0[333] + src0[334] + src0[335] + src0[336] + src0[337] + src0[338] + src0[339] + src0[340] + src0[341] + src0[342] + src0[343] + src0[344] + src0[345] + src0[346] + src0[347] + src0[348] + src0[349] + src0[350] + src0[351] + src0[352] + src0[353] + src0[354] + src0[355] + src0[356] + src0[357] + src0[358] + src0[359] + src0[360] + src0[361] + src0[362] + src0[363] + src0[364] + src0[365] + src0[366] + src0[367] + src0[368] + src0[369] + src0[370] + src0[371] + src0[372] + src0[373] + src0[374] + src0[375] + src0[376] + src0[377] + src0[378] + src0[379] + src0[380] + src0[381] + src0[382] + src0[383] + src0[384] + src0[385] + src0[386] + src0[387] + src0[388] + src0[389] + src0[390] + src0[391] + src0[392] + src0[393] + src0[394] + src0[395] + src0[396] + src0[397] + src0[398] + src0[399] + src0[400] + src0[401] + src0[402] + src0[403] + src0[404] + src0[405] + src0[406] + src0[407] + src0[408] + src0[409] + src0[410] + src0[411] + src0[412] + src0[413] + src0[414] + src0[415] + src0[416] + src0[417] + src0[418] + src0[419] + src0[420] + src0[421] + src0[422] + src0[423] + src0[424] + src0[425] + src0[426] + src0[427] + src0[428] + src0[429] + src0[430] + src0[431] + src0[432] + src0[433] + src0[434] + src0[435] + src0[436] + src0[437] + src0[438] + src0[439] + src0[440] + src0[441] + src0[442] + src0[443] + src0[444] + src0[445] + src0[446] + src0[447] + src0[448] + src0[449] + src0[450] + src0[451] + src0[452] + src0[453] + src0[454] + src0[455] + src0[456] + src0[457] + src0[458] + src0[459] + src0[460] + src0[461] + src0[462] + src0[463] + src0[464] + src0[465] + src0[466] + src0[467] + src0[468] + src0[469] + src0[470] + src0[471] + src0[472] + src0[473] + src0[474] + src0[475] + src0[476] + src0[477] + src0[478] + src0[479] + src0[480] + src0[481] + src0[482] + src0[483] + src0[484] + src0[485] + src0[486] + src0[487] + src0[488] + src0[489] + src0[490] + src0[491] + src0[492] + src0[493] + src0[494] + src0[495] + src0[496] + src0[497] + src0[498] + src0[499] + src0[500] + src0[501] + src0[502] + src0[503] + src0[504] + src0[505] + src0[506] + src0[507] + src0[508] + src0[509] + src0[510] + src0[511])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161] + src1[162] + src1[163] + src1[164] + src1[165] + src1[166] + src1[167] + src1[168] + src1[169] + src1[170] + src1[171] + src1[172] + src1[173] + src1[174] + src1[175] + src1[176] + src1[177] + src1[178] + src1[179] + src1[180] + src1[181] + src1[182] + src1[183] + src1[184] + src1[185] + src1[186] + src1[187] + src1[188] + src1[189] + src1[190] + src1[191] + src1[192] + src1[193] + src1[194] + src1[195] + src1[196] + src1[197] + src1[198] + src1[199] + src1[200] + src1[201] + src1[202] + src1[203] + src1[204] + src1[205] + src1[206] + src1[207] + src1[208] + src1[209] + src1[210] + src1[211] + src1[212] + src1[213] + src1[214] + src1[215] + src1[216] + src1[217] + src1[218] + src1[219] + src1[220] + src1[221] + src1[222] + src1[223] + src1[224] + src1[225] + src1[226] + src1[227] + src1[228] + src1[229] + src1[230] + src1[231] + src1[232] + src1[233] + src1[234] + src1[235] + src1[236] + src1[237] + src1[238] + src1[239] + src1[240] + src1[241] + src1[242] + src1[243] + src1[244] + src1[245] + src1[246] + src1[247] + src1[248] + src1[249] + src1[250] + src1[251] + src1[252] + src1[253] + src1[254] + src1[255] + src1[256] + src1[257] + src1[258] + src1[259] + src1[260] + src1[261] + src1[262] + src1[263] + src1[264] + src1[265] + src1[266] + src1[267] + src1[268] + src1[269] + src1[270] + src1[271] + src1[272] + src1[273] + src1[274] + src1[275] + src1[276] + src1[277] + src1[278] + src1[279] + src1[280] + src1[281] + src1[282] + src1[283] + src1[284] + src1[285] + src1[286] + src1[287] + src1[288] + src1[289] + src1[290] + src1[291] + src1[292] + src1[293] + src1[294] + src1[295] + src1[296] + src1[297] + src1[298] + src1[299] + src1[300] + src1[301] + src1[302] + src1[303] + src1[304] + src1[305] + src1[306] + src1[307] + src1[308] + src1[309] + src1[310] + src1[311] + src1[312] + src1[313] + src1[314] + src1[315] + src1[316] + src1[317] + src1[318] + src1[319] + src1[320] + src1[321] + src1[322] + src1[323] + src1[324] + src1[325] + src1[326] + src1[327] + src1[328] + src1[329] + src1[330] + src1[331] + src1[332] + src1[333] + src1[334] + src1[335] + src1[336] + src1[337] + src1[338] + src1[339] + src1[340] + src1[341] + src1[342] + src1[343] + src1[344] + src1[345] + src1[346] + src1[347] + src1[348] + src1[349] + src1[350] + src1[351] + src1[352] + src1[353] + src1[354] + src1[355] + src1[356] + src1[357] + src1[358] + src1[359] + src1[360] + src1[361] + src1[362] + src1[363] + src1[364] + src1[365] + src1[366] + src1[367] + src1[368] + src1[369] + src1[370] + src1[371] + src1[372] + src1[373] + src1[374] + src1[375] + src1[376] + src1[377] + src1[378] + src1[379] + src1[380] + src1[381] + src1[382] + src1[383] + src1[384] + src1[385] + src1[386] + src1[387] + src1[388] + src1[389] + src1[390] + src1[391] + src1[392] + src1[393] + src1[394] + src1[395] + src1[396] + src1[397] + src1[398] + src1[399] + src1[400] + src1[401] + src1[402] + src1[403] + src1[404] + src1[405] + src1[406] + src1[407] + src1[408] + src1[409] + src1[410] + src1[411] + src1[412] + src1[413] + src1[414] + src1[415] + src1[416] + src1[417] + src1[418] + src1[419] + src1[420] + src1[421] + src1[422] + src1[423] + src1[424] + src1[425] + src1[426] + src1[427] + src1[428] + src1[429] + src1[430] + src1[431] + src1[432] + src1[433] + src1[434] + src1[435] + src1[436] + src1[437] + src1[438] + src1[439] + src1[440] + src1[441] + src1[442] + src1[443] + src1[444] + src1[445] + src1[446] + src1[447] + src1[448] + src1[449] + src1[450] + src1[451] + src1[452] + src1[453] + src1[454] + src1[455] + src1[456] + src1[457] + src1[458] + src1[459] + src1[460] + src1[461] + src1[462] + src1[463] + src1[464] + src1[465] + src1[466] + src1[467] + src1[468] + src1[469] + src1[470] + src1[471] + src1[472] + src1[473] + src1[474] + src1[475] + src1[476] + src1[477] + src1[478] + src1[479] + src1[480] + src1[481] + src1[482] + src1[483] + src1[484] + src1[485] + src1[486] + src1[487] + src1[488] + src1[489] + src1[490] + src1[491] + src1[492] + src1[493] + src1[494] + src1[495] + src1[496] + src1[497] + src1[498] + src1[499] + src1[500] + src1[501] + src1[502] + src1[503] + src1[504] + src1[505] + src1[506] + src1[507] + src1[508] + src1[509] + src1[510] + src1[511])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161] + src2[162] + src2[163] + src2[164] + src2[165] + src2[166] + src2[167] + src2[168] + src2[169] + src2[170] + src2[171] + src2[172] + src2[173] + src2[174] + src2[175] + src2[176] + src2[177] + src2[178] + src2[179] + src2[180] + src2[181] + src2[182] + src2[183] + src2[184] + src2[185] + src2[186] + src2[187] + src2[188] + src2[189] + src2[190] + src2[191] + src2[192] + src2[193] + src2[194] + src2[195] + src2[196] + src2[197] + src2[198] + src2[199] + src2[200] + src2[201] + src2[202] + src2[203] + src2[204] + src2[205] + src2[206] + src2[207] + src2[208] + src2[209] + src2[210] + src2[211] + src2[212] + src2[213] + src2[214] + src2[215] + src2[216] + src2[217] + src2[218] + src2[219] + src2[220] + src2[221] + src2[222] + src2[223] + src2[224] + src2[225] + src2[226] + src2[227] + src2[228] + src2[229] + src2[230] + src2[231] + src2[232] + src2[233] + src2[234] + src2[235] + src2[236] + src2[237] + src2[238] + src2[239] + src2[240] + src2[241] + src2[242] + src2[243] + src2[244] + src2[245] + src2[246] + src2[247] + src2[248] + src2[249] + src2[250] + src2[251] + src2[252] + src2[253] + src2[254] + src2[255] + src2[256] + src2[257] + src2[258] + src2[259] + src2[260] + src2[261] + src2[262] + src2[263] + src2[264] + src2[265] + src2[266] + src2[267] + src2[268] + src2[269] + src2[270] + src2[271] + src2[272] + src2[273] + src2[274] + src2[275] + src2[276] + src2[277] + src2[278] + src2[279] + src2[280] + src2[281] + src2[282] + src2[283] + src2[284] + src2[285] + src2[286] + src2[287] + src2[288] + src2[289] + src2[290] + src2[291] + src2[292] + src2[293] + src2[294] + src2[295] + src2[296] + src2[297] + src2[298] + src2[299] + src2[300] + src2[301] + src2[302] + src2[303] + src2[304] + src2[305] + src2[306] + src2[307] + src2[308] + src2[309] + src2[310] + src2[311] + src2[312] + src2[313] + src2[314] + src2[315] + src2[316] + src2[317] + src2[318] + src2[319] + src2[320] + src2[321] + src2[322] + src2[323] + src2[324] + src2[325] + src2[326] + src2[327] + src2[328] + src2[329] + src2[330] + src2[331] + src2[332] + src2[333] + src2[334] + src2[335] + src2[336] + src2[337] + src2[338] + src2[339] + src2[340] + src2[341] + src2[342] + src2[343] + src2[344] + src2[345] + src2[346] + src2[347] + src2[348] + src2[349] + src2[350] + src2[351] + src2[352] + src2[353] + src2[354] + src2[355] + src2[356] + src2[357] + src2[358] + src2[359] + src2[360] + src2[361] + src2[362] + src2[363] + src2[364] + src2[365] + src2[366] + src2[367] + src2[368] + src2[369] + src2[370] + src2[371] + src2[372] + src2[373] + src2[374] + src2[375] + src2[376] + src2[377] + src2[378] + src2[379] + src2[380] + src2[381] + src2[382] + src2[383] + src2[384] + src2[385] + src2[386] + src2[387] + src2[388] + src2[389] + src2[390] + src2[391] + src2[392] + src2[393] + src2[394] + src2[395] + src2[396] + src2[397] + src2[398] + src2[399] + src2[400] + src2[401] + src2[402] + src2[403] + src2[404] + src2[405] + src2[406] + src2[407] + src2[408] + src2[409] + src2[410] + src2[411] + src2[412] + src2[413] + src2[414] + src2[415] + src2[416] + src2[417] + src2[418] + src2[419] + src2[420] + src2[421] + src2[422] + src2[423] + src2[424] + src2[425] + src2[426] + src2[427] + src2[428] + src2[429] + src2[430] + src2[431] + src2[432] + src2[433] + src2[434] + src2[435] + src2[436] + src2[437] + src2[438] + src2[439] + src2[440] + src2[441] + src2[442] + src2[443] + src2[444] + src2[445] + src2[446] + src2[447] + src2[448] + src2[449] + src2[450] + src2[451] + src2[452] + src2[453] + src2[454] + src2[455] + src2[456] + src2[457] + src2[458] + src2[459] + src2[460] + src2[461] + src2[462] + src2[463] + src2[464] + src2[465] + src2[466] + src2[467] + src2[468] + src2[469] + src2[470] + src2[471] + src2[472] + src2[473] + src2[474] + src2[475] + src2[476] + src2[477] + src2[478] + src2[479] + src2[480] + src2[481] + src2[482] + src2[483] + src2[484] + src2[485] + src2[486] + src2[487] + src2[488] + src2[489] + src2[490] + src2[491] + src2[492] + src2[493] + src2[494] + src2[495] + src2[496] + src2[497] + src2[498] + src2[499] + src2[500] + src2[501] + src2[502] + src2[503] + src2[504] + src2[505] + src2[506] + src2[507] + src2[508] + src2[509] + src2[510] + src2[511])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161] + src3[162] + src3[163] + src3[164] + src3[165] + src3[166] + src3[167] + src3[168] + src3[169] + src3[170] + src3[171] + src3[172] + src3[173] + src3[174] + src3[175] + src3[176] + src3[177] + src3[178] + src3[179] + src3[180] + src3[181] + src3[182] + src3[183] + src3[184] + src3[185] + src3[186] + src3[187] + src3[188] + src3[189] + src3[190] + src3[191] + src3[192] + src3[193] + src3[194] + src3[195] + src3[196] + src3[197] + src3[198] + src3[199] + src3[200] + src3[201] + src3[202] + src3[203] + src3[204] + src3[205] + src3[206] + src3[207] + src3[208] + src3[209] + src3[210] + src3[211] + src3[212] + src3[213] + src3[214] + src3[215] + src3[216] + src3[217] + src3[218] + src3[219] + src3[220] + src3[221] + src3[222] + src3[223] + src3[224] + src3[225] + src3[226] + src3[227] + src3[228] + src3[229] + src3[230] + src3[231] + src3[232] + src3[233] + src3[234] + src3[235] + src3[236] + src3[237] + src3[238] + src3[239] + src3[240] + src3[241] + src3[242] + src3[243] + src3[244] + src3[245] + src3[246] + src3[247] + src3[248] + src3[249] + src3[250] + src3[251] + src3[252] + src3[253] + src3[254] + src3[255] + src3[256] + src3[257] + src3[258] + src3[259] + src3[260] + src3[261] + src3[262] + src3[263] + src3[264] + src3[265] + src3[266] + src3[267] + src3[268] + src3[269] + src3[270] + src3[271] + src3[272] + src3[273] + src3[274] + src3[275] + src3[276] + src3[277] + src3[278] + src3[279] + src3[280] + src3[281] + src3[282] + src3[283] + src3[284] + src3[285] + src3[286] + src3[287] + src3[288] + src3[289] + src3[290] + src3[291] + src3[292] + src3[293] + src3[294] + src3[295] + src3[296] + src3[297] + src3[298] + src3[299] + src3[300] + src3[301] + src3[302] + src3[303] + src3[304] + src3[305] + src3[306] + src3[307] + src3[308] + src3[309] + src3[310] + src3[311] + src3[312] + src3[313] + src3[314] + src3[315] + src3[316] + src3[317] + src3[318] + src3[319] + src3[320] + src3[321] + src3[322] + src3[323] + src3[324] + src3[325] + src3[326] + src3[327] + src3[328] + src3[329] + src3[330] + src3[331] + src3[332] + src3[333] + src3[334] + src3[335] + src3[336] + src3[337] + src3[338] + src3[339] + src3[340] + src3[341] + src3[342] + src3[343] + src3[344] + src3[345] + src3[346] + src3[347] + src3[348] + src3[349] + src3[350] + src3[351] + src3[352] + src3[353] + src3[354] + src3[355] + src3[356] + src3[357] + src3[358] + src3[359] + src3[360] + src3[361] + src3[362] + src3[363] + src3[364] + src3[365] + src3[366] + src3[367] + src3[368] + src3[369] + src3[370] + src3[371] + src3[372] + src3[373] + src3[374] + src3[375] + src3[376] + src3[377] + src3[378] + src3[379] + src3[380] + src3[381] + src3[382] + src3[383] + src3[384] + src3[385] + src3[386] + src3[387] + src3[388] + src3[389] + src3[390] + src3[391] + src3[392] + src3[393] + src3[394] + src3[395] + src3[396] + src3[397] + src3[398] + src3[399] + src3[400] + src3[401] + src3[402] + src3[403] + src3[404] + src3[405] + src3[406] + src3[407] + src3[408] + src3[409] + src3[410] + src3[411] + src3[412] + src3[413] + src3[414] + src3[415] + src3[416] + src3[417] + src3[418] + src3[419] + src3[420] + src3[421] + src3[422] + src3[423] + src3[424] + src3[425] + src3[426] + src3[427] + src3[428] + src3[429] + src3[430] + src3[431] + src3[432] + src3[433] + src3[434] + src3[435] + src3[436] + src3[437] + src3[438] + src3[439] + src3[440] + src3[441] + src3[442] + src3[443] + src3[444] + src3[445] + src3[446] + src3[447] + src3[448] + src3[449] + src3[450] + src3[451] + src3[452] + src3[453] + src3[454] + src3[455] + src3[456] + src3[457] + src3[458] + src3[459] + src3[460] + src3[461] + src3[462] + src3[463] + src3[464] + src3[465] + src3[466] + src3[467] + src3[468] + src3[469] + src3[470] + src3[471] + src3[472] + src3[473] + src3[474] + src3[475] + src3[476] + src3[477] + src3[478] + src3[479] + src3[480] + src3[481] + src3[482] + src3[483] + src3[484] + src3[485] + src3[486] + src3[487] + src3[488] + src3[489] + src3[490] + src3[491] + src3[492] + src3[493] + src3[494] + src3[495] + src3[496] + src3[497] + src3[498] + src3[499] + src3[500] + src3[501] + src3[502] + src3[503] + src3[504] + src3[505] + src3[506] + src3[507] + src3[508] + src3[509] + src3[510] + src3[511])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161] + src4[162] + src4[163] + src4[164] + src4[165] + src4[166] + src4[167] + src4[168] + src4[169] + src4[170] + src4[171] + src4[172] + src4[173] + src4[174] + src4[175] + src4[176] + src4[177] + src4[178] + src4[179] + src4[180] + src4[181] + src4[182] + src4[183] + src4[184] + src4[185] + src4[186] + src4[187] + src4[188] + src4[189] + src4[190] + src4[191] + src4[192] + src4[193] + src4[194] + src4[195] + src4[196] + src4[197] + src4[198] + src4[199] + src4[200] + src4[201] + src4[202] + src4[203] + src4[204] + src4[205] + src4[206] + src4[207] + src4[208] + src4[209] + src4[210] + src4[211] + src4[212] + src4[213] + src4[214] + src4[215] + src4[216] + src4[217] + src4[218] + src4[219] + src4[220] + src4[221] + src4[222] + src4[223] + src4[224] + src4[225] + src4[226] + src4[227] + src4[228] + src4[229] + src4[230] + src4[231] + src4[232] + src4[233] + src4[234] + src4[235] + src4[236] + src4[237] + src4[238] + src4[239] + src4[240] + src4[241] + src4[242] + src4[243] + src4[244] + src4[245] + src4[246] + src4[247] + src4[248] + src4[249] + src4[250] + src4[251] + src4[252] + src4[253] + src4[254] + src4[255] + src4[256] + src4[257] + src4[258] + src4[259] + src4[260] + src4[261] + src4[262] + src4[263] + src4[264] + src4[265] + src4[266] + src4[267] + src4[268] + src4[269] + src4[270] + src4[271] + src4[272] + src4[273] + src4[274] + src4[275] + src4[276] + src4[277] + src4[278] + src4[279] + src4[280] + src4[281] + src4[282] + src4[283] + src4[284] + src4[285] + src4[286] + src4[287] + src4[288] + src4[289] + src4[290] + src4[291] + src4[292] + src4[293] + src4[294] + src4[295] + src4[296] + src4[297] + src4[298] + src4[299] + src4[300] + src4[301] + src4[302] + src4[303] + src4[304] + src4[305] + src4[306] + src4[307] + src4[308] + src4[309] + src4[310] + src4[311] + src4[312] + src4[313] + src4[314] + src4[315] + src4[316] + src4[317] + src4[318] + src4[319] + src4[320] + src4[321] + src4[322] + src4[323] + src4[324] + src4[325] + src4[326] + src4[327] + src4[328] + src4[329] + src4[330] + src4[331] + src4[332] + src4[333] + src4[334] + src4[335] + src4[336] + src4[337] + src4[338] + src4[339] + src4[340] + src4[341] + src4[342] + src4[343] + src4[344] + src4[345] + src4[346] + src4[347] + src4[348] + src4[349] + src4[350] + src4[351] + src4[352] + src4[353] + src4[354] + src4[355] + src4[356] + src4[357] + src4[358] + src4[359] + src4[360] + src4[361] + src4[362] + src4[363] + src4[364] + src4[365] + src4[366] + src4[367] + src4[368] + src4[369] + src4[370] + src4[371] + src4[372] + src4[373] + src4[374] + src4[375] + src4[376] + src4[377] + src4[378] + src4[379] + src4[380] + src4[381] + src4[382] + src4[383] + src4[384] + src4[385] + src4[386] + src4[387] + src4[388] + src4[389] + src4[390] + src4[391] + src4[392] + src4[393] + src4[394] + src4[395] + src4[396] + src4[397] + src4[398] + src4[399] + src4[400] + src4[401] + src4[402] + src4[403] + src4[404] + src4[405] + src4[406] + src4[407] + src4[408] + src4[409] + src4[410] + src4[411] + src4[412] + src4[413] + src4[414] + src4[415] + src4[416] + src4[417] + src4[418] + src4[419] + src4[420] + src4[421] + src4[422] + src4[423] + src4[424] + src4[425] + src4[426] + src4[427] + src4[428] + src4[429] + src4[430] + src4[431] + src4[432] + src4[433] + src4[434] + src4[435] + src4[436] + src4[437] + src4[438] + src4[439] + src4[440] + src4[441] + src4[442] + src4[443] + src4[444] + src4[445] + src4[446] + src4[447] + src4[448] + src4[449] + src4[450] + src4[451] + src4[452] + src4[453] + src4[454] + src4[455] + src4[456] + src4[457] + src4[458] + src4[459] + src4[460] + src4[461] + src4[462] + src4[463] + src4[464] + src4[465] + src4[466] + src4[467] + src4[468] + src4[469] + src4[470] + src4[471] + src4[472] + src4[473] + src4[474] + src4[475] + src4[476] + src4[477] + src4[478] + src4[479] + src4[480] + src4[481] + src4[482] + src4[483] + src4[484] + src4[485] + src4[486] + src4[487] + src4[488] + src4[489] + src4[490] + src4[491] + src4[492] + src4[493] + src4[494] + src4[495] + src4[496] + src4[497] + src4[498] + src4[499] + src4[500] + src4[501] + src4[502] + src4[503] + src4[504] + src4[505] + src4[506] + src4[507] + src4[508] + src4[509] + src4[510] + src4[511])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161] + src5[162] + src5[163] + src5[164] + src5[165] + src5[166] + src5[167] + src5[168] + src5[169] + src5[170] + src5[171] + src5[172] + src5[173] + src5[174] + src5[175] + src5[176] + src5[177] + src5[178] + src5[179] + src5[180] + src5[181] + src5[182] + src5[183] + src5[184] + src5[185] + src5[186] + src5[187] + src5[188] + src5[189] + src5[190] + src5[191] + src5[192] + src5[193] + src5[194] + src5[195] + src5[196] + src5[197] + src5[198] + src5[199] + src5[200] + src5[201] + src5[202] + src5[203] + src5[204] + src5[205] + src5[206] + src5[207] + src5[208] + src5[209] + src5[210] + src5[211] + src5[212] + src5[213] + src5[214] + src5[215] + src5[216] + src5[217] + src5[218] + src5[219] + src5[220] + src5[221] + src5[222] + src5[223] + src5[224] + src5[225] + src5[226] + src5[227] + src5[228] + src5[229] + src5[230] + src5[231] + src5[232] + src5[233] + src5[234] + src5[235] + src5[236] + src5[237] + src5[238] + src5[239] + src5[240] + src5[241] + src5[242] + src5[243] + src5[244] + src5[245] + src5[246] + src5[247] + src5[248] + src5[249] + src5[250] + src5[251] + src5[252] + src5[253] + src5[254] + src5[255] + src5[256] + src5[257] + src5[258] + src5[259] + src5[260] + src5[261] + src5[262] + src5[263] + src5[264] + src5[265] + src5[266] + src5[267] + src5[268] + src5[269] + src5[270] + src5[271] + src5[272] + src5[273] + src5[274] + src5[275] + src5[276] + src5[277] + src5[278] + src5[279] + src5[280] + src5[281] + src5[282] + src5[283] + src5[284] + src5[285] + src5[286] + src5[287] + src5[288] + src5[289] + src5[290] + src5[291] + src5[292] + src5[293] + src5[294] + src5[295] + src5[296] + src5[297] + src5[298] + src5[299] + src5[300] + src5[301] + src5[302] + src5[303] + src5[304] + src5[305] + src5[306] + src5[307] + src5[308] + src5[309] + src5[310] + src5[311] + src5[312] + src5[313] + src5[314] + src5[315] + src5[316] + src5[317] + src5[318] + src5[319] + src5[320] + src5[321] + src5[322] + src5[323] + src5[324] + src5[325] + src5[326] + src5[327] + src5[328] + src5[329] + src5[330] + src5[331] + src5[332] + src5[333] + src5[334] + src5[335] + src5[336] + src5[337] + src5[338] + src5[339] + src5[340] + src5[341] + src5[342] + src5[343] + src5[344] + src5[345] + src5[346] + src5[347] + src5[348] + src5[349] + src5[350] + src5[351] + src5[352] + src5[353] + src5[354] + src5[355] + src5[356] + src5[357] + src5[358] + src5[359] + src5[360] + src5[361] + src5[362] + src5[363] + src5[364] + src5[365] + src5[366] + src5[367] + src5[368] + src5[369] + src5[370] + src5[371] + src5[372] + src5[373] + src5[374] + src5[375] + src5[376] + src5[377] + src5[378] + src5[379] + src5[380] + src5[381] + src5[382] + src5[383] + src5[384] + src5[385] + src5[386] + src5[387] + src5[388] + src5[389] + src5[390] + src5[391] + src5[392] + src5[393] + src5[394] + src5[395] + src5[396] + src5[397] + src5[398] + src5[399] + src5[400] + src5[401] + src5[402] + src5[403] + src5[404] + src5[405] + src5[406] + src5[407] + src5[408] + src5[409] + src5[410] + src5[411] + src5[412] + src5[413] + src5[414] + src5[415] + src5[416] + src5[417] + src5[418] + src5[419] + src5[420] + src5[421] + src5[422] + src5[423] + src5[424] + src5[425] + src5[426] + src5[427] + src5[428] + src5[429] + src5[430] + src5[431] + src5[432] + src5[433] + src5[434] + src5[435] + src5[436] + src5[437] + src5[438] + src5[439] + src5[440] + src5[441] + src5[442] + src5[443] + src5[444] + src5[445] + src5[446] + src5[447] + src5[448] + src5[449] + src5[450] + src5[451] + src5[452] + src5[453] + src5[454] + src5[455] + src5[456] + src5[457] + src5[458] + src5[459] + src5[460] + src5[461] + src5[462] + src5[463] + src5[464] + src5[465] + src5[466] + src5[467] + src5[468] + src5[469] + src5[470] + src5[471] + src5[472] + src5[473] + src5[474] + src5[475] + src5[476] + src5[477] + src5[478] + src5[479] + src5[480] + src5[481] + src5[482] + src5[483] + src5[484] + src5[485] + src5[486] + src5[487] + src5[488] + src5[489] + src5[490] + src5[491] + src5[492] + src5[493] + src5[494] + src5[495] + src5[496] + src5[497] + src5[498] + src5[499] + src5[500] + src5[501] + src5[502] + src5[503] + src5[504] + src5[505] + src5[506] + src5[507] + src5[508] + src5[509] + src5[510] + src5[511])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161] + src6[162] + src6[163] + src6[164] + src6[165] + src6[166] + src6[167] + src6[168] + src6[169] + src6[170] + src6[171] + src6[172] + src6[173] + src6[174] + src6[175] + src6[176] + src6[177] + src6[178] + src6[179] + src6[180] + src6[181] + src6[182] + src6[183] + src6[184] + src6[185] + src6[186] + src6[187] + src6[188] + src6[189] + src6[190] + src6[191] + src6[192] + src6[193] + src6[194] + src6[195] + src6[196] + src6[197] + src6[198] + src6[199] + src6[200] + src6[201] + src6[202] + src6[203] + src6[204] + src6[205] + src6[206] + src6[207] + src6[208] + src6[209] + src6[210] + src6[211] + src6[212] + src6[213] + src6[214] + src6[215] + src6[216] + src6[217] + src6[218] + src6[219] + src6[220] + src6[221] + src6[222] + src6[223] + src6[224] + src6[225] + src6[226] + src6[227] + src6[228] + src6[229] + src6[230] + src6[231] + src6[232] + src6[233] + src6[234] + src6[235] + src6[236] + src6[237] + src6[238] + src6[239] + src6[240] + src6[241] + src6[242] + src6[243] + src6[244] + src6[245] + src6[246] + src6[247] + src6[248] + src6[249] + src6[250] + src6[251] + src6[252] + src6[253] + src6[254] + src6[255] + src6[256] + src6[257] + src6[258] + src6[259] + src6[260] + src6[261] + src6[262] + src6[263] + src6[264] + src6[265] + src6[266] + src6[267] + src6[268] + src6[269] + src6[270] + src6[271] + src6[272] + src6[273] + src6[274] + src6[275] + src6[276] + src6[277] + src6[278] + src6[279] + src6[280] + src6[281] + src6[282] + src6[283] + src6[284] + src6[285] + src6[286] + src6[287] + src6[288] + src6[289] + src6[290] + src6[291] + src6[292] + src6[293] + src6[294] + src6[295] + src6[296] + src6[297] + src6[298] + src6[299] + src6[300] + src6[301] + src6[302] + src6[303] + src6[304] + src6[305] + src6[306] + src6[307] + src6[308] + src6[309] + src6[310] + src6[311] + src6[312] + src6[313] + src6[314] + src6[315] + src6[316] + src6[317] + src6[318] + src6[319] + src6[320] + src6[321] + src6[322] + src6[323] + src6[324] + src6[325] + src6[326] + src6[327] + src6[328] + src6[329] + src6[330] + src6[331] + src6[332] + src6[333] + src6[334] + src6[335] + src6[336] + src6[337] + src6[338] + src6[339] + src6[340] + src6[341] + src6[342] + src6[343] + src6[344] + src6[345] + src6[346] + src6[347] + src6[348] + src6[349] + src6[350] + src6[351] + src6[352] + src6[353] + src6[354] + src6[355] + src6[356] + src6[357] + src6[358] + src6[359] + src6[360] + src6[361] + src6[362] + src6[363] + src6[364] + src6[365] + src6[366] + src6[367] + src6[368] + src6[369] + src6[370] + src6[371] + src6[372] + src6[373] + src6[374] + src6[375] + src6[376] + src6[377] + src6[378] + src6[379] + src6[380] + src6[381] + src6[382] + src6[383] + src6[384] + src6[385] + src6[386] + src6[387] + src6[388] + src6[389] + src6[390] + src6[391] + src6[392] + src6[393] + src6[394] + src6[395] + src6[396] + src6[397] + src6[398] + src6[399] + src6[400] + src6[401] + src6[402] + src6[403] + src6[404] + src6[405] + src6[406] + src6[407] + src6[408] + src6[409] + src6[410] + src6[411] + src6[412] + src6[413] + src6[414] + src6[415] + src6[416] + src6[417] + src6[418] + src6[419] + src6[420] + src6[421] + src6[422] + src6[423] + src6[424] + src6[425] + src6[426] + src6[427] + src6[428] + src6[429] + src6[430] + src6[431] + src6[432] + src6[433] + src6[434] + src6[435] + src6[436] + src6[437] + src6[438] + src6[439] + src6[440] + src6[441] + src6[442] + src6[443] + src6[444] + src6[445] + src6[446] + src6[447] + src6[448] + src6[449] + src6[450] + src6[451] + src6[452] + src6[453] + src6[454] + src6[455] + src6[456] + src6[457] + src6[458] + src6[459] + src6[460] + src6[461] + src6[462] + src6[463] + src6[464] + src6[465] + src6[466] + src6[467] + src6[468] + src6[469] + src6[470] + src6[471] + src6[472] + src6[473] + src6[474] + src6[475] + src6[476] + src6[477] + src6[478] + src6[479] + src6[480] + src6[481] + src6[482] + src6[483] + src6[484] + src6[485] + src6[486] + src6[487] + src6[488] + src6[489] + src6[490] + src6[491] + src6[492] + src6[493] + src6[494] + src6[495] + src6[496] + src6[497] + src6[498] + src6[499] + src6[500] + src6[501] + src6[502] + src6[503] + src6[504] + src6[505] + src6[506] + src6[507] + src6[508] + src6[509] + src6[510] + src6[511])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161] + src7[162] + src7[163] + src7[164] + src7[165] + src7[166] + src7[167] + src7[168] + src7[169] + src7[170] + src7[171] + src7[172] + src7[173] + src7[174] + src7[175] + src7[176] + src7[177] + src7[178] + src7[179] + src7[180] + src7[181] + src7[182] + src7[183] + src7[184] + src7[185] + src7[186] + src7[187] + src7[188] + src7[189] + src7[190] + src7[191] + src7[192] + src7[193] + src7[194] + src7[195] + src7[196] + src7[197] + src7[198] + src7[199] + src7[200] + src7[201] + src7[202] + src7[203] + src7[204] + src7[205] + src7[206] + src7[207] + src7[208] + src7[209] + src7[210] + src7[211] + src7[212] + src7[213] + src7[214] + src7[215] + src7[216] + src7[217] + src7[218] + src7[219] + src7[220] + src7[221] + src7[222] + src7[223] + src7[224] + src7[225] + src7[226] + src7[227] + src7[228] + src7[229] + src7[230] + src7[231] + src7[232] + src7[233] + src7[234] + src7[235] + src7[236] + src7[237] + src7[238] + src7[239] + src7[240] + src7[241] + src7[242] + src7[243] + src7[244] + src7[245] + src7[246] + src7[247] + src7[248] + src7[249] + src7[250] + src7[251] + src7[252] + src7[253] + src7[254] + src7[255] + src7[256] + src7[257] + src7[258] + src7[259] + src7[260] + src7[261] + src7[262] + src7[263] + src7[264] + src7[265] + src7[266] + src7[267] + src7[268] + src7[269] + src7[270] + src7[271] + src7[272] + src7[273] + src7[274] + src7[275] + src7[276] + src7[277] + src7[278] + src7[279] + src7[280] + src7[281] + src7[282] + src7[283] + src7[284] + src7[285] + src7[286] + src7[287] + src7[288] + src7[289] + src7[290] + src7[291] + src7[292] + src7[293] + src7[294] + src7[295] + src7[296] + src7[297] + src7[298] + src7[299] + src7[300] + src7[301] + src7[302] + src7[303] + src7[304] + src7[305] + src7[306] + src7[307] + src7[308] + src7[309] + src7[310] + src7[311] + src7[312] + src7[313] + src7[314] + src7[315] + src7[316] + src7[317] + src7[318] + src7[319] + src7[320] + src7[321] + src7[322] + src7[323] + src7[324] + src7[325] + src7[326] + src7[327] + src7[328] + src7[329] + src7[330] + src7[331] + src7[332] + src7[333] + src7[334] + src7[335] + src7[336] + src7[337] + src7[338] + src7[339] + src7[340] + src7[341] + src7[342] + src7[343] + src7[344] + src7[345] + src7[346] + src7[347] + src7[348] + src7[349] + src7[350] + src7[351] + src7[352] + src7[353] + src7[354] + src7[355] + src7[356] + src7[357] + src7[358] + src7[359] + src7[360] + src7[361] + src7[362] + src7[363] + src7[364] + src7[365] + src7[366] + src7[367] + src7[368] + src7[369] + src7[370] + src7[371] + src7[372] + src7[373] + src7[374] + src7[375] + src7[376] + src7[377] + src7[378] + src7[379] + src7[380] + src7[381] + src7[382] + src7[383] + src7[384] + src7[385] + src7[386] + src7[387] + src7[388] + src7[389] + src7[390] + src7[391] + src7[392] + src7[393] + src7[394] + src7[395] + src7[396] + src7[397] + src7[398] + src7[399] + src7[400] + src7[401] + src7[402] + src7[403] + src7[404] + src7[405] + src7[406] + src7[407] + src7[408] + src7[409] + src7[410] + src7[411] + src7[412] + src7[413] + src7[414] + src7[415] + src7[416] + src7[417] + src7[418] + src7[419] + src7[420] + src7[421] + src7[422] + src7[423] + src7[424] + src7[425] + src7[426] + src7[427] + src7[428] + src7[429] + src7[430] + src7[431] + src7[432] + src7[433] + src7[434] + src7[435] + src7[436] + src7[437] + src7[438] + src7[439] + src7[440] + src7[441] + src7[442] + src7[443] + src7[444] + src7[445] + src7[446] + src7[447] + src7[448] + src7[449] + src7[450] + src7[451] + src7[452] + src7[453] + src7[454] + src7[455] + src7[456] + src7[457] + src7[458] + src7[459] + src7[460] + src7[461] + src7[462] + src7[463] + src7[464] + src7[465] + src7[466] + src7[467] + src7[468] + src7[469] + src7[470] + src7[471] + src7[472] + src7[473] + src7[474] + src7[475] + src7[476] + src7[477] + src7[478] + src7[479] + src7[480] + src7[481] + src7[482] + src7[483] + src7[484] + src7[485] + src7[486] + src7[487] + src7[488] + src7[489] + src7[490] + src7[491] + src7[492] + src7[493] + src7[494] + src7[495] + src7[496] + src7[497] + src7[498] + src7[499] + src7[500] + src7[501] + src7[502] + src7[503] + src7[504] + src7[505] + src7[506] + src7[507] + src7[508] + src7[509] + src7[510] + src7[511])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161] + src8[162] + src8[163] + src8[164] + src8[165] + src8[166] + src8[167] + src8[168] + src8[169] + src8[170] + src8[171] + src8[172] + src8[173] + src8[174] + src8[175] + src8[176] + src8[177] + src8[178] + src8[179] + src8[180] + src8[181] + src8[182] + src8[183] + src8[184] + src8[185] + src8[186] + src8[187] + src8[188] + src8[189] + src8[190] + src8[191] + src8[192] + src8[193] + src8[194] + src8[195] + src8[196] + src8[197] + src8[198] + src8[199] + src8[200] + src8[201] + src8[202] + src8[203] + src8[204] + src8[205] + src8[206] + src8[207] + src8[208] + src8[209] + src8[210] + src8[211] + src8[212] + src8[213] + src8[214] + src8[215] + src8[216] + src8[217] + src8[218] + src8[219] + src8[220] + src8[221] + src8[222] + src8[223] + src8[224] + src8[225] + src8[226] + src8[227] + src8[228] + src8[229] + src8[230] + src8[231] + src8[232] + src8[233] + src8[234] + src8[235] + src8[236] + src8[237] + src8[238] + src8[239] + src8[240] + src8[241] + src8[242] + src8[243] + src8[244] + src8[245] + src8[246] + src8[247] + src8[248] + src8[249] + src8[250] + src8[251] + src8[252] + src8[253] + src8[254] + src8[255] + src8[256] + src8[257] + src8[258] + src8[259] + src8[260] + src8[261] + src8[262] + src8[263] + src8[264] + src8[265] + src8[266] + src8[267] + src8[268] + src8[269] + src8[270] + src8[271] + src8[272] + src8[273] + src8[274] + src8[275] + src8[276] + src8[277] + src8[278] + src8[279] + src8[280] + src8[281] + src8[282] + src8[283] + src8[284] + src8[285] + src8[286] + src8[287] + src8[288] + src8[289] + src8[290] + src8[291] + src8[292] + src8[293] + src8[294] + src8[295] + src8[296] + src8[297] + src8[298] + src8[299] + src8[300] + src8[301] + src8[302] + src8[303] + src8[304] + src8[305] + src8[306] + src8[307] + src8[308] + src8[309] + src8[310] + src8[311] + src8[312] + src8[313] + src8[314] + src8[315] + src8[316] + src8[317] + src8[318] + src8[319] + src8[320] + src8[321] + src8[322] + src8[323] + src8[324] + src8[325] + src8[326] + src8[327] + src8[328] + src8[329] + src8[330] + src8[331] + src8[332] + src8[333] + src8[334] + src8[335] + src8[336] + src8[337] + src8[338] + src8[339] + src8[340] + src8[341] + src8[342] + src8[343] + src8[344] + src8[345] + src8[346] + src8[347] + src8[348] + src8[349] + src8[350] + src8[351] + src8[352] + src8[353] + src8[354] + src8[355] + src8[356] + src8[357] + src8[358] + src8[359] + src8[360] + src8[361] + src8[362] + src8[363] + src8[364] + src8[365] + src8[366] + src8[367] + src8[368] + src8[369] + src8[370] + src8[371] + src8[372] + src8[373] + src8[374] + src8[375] + src8[376] + src8[377] + src8[378] + src8[379] + src8[380] + src8[381] + src8[382] + src8[383] + src8[384] + src8[385] + src8[386] + src8[387] + src8[388] + src8[389] + src8[390] + src8[391] + src8[392] + src8[393] + src8[394] + src8[395] + src8[396] + src8[397] + src8[398] + src8[399] + src8[400] + src8[401] + src8[402] + src8[403] + src8[404] + src8[405] + src8[406] + src8[407] + src8[408] + src8[409] + src8[410] + src8[411] + src8[412] + src8[413] + src8[414] + src8[415] + src8[416] + src8[417] + src8[418] + src8[419] + src8[420] + src8[421] + src8[422] + src8[423] + src8[424] + src8[425] + src8[426] + src8[427] + src8[428] + src8[429] + src8[430] + src8[431] + src8[432] + src8[433] + src8[434] + src8[435] + src8[436] + src8[437] + src8[438] + src8[439] + src8[440] + src8[441] + src8[442] + src8[443] + src8[444] + src8[445] + src8[446] + src8[447] + src8[448] + src8[449] + src8[450] + src8[451] + src8[452] + src8[453] + src8[454] + src8[455] + src8[456] + src8[457] + src8[458] + src8[459] + src8[460] + src8[461] + src8[462] + src8[463] + src8[464] + src8[465] + src8[466] + src8[467] + src8[468] + src8[469] + src8[470] + src8[471] + src8[472] + src8[473] + src8[474] + src8[475] + src8[476] + src8[477] + src8[478] + src8[479] + src8[480] + src8[481] + src8[482] + src8[483] + src8[484] + src8[485] + src8[486] + src8[487] + src8[488] + src8[489] + src8[490] + src8[491] + src8[492] + src8[493] + src8[494] + src8[495] + src8[496] + src8[497] + src8[498] + src8[499] + src8[500] + src8[501] + src8[502] + src8[503] + src8[504] + src8[505] + src8[506] + src8[507] + src8[508] + src8[509] + src8[510] + src8[511])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161] + src9[162] + src9[163] + src9[164] + src9[165] + src9[166] + src9[167] + src9[168] + src9[169] + src9[170] + src9[171] + src9[172] + src9[173] + src9[174] + src9[175] + src9[176] + src9[177] + src9[178] + src9[179] + src9[180] + src9[181] + src9[182] + src9[183] + src9[184] + src9[185] + src9[186] + src9[187] + src9[188] + src9[189] + src9[190] + src9[191] + src9[192] + src9[193] + src9[194] + src9[195] + src9[196] + src9[197] + src9[198] + src9[199] + src9[200] + src9[201] + src9[202] + src9[203] + src9[204] + src9[205] + src9[206] + src9[207] + src9[208] + src9[209] + src9[210] + src9[211] + src9[212] + src9[213] + src9[214] + src9[215] + src9[216] + src9[217] + src9[218] + src9[219] + src9[220] + src9[221] + src9[222] + src9[223] + src9[224] + src9[225] + src9[226] + src9[227] + src9[228] + src9[229] + src9[230] + src9[231] + src9[232] + src9[233] + src9[234] + src9[235] + src9[236] + src9[237] + src9[238] + src9[239] + src9[240] + src9[241] + src9[242] + src9[243] + src9[244] + src9[245] + src9[246] + src9[247] + src9[248] + src9[249] + src9[250] + src9[251] + src9[252] + src9[253] + src9[254] + src9[255] + src9[256] + src9[257] + src9[258] + src9[259] + src9[260] + src9[261] + src9[262] + src9[263] + src9[264] + src9[265] + src9[266] + src9[267] + src9[268] + src9[269] + src9[270] + src9[271] + src9[272] + src9[273] + src9[274] + src9[275] + src9[276] + src9[277] + src9[278] + src9[279] + src9[280] + src9[281] + src9[282] + src9[283] + src9[284] + src9[285] + src9[286] + src9[287] + src9[288] + src9[289] + src9[290] + src9[291] + src9[292] + src9[293] + src9[294] + src9[295] + src9[296] + src9[297] + src9[298] + src9[299] + src9[300] + src9[301] + src9[302] + src9[303] + src9[304] + src9[305] + src9[306] + src9[307] + src9[308] + src9[309] + src9[310] + src9[311] + src9[312] + src9[313] + src9[314] + src9[315] + src9[316] + src9[317] + src9[318] + src9[319] + src9[320] + src9[321] + src9[322] + src9[323] + src9[324] + src9[325] + src9[326] + src9[327] + src9[328] + src9[329] + src9[330] + src9[331] + src9[332] + src9[333] + src9[334] + src9[335] + src9[336] + src9[337] + src9[338] + src9[339] + src9[340] + src9[341] + src9[342] + src9[343] + src9[344] + src9[345] + src9[346] + src9[347] + src9[348] + src9[349] + src9[350] + src9[351] + src9[352] + src9[353] + src9[354] + src9[355] + src9[356] + src9[357] + src9[358] + src9[359] + src9[360] + src9[361] + src9[362] + src9[363] + src9[364] + src9[365] + src9[366] + src9[367] + src9[368] + src9[369] + src9[370] + src9[371] + src9[372] + src9[373] + src9[374] + src9[375] + src9[376] + src9[377] + src9[378] + src9[379] + src9[380] + src9[381] + src9[382] + src9[383] + src9[384] + src9[385] + src9[386] + src9[387] + src9[388] + src9[389] + src9[390] + src9[391] + src9[392] + src9[393] + src9[394] + src9[395] + src9[396] + src9[397] + src9[398] + src9[399] + src9[400] + src9[401] + src9[402] + src9[403] + src9[404] + src9[405] + src9[406] + src9[407] + src9[408] + src9[409] + src9[410] + src9[411] + src9[412] + src9[413] + src9[414] + src9[415] + src9[416] + src9[417] + src9[418] + src9[419] + src9[420] + src9[421] + src9[422] + src9[423] + src9[424] + src9[425] + src9[426] + src9[427] + src9[428] + src9[429] + src9[430] + src9[431] + src9[432] + src9[433] + src9[434] + src9[435] + src9[436] + src9[437] + src9[438] + src9[439] + src9[440] + src9[441] + src9[442] + src9[443] + src9[444] + src9[445] + src9[446] + src9[447] + src9[448] + src9[449] + src9[450] + src9[451] + src9[452] + src9[453] + src9[454] + src9[455] + src9[456] + src9[457] + src9[458] + src9[459] + src9[460] + src9[461] + src9[462] + src9[463] + src9[464] + src9[465] + src9[466] + src9[467] + src9[468] + src9[469] + src9[470] + src9[471] + src9[472] + src9[473] + src9[474] + src9[475] + src9[476] + src9[477] + src9[478] + src9[479] + src9[480] + src9[481] + src9[482] + src9[483] + src9[484] + src9[485] + src9[486] + src9[487] + src9[488] + src9[489] + src9[490] + src9[491] + src9[492] + src9[493] + src9[494] + src9[495] + src9[496] + src9[497] + src9[498] + src9[499] + src9[500] + src9[501] + src9[502] + src9[503] + src9[504] + src9[505] + src9[506] + src9[507] + src9[508] + src9[509] + src9[510] + src9[511])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161] + src10[162] + src10[163] + src10[164] + src10[165] + src10[166] + src10[167] + src10[168] + src10[169] + src10[170] + src10[171] + src10[172] + src10[173] + src10[174] + src10[175] + src10[176] + src10[177] + src10[178] + src10[179] + src10[180] + src10[181] + src10[182] + src10[183] + src10[184] + src10[185] + src10[186] + src10[187] + src10[188] + src10[189] + src10[190] + src10[191] + src10[192] + src10[193] + src10[194] + src10[195] + src10[196] + src10[197] + src10[198] + src10[199] + src10[200] + src10[201] + src10[202] + src10[203] + src10[204] + src10[205] + src10[206] + src10[207] + src10[208] + src10[209] + src10[210] + src10[211] + src10[212] + src10[213] + src10[214] + src10[215] + src10[216] + src10[217] + src10[218] + src10[219] + src10[220] + src10[221] + src10[222] + src10[223] + src10[224] + src10[225] + src10[226] + src10[227] + src10[228] + src10[229] + src10[230] + src10[231] + src10[232] + src10[233] + src10[234] + src10[235] + src10[236] + src10[237] + src10[238] + src10[239] + src10[240] + src10[241] + src10[242] + src10[243] + src10[244] + src10[245] + src10[246] + src10[247] + src10[248] + src10[249] + src10[250] + src10[251] + src10[252] + src10[253] + src10[254] + src10[255] + src10[256] + src10[257] + src10[258] + src10[259] + src10[260] + src10[261] + src10[262] + src10[263] + src10[264] + src10[265] + src10[266] + src10[267] + src10[268] + src10[269] + src10[270] + src10[271] + src10[272] + src10[273] + src10[274] + src10[275] + src10[276] + src10[277] + src10[278] + src10[279] + src10[280] + src10[281] + src10[282] + src10[283] + src10[284] + src10[285] + src10[286] + src10[287] + src10[288] + src10[289] + src10[290] + src10[291] + src10[292] + src10[293] + src10[294] + src10[295] + src10[296] + src10[297] + src10[298] + src10[299] + src10[300] + src10[301] + src10[302] + src10[303] + src10[304] + src10[305] + src10[306] + src10[307] + src10[308] + src10[309] + src10[310] + src10[311] + src10[312] + src10[313] + src10[314] + src10[315] + src10[316] + src10[317] + src10[318] + src10[319] + src10[320] + src10[321] + src10[322] + src10[323] + src10[324] + src10[325] + src10[326] + src10[327] + src10[328] + src10[329] + src10[330] + src10[331] + src10[332] + src10[333] + src10[334] + src10[335] + src10[336] + src10[337] + src10[338] + src10[339] + src10[340] + src10[341] + src10[342] + src10[343] + src10[344] + src10[345] + src10[346] + src10[347] + src10[348] + src10[349] + src10[350] + src10[351] + src10[352] + src10[353] + src10[354] + src10[355] + src10[356] + src10[357] + src10[358] + src10[359] + src10[360] + src10[361] + src10[362] + src10[363] + src10[364] + src10[365] + src10[366] + src10[367] + src10[368] + src10[369] + src10[370] + src10[371] + src10[372] + src10[373] + src10[374] + src10[375] + src10[376] + src10[377] + src10[378] + src10[379] + src10[380] + src10[381] + src10[382] + src10[383] + src10[384] + src10[385] + src10[386] + src10[387] + src10[388] + src10[389] + src10[390] + src10[391] + src10[392] + src10[393] + src10[394] + src10[395] + src10[396] + src10[397] + src10[398] + src10[399] + src10[400] + src10[401] + src10[402] + src10[403] + src10[404] + src10[405] + src10[406] + src10[407] + src10[408] + src10[409] + src10[410] + src10[411] + src10[412] + src10[413] + src10[414] + src10[415] + src10[416] + src10[417] + src10[418] + src10[419] + src10[420] + src10[421] + src10[422] + src10[423] + src10[424] + src10[425] + src10[426] + src10[427] + src10[428] + src10[429] + src10[430] + src10[431] + src10[432] + src10[433] + src10[434] + src10[435] + src10[436] + src10[437] + src10[438] + src10[439] + src10[440] + src10[441] + src10[442] + src10[443] + src10[444] + src10[445] + src10[446] + src10[447] + src10[448] + src10[449] + src10[450] + src10[451] + src10[452] + src10[453] + src10[454] + src10[455] + src10[456] + src10[457] + src10[458] + src10[459] + src10[460] + src10[461] + src10[462] + src10[463] + src10[464] + src10[465] + src10[466] + src10[467] + src10[468] + src10[469] + src10[470] + src10[471] + src10[472] + src10[473] + src10[474] + src10[475] + src10[476] + src10[477] + src10[478] + src10[479] + src10[480] + src10[481] + src10[482] + src10[483] + src10[484] + src10[485] + src10[486] + src10[487] + src10[488] + src10[489] + src10[490] + src10[491] + src10[492] + src10[493] + src10[494] + src10[495] + src10[496] + src10[497] + src10[498] + src10[499] + src10[500] + src10[501] + src10[502] + src10[503] + src10[504] + src10[505] + src10[506] + src10[507] + src10[508] + src10[509] + src10[510] + src10[511])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161] + src11[162] + src11[163] + src11[164] + src11[165] + src11[166] + src11[167] + src11[168] + src11[169] + src11[170] + src11[171] + src11[172] + src11[173] + src11[174] + src11[175] + src11[176] + src11[177] + src11[178] + src11[179] + src11[180] + src11[181] + src11[182] + src11[183] + src11[184] + src11[185] + src11[186] + src11[187] + src11[188] + src11[189] + src11[190] + src11[191] + src11[192] + src11[193] + src11[194] + src11[195] + src11[196] + src11[197] + src11[198] + src11[199] + src11[200] + src11[201] + src11[202] + src11[203] + src11[204] + src11[205] + src11[206] + src11[207] + src11[208] + src11[209] + src11[210] + src11[211] + src11[212] + src11[213] + src11[214] + src11[215] + src11[216] + src11[217] + src11[218] + src11[219] + src11[220] + src11[221] + src11[222] + src11[223] + src11[224] + src11[225] + src11[226] + src11[227] + src11[228] + src11[229] + src11[230] + src11[231] + src11[232] + src11[233] + src11[234] + src11[235] + src11[236] + src11[237] + src11[238] + src11[239] + src11[240] + src11[241] + src11[242] + src11[243] + src11[244] + src11[245] + src11[246] + src11[247] + src11[248] + src11[249] + src11[250] + src11[251] + src11[252] + src11[253] + src11[254] + src11[255] + src11[256] + src11[257] + src11[258] + src11[259] + src11[260] + src11[261] + src11[262] + src11[263] + src11[264] + src11[265] + src11[266] + src11[267] + src11[268] + src11[269] + src11[270] + src11[271] + src11[272] + src11[273] + src11[274] + src11[275] + src11[276] + src11[277] + src11[278] + src11[279] + src11[280] + src11[281] + src11[282] + src11[283] + src11[284] + src11[285] + src11[286] + src11[287] + src11[288] + src11[289] + src11[290] + src11[291] + src11[292] + src11[293] + src11[294] + src11[295] + src11[296] + src11[297] + src11[298] + src11[299] + src11[300] + src11[301] + src11[302] + src11[303] + src11[304] + src11[305] + src11[306] + src11[307] + src11[308] + src11[309] + src11[310] + src11[311] + src11[312] + src11[313] + src11[314] + src11[315] + src11[316] + src11[317] + src11[318] + src11[319] + src11[320] + src11[321] + src11[322] + src11[323] + src11[324] + src11[325] + src11[326] + src11[327] + src11[328] + src11[329] + src11[330] + src11[331] + src11[332] + src11[333] + src11[334] + src11[335] + src11[336] + src11[337] + src11[338] + src11[339] + src11[340] + src11[341] + src11[342] + src11[343] + src11[344] + src11[345] + src11[346] + src11[347] + src11[348] + src11[349] + src11[350] + src11[351] + src11[352] + src11[353] + src11[354] + src11[355] + src11[356] + src11[357] + src11[358] + src11[359] + src11[360] + src11[361] + src11[362] + src11[363] + src11[364] + src11[365] + src11[366] + src11[367] + src11[368] + src11[369] + src11[370] + src11[371] + src11[372] + src11[373] + src11[374] + src11[375] + src11[376] + src11[377] + src11[378] + src11[379] + src11[380] + src11[381] + src11[382] + src11[383] + src11[384] + src11[385] + src11[386] + src11[387] + src11[388] + src11[389] + src11[390] + src11[391] + src11[392] + src11[393] + src11[394] + src11[395] + src11[396] + src11[397] + src11[398] + src11[399] + src11[400] + src11[401] + src11[402] + src11[403] + src11[404] + src11[405] + src11[406] + src11[407] + src11[408] + src11[409] + src11[410] + src11[411] + src11[412] + src11[413] + src11[414] + src11[415] + src11[416] + src11[417] + src11[418] + src11[419] + src11[420] + src11[421] + src11[422] + src11[423] + src11[424] + src11[425] + src11[426] + src11[427] + src11[428] + src11[429] + src11[430] + src11[431] + src11[432] + src11[433] + src11[434] + src11[435] + src11[436] + src11[437] + src11[438] + src11[439] + src11[440] + src11[441] + src11[442] + src11[443] + src11[444] + src11[445] + src11[446] + src11[447] + src11[448] + src11[449] + src11[450] + src11[451] + src11[452] + src11[453] + src11[454] + src11[455] + src11[456] + src11[457] + src11[458] + src11[459] + src11[460] + src11[461] + src11[462] + src11[463] + src11[464] + src11[465] + src11[466] + src11[467] + src11[468] + src11[469] + src11[470] + src11[471] + src11[472] + src11[473] + src11[474] + src11[475] + src11[476] + src11[477] + src11[478] + src11[479] + src11[480] + src11[481] + src11[482] + src11[483] + src11[484] + src11[485] + src11[486] + src11[487] + src11[488] + src11[489] + src11[490] + src11[491] + src11[492] + src11[493] + src11[494] + src11[495] + src11[496] + src11[497] + src11[498] + src11[499] + src11[500] + src11[501] + src11[502] + src11[503] + src11[504] + src11[505] + src11[506] + src11[507] + src11[508] + src11[509] + src11[510] + src11[511])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161] + src12[162] + src12[163] + src12[164] + src12[165] + src12[166] + src12[167] + src12[168] + src12[169] + src12[170] + src12[171] + src12[172] + src12[173] + src12[174] + src12[175] + src12[176] + src12[177] + src12[178] + src12[179] + src12[180] + src12[181] + src12[182] + src12[183] + src12[184] + src12[185] + src12[186] + src12[187] + src12[188] + src12[189] + src12[190] + src12[191] + src12[192] + src12[193] + src12[194] + src12[195] + src12[196] + src12[197] + src12[198] + src12[199] + src12[200] + src12[201] + src12[202] + src12[203] + src12[204] + src12[205] + src12[206] + src12[207] + src12[208] + src12[209] + src12[210] + src12[211] + src12[212] + src12[213] + src12[214] + src12[215] + src12[216] + src12[217] + src12[218] + src12[219] + src12[220] + src12[221] + src12[222] + src12[223] + src12[224] + src12[225] + src12[226] + src12[227] + src12[228] + src12[229] + src12[230] + src12[231] + src12[232] + src12[233] + src12[234] + src12[235] + src12[236] + src12[237] + src12[238] + src12[239] + src12[240] + src12[241] + src12[242] + src12[243] + src12[244] + src12[245] + src12[246] + src12[247] + src12[248] + src12[249] + src12[250] + src12[251] + src12[252] + src12[253] + src12[254] + src12[255] + src12[256] + src12[257] + src12[258] + src12[259] + src12[260] + src12[261] + src12[262] + src12[263] + src12[264] + src12[265] + src12[266] + src12[267] + src12[268] + src12[269] + src12[270] + src12[271] + src12[272] + src12[273] + src12[274] + src12[275] + src12[276] + src12[277] + src12[278] + src12[279] + src12[280] + src12[281] + src12[282] + src12[283] + src12[284] + src12[285] + src12[286] + src12[287] + src12[288] + src12[289] + src12[290] + src12[291] + src12[292] + src12[293] + src12[294] + src12[295] + src12[296] + src12[297] + src12[298] + src12[299] + src12[300] + src12[301] + src12[302] + src12[303] + src12[304] + src12[305] + src12[306] + src12[307] + src12[308] + src12[309] + src12[310] + src12[311] + src12[312] + src12[313] + src12[314] + src12[315] + src12[316] + src12[317] + src12[318] + src12[319] + src12[320] + src12[321] + src12[322] + src12[323] + src12[324] + src12[325] + src12[326] + src12[327] + src12[328] + src12[329] + src12[330] + src12[331] + src12[332] + src12[333] + src12[334] + src12[335] + src12[336] + src12[337] + src12[338] + src12[339] + src12[340] + src12[341] + src12[342] + src12[343] + src12[344] + src12[345] + src12[346] + src12[347] + src12[348] + src12[349] + src12[350] + src12[351] + src12[352] + src12[353] + src12[354] + src12[355] + src12[356] + src12[357] + src12[358] + src12[359] + src12[360] + src12[361] + src12[362] + src12[363] + src12[364] + src12[365] + src12[366] + src12[367] + src12[368] + src12[369] + src12[370] + src12[371] + src12[372] + src12[373] + src12[374] + src12[375] + src12[376] + src12[377] + src12[378] + src12[379] + src12[380] + src12[381] + src12[382] + src12[383] + src12[384] + src12[385] + src12[386] + src12[387] + src12[388] + src12[389] + src12[390] + src12[391] + src12[392] + src12[393] + src12[394] + src12[395] + src12[396] + src12[397] + src12[398] + src12[399] + src12[400] + src12[401] + src12[402] + src12[403] + src12[404] + src12[405] + src12[406] + src12[407] + src12[408] + src12[409] + src12[410] + src12[411] + src12[412] + src12[413] + src12[414] + src12[415] + src12[416] + src12[417] + src12[418] + src12[419] + src12[420] + src12[421] + src12[422] + src12[423] + src12[424] + src12[425] + src12[426] + src12[427] + src12[428] + src12[429] + src12[430] + src12[431] + src12[432] + src12[433] + src12[434] + src12[435] + src12[436] + src12[437] + src12[438] + src12[439] + src12[440] + src12[441] + src12[442] + src12[443] + src12[444] + src12[445] + src12[446] + src12[447] + src12[448] + src12[449] + src12[450] + src12[451] + src12[452] + src12[453] + src12[454] + src12[455] + src12[456] + src12[457] + src12[458] + src12[459] + src12[460] + src12[461] + src12[462] + src12[463] + src12[464] + src12[465] + src12[466] + src12[467] + src12[468] + src12[469] + src12[470] + src12[471] + src12[472] + src12[473] + src12[474] + src12[475] + src12[476] + src12[477] + src12[478] + src12[479] + src12[480] + src12[481] + src12[482] + src12[483] + src12[484] + src12[485] + src12[486] + src12[487] + src12[488] + src12[489] + src12[490] + src12[491] + src12[492] + src12[493] + src12[494] + src12[495] + src12[496] + src12[497] + src12[498] + src12[499] + src12[500] + src12[501] + src12[502] + src12[503] + src12[504] + src12[505] + src12[506] + src12[507] + src12[508] + src12[509] + src12[510] + src12[511])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161] + src13[162] + src13[163] + src13[164] + src13[165] + src13[166] + src13[167] + src13[168] + src13[169] + src13[170] + src13[171] + src13[172] + src13[173] + src13[174] + src13[175] + src13[176] + src13[177] + src13[178] + src13[179] + src13[180] + src13[181] + src13[182] + src13[183] + src13[184] + src13[185] + src13[186] + src13[187] + src13[188] + src13[189] + src13[190] + src13[191] + src13[192] + src13[193] + src13[194] + src13[195] + src13[196] + src13[197] + src13[198] + src13[199] + src13[200] + src13[201] + src13[202] + src13[203] + src13[204] + src13[205] + src13[206] + src13[207] + src13[208] + src13[209] + src13[210] + src13[211] + src13[212] + src13[213] + src13[214] + src13[215] + src13[216] + src13[217] + src13[218] + src13[219] + src13[220] + src13[221] + src13[222] + src13[223] + src13[224] + src13[225] + src13[226] + src13[227] + src13[228] + src13[229] + src13[230] + src13[231] + src13[232] + src13[233] + src13[234] + src13[235] + src13[236] + src13[237] + src13[238] + src13[239] + src13[240] + src13[241] + src13[242] + src13[243] + src13[244] + src13[245] + src13[246] + src13[247] + src13[248] + src13[249] + src13[250] + src13[251] + src13[252] + src13[253] + src13[254] + src13[255] + src13[256] + src13[257] + src13[258] + src13[259] + src13[260] + src13[261] + src13[262] + src13[263] + src13[264] + src13[265] + src13[266] + src13[267] + src13[268] + src13[269] + src13[270] + src13[271] + src13[272] + src13[273] + src13[274] + src13[275] + src13[276] + src13[277] + src13[278] + src13[279] + src13[280] + src13[281] + src13[282] + src13[283] + src13[284] + src13[285] + src13[286] + src13[287] + src13[288] + src13[289] + src13[290] + src13[291] + src13[292] + src13[293] + src13[294] + src13[295] + src13[296] + src13[297] + src13[298] + src13[299] + src13[300] + src13[301] + src13[302] + src13[303] + src13[304] + src13[305] + src13[306] + src13[307] + src13[308] + src13[309] + src13[310] + src13[311] + src13[312] + src13[313] + src13[314] + src13[315] + src13[316] + src13[317] + src13[318] + src13[319] + src13[320] + src13[321] + src13[322] + src13[323] + src13[324] + src13[325] + src13[326] + src13[327] + src13[328] + src13[329] + src13[330] + src13[331] + src13[332] + src13[333] + src13[334] + src13[335] + src13[336] + src13[337] + src13[338] + src13[339] + src13[340] + src13[341] + src13[342] + src13[343] + src13[344] + src13[345] + src13[346] + src13[347] + src13[348] + src13[349] + src13[350] + src13[351] + src13[352] + src13[353] + src13[354] + src13[355] + src13[356] + src13[357] + src13[358] + src13[359] + src13[360] + src13[361] + src13[362] + src13[363] + src13[364] + src13[365] + src13[366] + src13[367] + src13[368] + src13[369] + src13[370] + src13[371] + src13[372] + src13[373] + src13[374] + src13[375] + src13[376] + src13[377] + src13[378] + src13[379] + src13[380] + src13[381] + src13[382] + src13[383] + src13[384] + src13[385] + src13[386] + src13[387] + src13[388] + src13[389] + src13[390] + src13[391] + src13[392] + src13[393] + src13[394] + src13[395] + src13[396] + src13[397] + src13[398] + src13[399] + src13[400] + src13[401] + src13[402] + src13[403] + src13[404] + src13[405] + src13[406] + src13[407] + src13[408] + src13[409] + src13[410] + src13[411] + src13[412] + src13[413] + src13[414] + src13[415] + src13[416] + src13[417] + src13[418] + src13[419] + src13[420] + src13[421] + src13[422] + src13[423] + src13[424] + src13[425] + src13[426] + src13[427] + src13[428] + src13[429] + src13[430] + src13[431] + src13[432] + src13[433] + src13[434] + src13[435] + src13[436] + src13[437] + src13[438] + src13[439] + src13[440] + src13[441] + src13[442] + src13[443] + src13[444] + src13[445] + src13[446] + src13[447] + src13[448] + src13[449] + src13[450] + src13[451] + src13[452] + src13[453] + src13[454] + src13[455] + src13[456] + src13[457] + src13[458] + src13[459] + src13[460] + src13[461] + src13[462] + src13[463] + src13[464] + src13[465] + src13[466] + src13[467] + src13[468] + src13[469] + src13[470] + src13[471] + src13[472] + src13[473] + src13[474] + src13[475] + src13[476] + src13[477] + src13[478] + src13[479] + src13[480] + src13[481] + src13[482] + src13[483] + src13[484] + src13[485] + src13[486] + src13[487] + src13[488] + src13[489] + src13[490] + src13[491] + src13[492] + src13[493] + src13[494] + src13[495] + src13[496] + src13[497] + src13[498] + src13[499] + src13[500] + src13[501] + src13[502] + src13[503] + src13[504] + src13[505] + src13[506] + src13[507] + src13[508] + src13[509] + src13[510] + src13[511])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161] + src14[162] + src14[163] + src14[164] + src14[165] + src14[166] + src14[167] + src14[168] + src14[169] + src14[170] + src14[171] + src14[172] + src14[173] + src14[174] + src14[175] + src14[176] + src14[177] + src14[178] + src14[179] + src14[180] + src14[181] + src14[182] + src14[183] + src14[184] + src14[185] + src14[186] + src14[187] + src14[188] + src14[189] + src14[190] + src14[191] + src14[192] + src14[193] + src14[194] + src14[195] + src14[196] + src14[197] + src14[198] + src14[199] + src14[200] + src14[201] + src14[202] + src14[203] + src14[204] + src14[205] + src14[206] + src14[207] + src14[208] + src14[209] + src14[210] + src14[211] + src14[212] + src14[213] + src14[214] + src14[215] + src14[216] + src14[217] + src14[218] + src14[219] + src14[220] + src14[221] + src14[222] + src14[223] + src14[224] + src14[225] + src14[226] + src14[227] + src14[228] + src14[229] + src14[230] + src14[231] + src14[232] + src14[233] + src14[234] + src14[235] + src14[236] + src14[237] + src14[238] + src14[239] + src14[240] + src14[241] + src14[242] + src14[243] + src14[244] + src14[245] + src14[246] + src14[247] + src14[248] + src14[249] + src14[250] + src14[251] + src14[252] + src14[253] + src14[254] + src14[255] + src14[256] + src14[257] + src14[258] + src14[259] + src14[260] + src14[261] + src14[262] + src14[263] + src14[264] + src14[265] + src14[266] + src14[267] + src14[268] + src14[269] + src14[270] + src14[271] + src14[272] + src14[273] + src14[274] + src14[275] + src14[276] + src14[277] + src14[278] + src14[279] + src14[280] + src14[281] + src14[282] + src14[283] + src14[284] + src14[285] + src14[286] + src14[287] + src14[288] + src14[289] + src14[290] + src14[291] + src14[292] + src14[293] + src14[294] + src14[295] + src14[296] + src14[297] + src14[298] + src14[299] + src14[300] + src14[301] + src14[302] + src14[303] + src14[304] + src14[305] + src14[306] + src14[307] + src14[308] + src14[309] + src14[310] + src14[311] + src14[312] + src14[313] + src14[314] + src14[315] + src14[316] + src14[317] + src14[318] + src14[319] + src14[320] + src14[321] + src14[322] + src14[323] + src14[324] + src14[325] + src14[326] + src14[327] + src14[328] + src14[329] + src14[330] + src14[331] + src14[332] + src14[333] + src14[334] + src14[335] + src14[336] + src14[337] + src14[338] + src14[339] + src14[340] + src14[341] + src14[342] + src14[343] + src14[344] + src14[345] + src14[346] + src14[347] + src14[348] + src14[349] + src14[350] + src14[351] + src14[352] + src14[353] + src14[354] + src14[355] + src14[356] + src14[357] + src14[358] + src14[359] + src14[360] + src14[361] + src14[362] + src14[363] + src14[364] + src14[365] + src14[366] + src14[367] + src14[368] + src14[369] + src14[370] + src14[371] + src14[372] + src14[373] + src14[374] + src14[375] + src14[376] + src14[377] + src14[378] + src14[379] + src14[380] + src14[381] + src14[382] + src14[383] + src14[384] + src14[385] + src14[386] + src14[387] + src14[388] + src14[389] + src14[390] + src14[391] + src14[392] + src14[393] + src14[394] + src14[395] + src14[396] + src14[397] + src14[398] + src14[399] + src14[400] + src14[401] + src14[402] + src14[403] + src14[404] + src14[405] + src14[406] + src14[407] + src14[408] + src14[409] + src14[410] + src14[411] + src14[412] + src14[413] + src14[414] + src14[415] + src14[416] + src14[417] + src14[418] + src14[419] + src14[420] + src14[421] + src14[422] + src14[423] + src14[424] + src14[425] + src14[426] + src14[427] + src14[428] + src14[429] + src14[430] + src14[431] + src14[432] + src14[433] + src14[434] + src14[435] + src14[436] + src14[437] + src14[438] + src14[439] + src14[440] + src14[441] + src14[442] + src14[443] + src14[444] + src14[445] + src14[446] + src14[447] + src14[448] + src14[449] + src14[450] + src14[451] + src14[452] + src14[453] + src14[454] + src14[455] + src14[456] + src14[457] + src14[458] + src14[459] + src14[460] + src14[461] + src14[462] + src14[463] + src14[464] + src14[465] + src14[466] + src14[467] + src14[468] + src14[469] + src14[470] + src14[471] + src14[472] + src14[473] + src14[474] + src14[475] + src14[476] + src14[477] + src14[478] + src14[479] + src14[480] + src14[481] + src14[482] + src14[483] + src14[484] + src14[485] + src14[486] + src14[487] + src14[488] + src14[489] + src14[490] + src14[491] + src14[492] + src14[493] + src14[494] + src14[495] + src14[496] + src14[497] + src14[498] + src14[499] + src14[500] + src14[501] + src14[502] + src14[503] + src14[504] + src14[505] + src14[506] + src14[507] + src14[508] + src14[509] + src14[510] + src14[511])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161] + src15[162] + src15[163] + src15[164] + src15[165] + src15[166] + src15[167] + src15[168] + src15[169] + src15[170] + src15[171] + src15[172] + src15[173] + src15[174] + src15[175] + src15[176] + src15[177] + src15[178] + src15[179] + src15[180] + src15[181] + src15[182] + src15[183] + src15[184] + src15[185] + src15[186] + src15[187] + src15[188] + src15[189] + src15[190] + src15[191] + src15[192] + src15[193] + src15[194] + src15[195] + src15[196] + src15[197] + src15[198] + src15[199] + src15[200] + src15[201] + src15[202] + src15[203] + src15[204] + src15[205] + src15[206] + src15[207] + src15[208] + src15[209] + src15[210] + src15[211] + src15[212] + src15[213] + src15[214] + src15[215] + src15[216] + src15[217] + src15[218] + src15[219] + src15[220] + src15[221] + src15[222] + src15[223] + src15[224] + src15[225] + src15[226] + src15[227] + src15[228] + src15[229] + src15[230] + src15[231] + src15[232] + src15[233] + src15[234] + src15[235] + src15[236] + src15[237] + src15[238] + src15[239] + src15[240] + src15[241] + src15[242] + src15[243] + src15[244] + src15[245] + src15[246] + src15[247] + src15[248] + src15[249] + src15[250] + src15[251] + src15[252] + src15[253] + src15[254] + src15[255] + src15[256] + src15[257] + src15[258] + src15[259] + src15[260] + src15[261] + src15[262] + src15[263] + src15[264] + src15[265] + src15[266] + src15[267] + src15[268] + src15[269] + src15[270] + src15[271] + src15[272] + src15[273] + src15[274] + src15[275] + src15[276] + src15[277] + src15[278] + src15[279] + src15[280] + src15[281] + src15[282] + src15[283] + src15[284] + src15[285] + src15[286] + src15[287] + src15[288] + src15[289] + src15[290] + src15[291] + src15[292] + src15[293] + src15[294] + src15[295] + src15[296] + src15[297] + src15[298] + src15[299] + src15[300] + src15[301] + src15[302] + src15[303] + src15[304] + src15[305] + src15[306] + src15[307] + src15[308] + src15[309] + src15[310] + src15[311] + src15[312] + src15[313] + src15[314] + src15[315] + src15[316] + src15[317] + src15[318] + src15[319] + src15[320] + src15[321] + src15[322] + src15[323] + src15[324] + src15[325] + src15[326] + src15[327] + src15[328] + src15[329] + src15[330] + src15[331] + src15[332] + src15[333] + src15[334] + src15[335] + src15[336] + src15[337] + src15[338] + src15[339] + src15[340] + src15[341] + src15[342] + src15[343] + src15[344] + src15[345] + src15[346] + src15[347] + src15[348] + src15[349] + src15[350] + src15[351] + src15[352] + src15[353] + src15[354] + src15[355] + src15[356] + src15[357] + src15[358] + src15[359] + src15[360] + src15[361] + src15[362] + src15[363] + src15[364] + src15[365] + src15[366] + src15[367] + src15[368] + src15[369] + src15[370] + src15[371] + src15[372] + src15[373] + src15[374] + src15[375] + src15[376] + src15[377] + src15[378] + src15[379] + src15[380] + src15[381] + src15[382] + src15[383] + src15[384] + src15[385] + src15[386] + src15[387] + src15[388] + src15[389] + src15[390] + src15[391] + src15[392] + src15[393] + src15[394] + src15[395] + src15[396] + src15[397] + src15[398] + src15[399] + src15[400] + src15[401] + src15[402] + src15[403] + src15[404] + src15[405] + src15[406] + src15[407] + src15[408] + src15[409] + src15[410] + src15[411] + src15[412] + src15[413] + src15[414] + src15[415] + src15[416] + src15[417] + src15[418] + src15[419] + src15[420] + src15[421] + src15[422] + src15[423] + src15[424] + src15[425] + src15[426] + src15[427] + src15[428] + src15[429] + src15[430] + src15[431] + src15[432] + src15[433] + src15[434] + src15[435] + src15[436] + src15[437] + src15[438] + src15[439] + src15[440] + src15[441] + src15[442] + src15[443] + src15[444] + src15[445] + src15[446] + src15[447] + src15[448] + src15[449] + src15[450] + src15[451] + src15[452] + src15[453] + src15[454] + src15[455] + src15[456] + src15[457] + src15[458] + src15[459] + src15[460] + src15[461] + src15[462] + src15[463] + src15[464] + src15[465] + src15[466] + src15[467] + src15[468] + src15[469] + src15[470] + src15[471] + src15[472] + src15[473] + src15[474] + src15[475] + src15[476] + src15[477] + src15[478] + src15[479] + src15[480] + src15[481] + src15[482] + src15[483] + src15[484] + src15[485] + src15[486] + src15[487] + src15[488] + src15[489] + src15[490] + src15[491] + src15[492] + src15[493] + src15[494] + src15[495] + src15[496] + src15[497] + src15[498] + src15[499] + src15[500] + src15[501] + src15[502] + src15[503] + src15[504] + src15[505] + src15[506] + src15[507] + src15[508] + src15[509] + src15[510] + src15[511])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he3e528552ebfb77f15906973ccfef3407c84b90f324f981f37fd79988c74759ad9cb10c7c072858d29260a7712fca0f73ea43c55d4f7dc6bd9983e2fde0234721cb698a03d368fe6ae3445d6b456c063a0356f610be3ec0f69f1edb447dfc17c2f0b8cbf83f09aa091e65eaf15fc87cbd60e9e77d726cf58e3239e031e7f363e9b4bebd52ef6d3dccf8a5858660e989782547e8eda98f22fabdb4436a547c87af7824092d63cddb8abbcc6a5530b780c7c570e75d71889269c49e74351f6114fcfbff6043ff1d49208ec37b1417a9f14a06a8c99dc84ccb433f284d5ce1952f989c52bed7c3e3ae6917ca2f400c82f439531cbf6dbaa81b4d02be3159b365fc1ec00e22ec75baa07f97884e12c9a2c95122d49ce833c30f8641b0853201f9913259f504516b7f8dfdc29a947e4d7c071cc7c923e7d0e3a5d8cfe9c16659a2b54952180ad48b687c71eab0bea94014977d2b18a97038c2e49d3eb3dd3c1efc5b22b12e1da1f9e6f1994a9983fc0be51cfa1519c8aea123ed47ed1a143d977695e8bbfa3079f077b5034b1f7fc8d79f7da7f91dc715d96b45d86cd630b1946da82c3c22d112736da8795851db7040ce9bd326b9b923d31eb3beb84c5182e8361ef1af7106ca2fd2853f485163ebcc7a5bf5755a83b5be5a0cdb3ec41983ff59871b6aa215aeca621c40c64dad6b5b81497a86ddc792def8381dcfb5afcb8ffe371a71f3d941ac4793932739174fbb042c88f2c8296682994668e832c16b73bbb1c187a6b98be74ea0e3b929a6ef469e1a02952282b75e0e8e0a0d38b2ddbe2f6c4f4d47b9d427ab0eb843336c1eeb7aea431f6409fd137fac503a0a5925d17cd6c0a0095bc556ad7961d82bd0fd0ec38af2b0854fa3c24b4b16d9e756f281db2ac1002356dfb0ae6f620208d07315bca488df95fbcb81626b35b7211769d4d907a74a5872a79106c321d9d74c529df63f99f03ebd55058cc71cfab55909cec0dfdbd47811f8c5e97d14ad5e8fc372382180d322a0622688c7a1ce751fbab7c0579bdf1183f8a25e8d8ffaf132669181983628d9a2d59686db47eafd320d6779dedc75bbbd09ab1da4ab197c5b3fa6cf57e09ec11938e0081cf4c427053696583f992692327efbd26c6a750e19abc3f1c3690de753b27b69c221e749c7390a05828f0ce659109cd16e0342baff91bfc42564759b86f914348fff5406a85013d58ac1b45697609f547a85406f280a7034b16465b7d08262487e95c02d8ae29d847be19911213548945112071620acbbf93b7466e2d5cfd171f13ab042679db818ddb0846ba5ee72d81923d35a0b9734bae86747f5f73121129377a02cae69434c8fb4cc72e414402af10a1a2ed25d7cc02bf7c1da8db9e36888d3d8425b5cfcd85128162906cc458600ff65e88765b77f210f5e19164cc618584caeedf78953d8208;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h83ab94ecf036bafc8a94fd45cb9fc6efd43a2fc721cfafc5c77635b3eb2ffe5bd85b4071341597dc61b9e88e83d10be9a572deba91648befccfc5d29d74d01d701668347a0503c1aa16c6484019717adfe2c66e239e6a07ecee240fce492a5299ac9611e259e6698f5bcd4cca189012b6dc7a339bc94d21f54b5e3bed3703210cc319e8d29a26a976a52382d5984d85f01cc04cb918e644cc4eb9d24e59181a4715b49b4a4c5b31638932af5e152c0626bcafcca2149ce6ba3c2808ed7870158e068f0397291b2455ae44112d06350bdd00205954dfb1d02d245545bc0ef8e5db3e29cbc7f4edb649dbc8d1001049b4c1d5c31a0040b9a9ae2d55669238e2ab373daa9541cc8407293de60dce3fd8e45e749bac3f99109fc4e34f3f91478cbaf43ff993f05c3ac33d1614199774bacb67e1ea4bdfd073e53976cc7d9602ed457961e2ad1aae4bb2fc873a285ef2bf4128cd270a5cca5697e7e1fbddb68824291d0f0dcfb684278406961cdbe1cae813c6c11543f6e7b06522149ff59f91b5379165b71def1aed98da6adbf075ab86525428f979672b0a9c63b5357e09990bd760b9ca951ee429491c37f30b264af506592ad035218a3caaf009a6f100f518f13cfb11056a1e9e6ab5e571124cfbbe52d8cb3c15c0d18b7db365d5745755d6cf18a055b80ed77d9ab7ab0b05e7e1171eaa6fa49e1ca23b4fed19165e210ca3f13526fc2eee32b6321f56d247e85491083aeec0dd0b5e30d391076b5085742e9a61db4787575a0e0e3b9c3575161f354da72875cc57d87a8f0548a7ebba5e9a8a5f4a88728ea7396cd176b0a45dacdaf407c720c9198fb827046e4bca971284ada732bd3822540e9c6b5b1ee3a61200005e0ac98de0fba1b639ed7d59984e275d28366c2f0350156ee0ddfe7a2e2d6b7569d9d986206c27817a12852710210f97a3425f4aed377a1aacf5357ce187f0ac4f047a113e6ae709d31dad6aa9ad72bacc884bd43e03840b65676699931e7b6a0fa77ff3d61d0a245d952a2be242b39eb9ebc07da215a6bcfca0b845273f14c693af6d72e02cfc7b6425738b94ebe163dc0226243cd15d3c71ffc345230c9cc2faf6453e6a858022db08806e6ee1bf399e0b9ac316d5c0fa8ae0416460b3edd2f1d06c779be569662d1bbc091261df42ccd622b8f25735e73b41d8cc3997d085da42a32e10414ed94ff677d4acaf5f4bbe5e687f5a18f819eca05dd898cfba16e2a6a47b60838b850364f7d59dae1d100a467c565ed21d29ad8979962a153a2d55408940d4b189793332be971a525e86c3d9840be61803ca9fa9f575fda7f78f0456c6d527c8684b87308b5f57813c73892cd932717e29d3ab016e7861cdb11aa0c1b708c96b725bc4250d4863ae75f79d0dfa490512809a4160f44c8dab2571241a3b3c3fc7c59a5c808d605bcab97d8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he89bb9a91c4c6c76f24c08bf883b76ff7bba6943f91ae66cb644e24add1c99a2262a73289a8fb9ec2eb6932f87526cf1ee76f6fe39d989c9c2c57d4550b37a8c071ae2152d924f57c6e6266e3b4d40de73ff12dcb83d6b13e9dbcfad093c6b7aa884715bac96dc14f6336f4ac7ac270ab8607f55d3075d8333abed1b31fdb0f310b637922a3ee5012b8466b4c4441c0f70b4ce60d94ebcda46749ae52f78278b73339e80971461fbe17735ebaffd1daa13f6dcea566a211516fe94f7a44a05073e3e54b37b52bc2d2dfc5b29c23528102b66c80b998ea4beee64abeee429eebd0e7f6a7709b7ba7e3f6f841ac499464642aa2d1471a5adfcc75e09c1a19e310923859def23788a2e0d3c2746411cab3766441637fe68d8d84434f61124712e0e18a16ae4f68b37d1b8370e2d4dfb1c4c4812569dec0e72a96dd9f03c5b1fb49a73a471524bf132943971e1946993a480e2c4969ac33f69e83e29cfdc94ece63541d434a0e6c023a8d645e86c8d4c05d05fb2cc7a6de3cc96f66c933e5ad96a8084d19b5c3e266215c25a6b0c01581fec87b8f802693fdd6bbb41fc7eb0257b845475684c754c51c5c72baa9c8902f1c448c42d6e2d6a07c3a9c16b3150e23c3fb4a4bab08e52ab2632b02dcdbc8b951434fe22514353d25636c3bbcc3f577c991c90db1f0900016eee01b776f463cd4018dfc8f47557896805dc710347b7d880fb5c5fb8ebb5ec952bedb0c5747e8fbf3039586b05ed819a649f8a04e52b720d1d11dbc445b14f69066644419f0c2fd5fe937c809317fdc5d6c9e1946fd769f89c9c99d6d4227514aa334aeb507bba9962a30d77d5e63eac2f819d5bc8c7cda3a90a87e59acea899d0de228238823e91c077021fd7714b7147a6f8872d621f58fa5631b8ef37656b15046df7038d5a64480d0f69adde01a66938719745c871fe6e26f5467cb62f78b0a29e32f499a2e0382ce4a029a7b9c945e96e1d7b2abbed6ede43ed4632baf9f558e4a30bd91758aa767dfedbecfc77562634cb6ff41c2b57cab137c39204d8b7d5b0fc2ad11716fbadd177634d9705319f5af4989ce1b5d153ee6b8560d31574457b8978995d250ae8635cbbb0699bab4b0b95a262716787ad52b13b385a948550d5e9eb2576e9dd5da5069ed176c0aa788369c5a7274eead3bb6c25a7f8f54bc203810d62ff6b14b35bc1fb3b1d8301f487da9feeade07fcc10f323273abba8423bfe617f708194d2ec250dd38f013aa2596f78f0356b08b80a2a18806d4a3a71106f35182e567648652d657680aa17531b8f14ecbb3a514014493d8779db63e58780a84fed8f00bc00e61fedbdcff4178c2fd82201d0ce99aaa1ae367e9629774dad103287704feff1852a6221213b58cc4bb48710ba22769164e93fd33f64692cdbd83b019f77dfa43f70d4588f3252f3b3c4cec853;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7bd204b0b807593efd120b9ee1ed31e8e90bf399c6cd0fde2a34d68af8a2bbee4e3c73863e8500a768740f96e10c6ce7d29fa868c11598b3197fe80101bfb85f5a293433c222d1ebf5801f97a0f93774959ccb25b71aeffa19b9f9b1bd7c158f3591d3ae6471fed91e0cd6b89b3b4a9deff6ca05205129d1b51ef452fe96edf2b50386e4f457cd217e9c286c70bb4cccee54c36fb246407ba302c25b7d881de20fb58d819e0e782eaa513df60469e4480e201bb7b416f78ebd99f1d3cec13ab9ef0ff45b02006bd26c6e07cdb72631811738344264d14262772d5980ce6b7a690ca124fd8b7625e19b2f76f99fd12eec61ed4ef1231fd78f1167a54b20ff69b0549bc5217cb1bf1574d6f8fde9f17a8d7e4e84b70ed810e1ee4670f1d9a7fa87743eb4a88a8c6603d74b6df5e4b6f591457020d1e94c2c67e964192652f79e4d0b32d0587c959aae035a71049cc869433f319a333f615db09336886bafdd57728b8a44b74bee41f9e148c423f813b5170302fa20be68ac9e8c90a1dafd47d1bdf4d81804ec1c67c8e08f54d99536dba4f34c199837f95e478a5dd9daa0e3a2378abca5cedb23493a168676f2ebf1d859b4069abcfdb8fffe53ea79207a57516b4195624b66542f94b6b01c5b50bba6372bf74ac2185c637ad0ffd5ea952acb5ce16307067f0d875d449696289f01a3c21784a9604038a4c45abae7786f05bd50b308ab9d53ab320b3799a0dd8b445b3f01fd7b79f2639b5ddda5e476243e4995757bf70954c975762e17ec3abc533757bf2619ff9bba0bc5ce8f2c2c514b05f592e21a04387932a2bf75e04abdbbcd975f96ba9a5586c72bff5d239af5efdedb5a435eeb15adf9cb137aebfeb023420b80c429b9bde3f0c07263af046207f9df6d8cb84c2fddec9ee04389e6e7ccd19dc1b0277d55006ae02d7df955493c135a4d293165f0c5759e0f15ff35b3ba88cd96366480b1bded6a37d9246f3879e3acd96af102276864f6fa38a83345a90120946b3ccde4c8f6a34ddced1ec2ad00782f9a7459de756bb0d52260d88a5555d072e7c7cacc1e492798cc9201af3bc14203e50debf015393331a742589bd49a6d2933719de6d6be5ac0fd766763782928346a0704c524adc7bd418f60d7d8fdd9f34bead4c8a2666b63bfd1c395d59df9e14b9a97096d1f581717f4814fee35e26c70d5b6024ffc3f6cbac518e1292293a4278c05832b885d130c245ff4b0d594425adf88424d8b0f16330b9ad385c3959831cccee312b5e957c9a1f308c72abfb902f62d37f1ee85c5de10f064e123cb92d54089c13117ea2a47626f53bd2be8455252f2a9bbeeb61e048fe5f5e16d4ca913e94b4ebb860ed30f891c37d5f1f7f61cc0eebce8ad548063e9283064c227c120c2ef83aec6d5be523eb1fff8415411ffde70365abf169660e70e85e33bcc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he0bb8c8270ba5c14ae66706b5076e0186a8c285d6ce1bfc8903c8a09041e9969423ccd02aee079c4a42fdb45f2f2b15eab2ac2d3acabf86745b8759c483204333a696e4c1f85802bbe501cfb180a31a160665655ca50ecb5a4c3d078d72ca13bbb30a25737968823bb458262ef1d919c8eee34a8716ffe598966c0935140a043d6d8d39692d1dd2168ca30b0d85413e2e6c389a4eb0edb869e2979766fb8d396e69173d6db603295ce6687fa476a54b6b39f94d2706941f2dc85c1ebe3bcf2b88382d8e52b47307eb17b944c7d8577822e108915612d840528033b238d1f6e0697d8c114ccca20b5ace8531c07670d2019d23f6705b41c31706e74af36a971c0509045451d86ce60e55b58c3e7334051265cd859a20b0bf43b4cd69c4527b06f3d7cdb28d97d3f477c830909747e9e4886246a673e42ad3e0286609274caad76938cb1c28a0f05bb7d780bf0c2de20997fc4de419ff699e722e639d7abefaf8b5060281fef3cff2618e5c2e21d18721c3d54af5e39f695ebc50e4d808587e0481a9f922f40411995ac2fcde36882bf3a75b7fe59ec782cfd1508575505f2bf8329460ee3ed0f48643f09532a63cc88d0347f89379f507e63d5e2cffadc7babffc0ba10906491890684bb085673f0291ef0827c989b79662372ab6447c87a22c30ffa676610cae6c66b907a8f83d97802df28f3877701c3b2eb130d4cfca326bc415de9eaf93042468fd698b592dfb53e8a4638712267d30a648ba9b75b6087f98642eee0527f865e676f5c487eeaaefcbdfca5ac07501c5fd9aa21b1ce32ae45d344ed01bd4c01dac6a4ad3ea585084be869c7b780fe525e48c1236dd5264db79b53c12d13422d94654e2d2c90621634c85a50cd2d6c639f6dfed96d968c23d37385918b4f88892b0c742cbaa07e026c8598ce03c2c929f9f10866979ed1e963e8ecdc2af0e1c6192f24ff3e84533dcc2a7397b51ce994e11d976f6a6184bb55c132a6d02471d3ce68aaf4c5bcf8dd2be9d5316fcae4bf6cf737fd67d5e76018885cd71e599dba92e426109eea2677fcf7b719e49143ebcff3aae9491d51ce35857c31a66183ec69c2ce8bfa8e5526e6cad77045697c3398d3f78e60866e597ce26edbd3f0219831e8da7014cad1be1f6f3f3e5c28a10332b019cd3364ceb8ee53218e530d8719023b04ee3655857372ff200d5492f2c45e7b91f9fa8854c4d559074797feada4a28015d634c62c19c6f12b9a56418360d33168f762177e476670b6160338aa90bf622f33fce4419da40872b06f4bd47a60d9cf0b0aa92f2cbbff34488907de6fa05774104b80c8c2dc9934fa023b7400bdb59c027c6634ed606a747127bbb46202dd4995f7c753abcf4f78d63d363cce6ffe653a5eb7bd10a6d1fb8f8901a9fac21df1d3b5c9c64051359298c17d882b9af3cecc8de04929b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha83eb9e8973dfdb5ad4d3314d90786e5fd943cf7ea39883d19295665eb01e0ee31b6fc29cff23a62109bea7d9b546321a5949fd815f8637cbc876266a618f3ac57244094b2aaad75ccac811c619b40bfe02610f35c88c11ac98b4687f69d93441d15bbb250b7b4415eca1ae27c6fae7735f354bf89a36f343fb455b1e6f1b56a66c161c420ca742180548decaac886a1adb899cfac29d50b0b5fb96413c8817eba7d50ac63c999fbd66fb6d798983deb82d413966df286e000bc9907f65a0538403d5743ec57b1951b3d6b51a67fb7d930d58496a9aba6a380c244f761df59476a7f167efc2efd52f55586590d7ca1531afa41369b33b12367c883e699ec3f0e5bf4f37de8f0ea91c8162c61f0c28f3da9c3ec09484147254857e7a46d6a989512f36c7ce3aca863ddab28d2d2e394d8dd1c3c259d645e760d8334456c1e151b36c982186c358ec0e8e318a1aca1f6b44b79bf9c9965d85ad856eccc93f0c48de83d7d3b22c7ebcebb4963b9fce3eed0146a08965cd8a404687724191d948cc5060fc42adbd9937c4d69023317d7c0a524fee9f82b24dba3f393f1f682d93a3bb59492d3b6490392438008ef29015046b2152c66f414f56543ae85257ae7cac7321f041fe0a709df5a82071d12bb4274824232c74d3e299dc0c6ef3545d6cd262f82ccb3eb2dc8f3fa934edcbe273b41759f4fc9c3b718a2c33f28c7f89e90712d865c39a433efcf1471042f30e6c5423843c1a314f049e4e1f29b0e897f28490cf0fc4398372ac6dd979627b2952c303f928d0363556a10ee94f3404d96f548e0a24501ae82216d007aba742dc69aa9d54892fe20deb62ca11d79aa35947b43447d6a7db6dff707ea8bf125096fe5962938f43bca542046e8d04ae362abe171e6e640e3e9f03e9f65e4a27824c875da54701b099cd8ef1c72c118fcad190d4fc0554ea40fdee4fd1fc3803b6262d5616d1059dca45d732018c18eb9838f64e2a9154f70e4ce47ca96ae9fbb20367a898196b7a2125b774a729b75fc9d1674691caf61d8b958e6c8a94d38ba00b506a8c0b1eb724b435568e0c76a9fe827ecc5f18073458d495139691d93e251c1b86909112025312cb8c638d122f7c580cdaf1ac8c1723772fc3a19ee4805490d674725a4bd436db9e28a405889e6bfa9f2cb02141dae096df397f355012428bf5abc0b485252b0ad6c68c266dd2d33c2874ea3ce46f89793055896ca1a42ae0cd88d437149dc2f24ec460aa6873cd5cc596deb2a79b177d1b6f0a84a2a42c9e5c8d4b2bcee05c2645512fd67ad0404ffd94dbe50180964927593e1b389e649578dc680de6507c8f46868ae2f9d13ab2ff62467bb1a91f6daa61c4e70b1031a98239799068b602d6787db2631e26c8e7c545267f72cfb5835f45cb188d7acde052904a1e74573ef001492e71bd944a2f4a00f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc74801d58a6d3776babce2a710f369b6703a3689d84d87b0afa7b1141fc6d1b0b061b8dc69adc7152169a2402af2f9207fcd3c9a1b5237b9a897af1440bd13a200fc16ee30ce2e668a3f6c9167bc1f36e5ba612fd73f06d67db5d22d71f3efb9f7946cd977e73225547492304d346b499e887cea7d97afba5b6e85b66941373ced4bcff90f758087ebc50fc49b0328b40ac309ebb01b43c5c9ccf3be1af2f706e8f8b53f410d257d42531b6713e81b4e7bbfa8aba65bfbdf926f30d7224eae533b46e4a05d548fdccef358b533e61063feee7088018ff034345a883b8b5bb50832cb2a280ceeabc13fbb1a5275d3dc11695ce613f5dc208ffbc093223b6f82a1a1937b0afe040ad2de6f4daaa2b230596bd766d0c1cb12401fbf09458a26c4d16e8db7c13bfbb3b6dca465212519e23bf52144c7bfcd2651c00c99ad3fede112140eb7e8b60eafe84adff69627610e56d1c6131609ce499944dd4174973378422404a90a52c68660a2087d4d100824be4c0e67bff56509b422d859d3e7b8ef66b5f727115fa99e677ec08f8785702cfdd1c743da176c519a17c2a7097c503701ca6866ec59b4cc3c9f478685f236c52584f218c13ec107944279d776e393111030b559f1c0eee0beaabf8c71e1025292741bcd6b53a14b4ba0d29fac2a571db976ba38881970fb9f99c87e09a6be722707c7128e95ab3aa6d660a8a618b36c449251a80ed4f8c21f251407a5e88b44d506ad515e3acc80e29e1997e966402f76a0c6c1a1156d7c73ccb8666efc566b6af1719cc72816d09427017049dd4dc488ee17185f0cdb92e6832424939a1f018a5f8ab824988f861d76c75c70afd6172fe868af9bccfef01a8925caa58bc154397992a2c571f8c49d54e0ed28122e16f42b6b086bb83a2a4dd04ee0c0141d8978f06e767f0106bf8a9e08447e389be316e49a22b39eecd3af961de28718d14d6e863e90310ccd243d4100e826a4df9000ac03e0aac342c3e03049ed7dfbbe06620d0110e423ae446007e7425cb1ee728c5d75c01ec4aa675952099132fef33872f05fd359e9c8333c54e594c49ebb3b1b3c4a617ff4e0d9e84fa1dba434bddb108f40f5ac5b14db1f2087db9c3ca9c97804b07b616c6df2eea0e5f9218114046e1b8b42a2ffcf3a29d3565976e8aaf04f09dfb035ef71fa3567f5d51994b34284d4f0f40609e051f19d5f279dd7e666847a28805a7260cf00686b9b196d9d3af800f47dacd51518b972d724f35a062fd3f5a518d9aeb04abe565269b5dedccfbd787a7227c28645ce2a0c88cc8654c713e1af59438d60b4c36c18e38284dc9b7d8eebc283b49138f85fa0d459ffa5bb1e57da7f51d155f12a347a88f8ebb2a0477b07286132e9d361107f648243c9af531a64e15a568abf27a4ca9fa02ba6fe00d5f333644f6bdafecd6152e71f373c5a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h844a186b3d0c74beee04af0edbd71343a37d43e268f1490cb41d1d4bb9c6a4ea3fe3093a9a4a152f6ba496979546419904377cffe67e2c859d35177832a8e279b20d6c433cab8eaed5d570b2d441d65e119dc00a44077a17aef844beb42ce7efef6cf141a0930e9df60c72b3a59c16b2f770a06136303620a74d9f444095105bd88c2f3fe52d4ca20e5f1235b94e4f756b862f3670fedd7b008a993c67a11b4a7c8dbb97f6f0ae18ff199334c87b380ffd2adb818964ba248edd913d5e78a4ad134386b2dcabc2e9b6331e2228e0b8ea0bdc5382b4ff60873161db4934f1d7dd37be5f43713a441874d4601b65559437b7fb32b07753f30a048e416dd668107db07f8ec99ffa70734ed52c3579d200d5ff9c771e935d4a088e8cef729c6310a954ecf70d15e3ecff99e185e3ad66c2ffc843919ed4f22e82ce6e4702a6ea71a6c2094080fd722c9fd9df629ca395e8966531dd253523f5f8eec6c39f61c8856efb4711f9b5558a0ccac6b039a5ac4e0da4cd4e9e4a9f383db37ea3e40034785db508877df05a275787e39f7bca0453923be2210fe9691f7c67bdd06f1577d6d9c8f258232fa7c6fc216ddc6fa455b0c0e2095d3df9216be6905555cfaf20cd0de15e93b5a5ec1a5d82e4b901c830d698978e5075acd53cef9d38157164f591ec1845d6852750a262ced3cdd674005351a56f5bf39bb11c685cbca5493dce6eeb9ecbf7e02a5f636849974a9267bc019cb9e1b1ec1c9b895dfaa1b9d4dc9674d291aa1bde716ab733a6017fa9ad5c8567312007ef2c1d1a25245fbd05d65d67d63471b4669c5acc9e4ffdda7c1224aa52b63369a259303df535b79744b983d6a975a6296c10af6e9806bbea870d4a8908fef0d7fbfd5cb90d308192d946e369e639d30d3f0bc0994f1662801ed55b2c597aaf6bebdb1dc76926053acf42c8098f288fa4cc73147db761a46c928a8f1dc8d5512d31d33ddb79920d4695d4d10e91baa3bf74e90c0753c1f032eff490fa6be7dc1fbd1f5fc434b84eb1ca96102a22cc18bc199969b4dc5396982e6d75e8e9372cf9536a44e69be9c43a7ef924098226d601bf62334d62dd923a908be2ddbe5f7cd6f2177282895e7c4daba1a256c550dfddbe041b08d481772d1af0978c4800208647ad090fec8b76aef995b935750418145ba5dabdd6eb453fe2251256a115532c08f5180b9a751c4f10c8e9d376feed4351bafe2f4c479f05b5730203ba41872dda6bbff00a55e99374bf0785a88f5f4634cfecf53c39e12ddfcc2987612538e9472e7a76eb11372b5c2c0cdc75d7ec556d437a217b62fd961bcdd607efa7b7259cf499a687c6da0e6dbfdd7c245c43c7beefc84603cb962849406bae3ce5f4bbe6f58900d861a8cca095c9f2cf8cb7774ba5dd3185be47504f54ab79911279169941557d96f1e6c62dd6d45c9c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9d7c2b0075dc6950557c68b307712525ac319fd90f318d90c118012f46a24a89ad3235980b268c619e6577cf5ef6917f021bf5f7ea11d1c7548db7c6faf57537b0bd5f5e5a321f12f8e678f7970b2d99cb7e043a45c9f415860e7a911327605c097857fb94a6b5c069e0c282da8d67057397d46824663098fcaac43f06632deee343859d4c4a672551d9e23587a827071f44821630e90a8a8c81f41d8d3047fbc2a05817d465fb9b2515ff7c5bc0dca6974c00031df3fa9ff44beb0e8bde63e9c1e132dda7162ea99cce38431c4792491dfbfb535e8a6d68df890083edfe24d1a7499500db609f0dd842cb8631701fc3d1b5f122199f082460f0d6e40deda57e189b6bebb63c5824aaba973c417ab1e69f6e3492078957b614f074327508391eca9b7883f6aa43e8840164f6f810cfa325fc4911637184f8cd81b1a37386975e2cefb0c52955e76dc8eceb5393e709dd43f5ab807853976581e6c8c8a7e3578713230abcb1f508eb5868fe5f96c12ee1fe4259c70897103aadfe40bc3f3ee386c223503313bf79413a873d685f9f04f85618fb9dfa1776650f78f58a4208b6f8f6c590ce0ebaa5f2ad0ab751168a2ecbc4901032fc9587c53cf42e21e6267993639a1aefe5213b0a4ea6d871da67069a9e7f9e86543418b61b257a094341abd210309842f324d65af9076f21f4d975b0c31fc1a5d94967f28a9506dd281ad855dfea9877fe8a465fc891c1d04359d82c0804456ef2421a361f0b4cce6a9b40d6bd45fd707d90ab781de94d04b54f25bfe83221d1852570288424a400f77eaebe9f96ce81738a91f659a519caa7a233ff1b0d81720623545a4366e043596d16bcaccb07c5c6484ff46b7e41221b89303d1228b2d7ce867f1a2c8ab6d2dae9929fc198cbb4f34a48a0c607478c3ddbcad9b29d7db4f26d51fcbbbf16209470dbff65d1df2bb0fa66dcf4070fd98523055977f41a1162f53f76970554f975e06841a2264a15405cb9c5f3dab0e02a7e1ba7d7765220d677716990ca37571a65c716d37529d644f98b30512bae875de8922b23fcb3bfae080353f854c495d5856e11d861c3eb08c36f85058199894f29b660cae38c4c3ecb3fd9b791099c4d82bc02361fd77409b09fb98e878d593aee6ddc36e6d4d2acdc055a29ad501cdfaf8319934a9f86486178bffb9b99a0981cae7ffda352e7281365f08073e14a26bb0ee9f2cc119fb0b647f1cd143234b8540529492a7ee6df8084484be5e36189248c0df47ce813b78e66bfdc47ead98c0be59485577d06d7c78afff421caaf3a99e2306b31253d826d6c8a3dca25dc9b2bdc3b1b4f57cb4d9407de6f355c81c87949a2fc173aad8a9177ab26ef8de3e22719102320d0fa7017ea3680b51e3ca21f8cf4ef67695eeada69635b0ccebfec756bd28d34a3cf34e3d92869d036a4f4a61f1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc6d3138201cbaf7995dadcbef9bbd1a9eb5b082d6f3fcbc4ca80127b9e3100db3d8aa66b2be9a6533b1cccba6614654865fc2f7511fa14e51cb95573fea6848bcdaff09b3a4094a9b83fe874ea8b7eeb82f887b4de836fa84162db0677ef6c0b29626b127d4554092cbe8940de137baf829cc52d1792614ef90eedcc646b4ed8682d63167d1caa0a54613d2fed755ffcf7194d42a33283ec9a3297da24f36437781689d02d4b69c4afccc8eb692e4592c0e7243f6d5324875fc197fa7641278bee1fd1ed3ff4ee865803516d79851a33ea408a7a2ad4700b904520bc6f6472a6f503e44a813aa9eef056a93d16cbb04912a99e3aa6b8f7552f0332e45fc3bf5f9cf17addbd3b67d0c69554e5f53ea00681d072e8344a27dcd66603e6bae3330a98a50ed8d6c36254e648589ffded37fea5eaca8d94b0651783ab6f7f1948037f2a4a58546de1b11f5e4ee02b957072786b2a5e4dbfe7a77b28ef8c0507ffe765d4238e1bf5263d7669781f22f02c1bec5ed5e27effc865d87707db21a988c95c6327a02452c906057789f78944f181257f7df29f8f237a264f50ce5965361e60495505dffcefd2e3858deac0342550ac593afaf4a692d60cda5b37262081330f3d7bce39c874fcbbdd49860b3f5b892626b2add8fc7bb3222c72250b58a00cfe1488e34b6f392180b520727310510e8934072622dfa67383aa8d42a485be2d0abf15a70c6654a0b838dcb6b38a4b6babda63bbdf6c9918108600f4290ee664d62b8dd0365eee89c31e7d29e644a000b402ae63316f620ae31cedd6e3b496e16c8d91c5e293c09de19b2b1ab703c853176050721f17eedf6f45af00136498ced94625a52b3111ab2bf54a980244e6d75e0b6eb7e8ccf18b9c8ced5115744c6937f00e4958322f806fa15d74f61d840c945c9cb2e28dbb09ba46f3dba6b9b03509ee6d7234295e02e44130ca05560569fa75e01432675435be0a8fde4e6c11b1c338ea070fc3d11386868bdc9004a30f3bcfd483ac9d6b03871d717ad52a170b1d28fa557a8e51167d529a008e6d553a8dffdff5aa9adbf6625ce6a20709c35d7657b4331eb35473dda7da611036ae9e9ed35f1c6e11156de754c2de2a4981f9f155462ac9b251062c7126fe3fbad8afe697e5bbaf9cf8dac2ddd1b70c685ca66de05b4c25307d0d7333bb63125164d89b5bad8b1d6d0bf3a81c3ee8645969ac979c21339fc2a3904a45488384ecf376182da1728d6c942cfa70b524567b0727411970c55b4c1cb3f5f3ec3e5de6bf3e2546b7e44e8e5577976238437d018183b0bbf56fa46387f95d22e303135558409f2c7c3fb4bd28e12c5835d20e0b59734b881f2f65b284012e43dd83317ca5b3f0d57e95f136dfa133939a38acf235f8e7a757a5c80519254aefadc494e60c10ae521b59432316ff5c3a7611ed3f533b91;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h94b1e5c8e9c021beeae62825b8b7e8b1bb1f5acfbbd5ef201d350efcd7611958d7603cfe9279090e867444d5ba046833c47c079ceea0d537a92a1ab1b91ab6656004157afff3839661237b2191c2180d759f856c9f244be82c7629e2b0b5248a4ac801b051f96871ae7d428e3084fe390e22bd98379135b1826b264c4a06ea1fd3e8ffeb30d6cf970f6f630d365e47cbbc9dc9988ecaa3a06871a4e11b02dc0c41ad2d36d0726237dedb4733c8e14299e1ad1ff7a944fd3bb8514fef52bd7647473b9439f5c129279ebe79883acf0f0533bf40dde88e64b00a6a32d475d3ceb98c9653930e034d4add78a89fdabe1002f9117cd4c9584dde689364a8e3b474827533e5fb98932cab71a9fb982f638a4480b7b99f154f41326bf17068e8bd76434b333a5b70fa799a61ee5d10cf4886eccb996844e43b1a04f483e063818f43f5e45db825b700bef7a1b6fec08e4412d70279700e19419cb20b296b0c8eb9af777b1e40ade688aaea77476227cdc9b210b5365b4485b9826ea433d6b68f76694be601c96f4f487080819d26ac3018b45fb99a2499f7a02e77d735ca07ce5bafc6f15c90eab2d9271c456991f1aebd8750b5c9cc4876d18d84b15451cba84696b1022cdabf7523b47b6aaa195d67e071b9da95390325cc9f33c3db3327ce8caa5553f02bdc2903543b28089d643ae09987039e5de202ae441c567c240d5b6edcb5783cd4d98dad1687e9239863339d980e7ba43923f6c1f079002dbc990bd813c6cd92d5b26b4dce929b3dd30156c28f2bc2eaa9e4436e27956c1c75f4b4a7c42a2c1be366bcca0ac73d1087ff5fc848ec050a4f75747b4152da723f585a6ed81a8cc3ca1a74c9568e31a3283453d25b845a95a053516c507d7fd79be12dd11a2a52cfafd5fd6ddc49fc89349366f50df9d527e6fe5b702f9bf86fe5cfbb3a78cee9d73a04baca27a3605a0c05e8811272e7b522bff3f217e6a93225e086a24463296576f264ba74d7ab38e7b6ea1c1f95727937e503ee6c6d723aa715fc155defe3ac21cad6d9666f457124863c38587069aa7028d682575bab6bf4dd25598e85fde9fe72148198c10d555bccc0708a9fdbc46cdf64b1040355e5abc1e2a7901cecd51c0ad743072e2a884be55b40901a1cdee192798922261ec2d4fc0127cfb31bc080db748809ecbdde715483e098806844b867832177054d99b94b6d1dd132454abebc7ee063ca92dc2117f41d313741b1df75a55219caa4476624ebe843ec7b308de1208920dc62fee34d6b72cdece259cf8012f5e2768ee37c5737f1e26ee24555a8cc0cc5cac095539f7bf2dcc4e500f352775b4075dff7ef7209346d200276ad5f2325b83c0dc366029107138fb4f60494ab6776c2e9dd0767c51949d2b5c6e95bb54a12385ee87d37dac1e9a937e953618bcf019591c2fb0bbcf3c210;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc4a2cde04f60da16f10d720fa0fed20e5394b41f11bf8f0217a80227e8bd295e41970c9e49e4a309a1e63ee583b51e70f344a44670e25ac183b6c29aa1efc4db8a01426f896b82244999e9b514c1c090dfbf7afb9e33bbdba335249ae83ee9def0388dde96bc47936b9c6b2fb9833e4e3230736d8f173e32940f3c703b8a20ba6d01a3f9f613c60c2c010790fed0a3b6f19b9bb1ffba1ae5dc8dd8b770572cc366c9f3f74ca25b6b7e7d9198b0987735350c3f94a5d412a4f951836ecdd459dbde0b9bc61b6dbd7838417f9e8d73e5c427e6ea4ec9533a5232010a8716c0f091f3b05338ed9bc0a0de8439fb0f1ee0dc3d8976ff58c543df2711005d897eab6eec783f457b47a597c62d36b720d38d530a0a85e4c6e5f585eec557e49122032424ffb5d80a6304feb41f9d67e1cf0eac39020097926421b14933aa28595569c3d55c04181eb61a8f73c18e9afec3e92a217a314df0a5ac45a2c68803cffe4ec33540b39b9dc9dafb97c78adc023b5cdf0203c16a784c9fe4b34fd00a95cd4db655adcec898044192b2338f529c4dd74871a7a284aa3b96f7ab5f66badf271296f2970773fc9f45296ffed16aad858c7bd3b5668f216a8ee3463f85bf7e464c8e7fb916a8713d4b453e16c382678c81d1ce2be435d15b5a0c2351f97725f4d8cb7cc025ee63c75023daf29630f7f7d3c09f1270a299b794ee1e8bf3424b69483f3fb01d7ba46cd8e6d83213c1c0b4b2bd3b54fb01636772e418e1f961b23542bd9f75b65dbcd254a55f91c2edfd18f13f0a3084cf8a7994d860bda41cd141e2c458c7997fc3460f1794fe524a866cb24ed091d13f392219ea359634dc6609c3a6d2c997624fe6410fbac41d2b1c55ef48295b6013bb25c7e287d5dcb71daa168dd9a3def7833e3241a7020b8698d8463ea98907fe43d55141235f316549fb94427ca1ece060db3956694a595fbb43986ffea2ec35678a79f6628c152c709540cc2234e92cc1c9a2e4cbd1a8fa9448f69ec756c069694cfeae652cbf9c2ec97c30f5234ea503a4083b9002c47e90b5cd8fc107b7072cad81e1007e6d80730d547ed8e45b23813f2d1041a5b7255f7c32bc6600f5bc1d1c7e7ae1e5649e1d99e109b691b102f3a7cde00a8113b54078e0d44928fbb76d74ab5f708a3e484953bffdfe8c39c8a1646147212c8506bfffb4cc730c67df1a1cc73c6574236f2db0101672c1cd9f829505860b449b6f10cd401f3af173ae3573eab7e1b9cd312949c2903464ec64126fc8abf633c52c9779c847943a62c61723e89d0f404cb2c4fb299dda0fe1d55fcdc1173384f1c370ce8ea1fa328f1dbaf7095a97474cdcb903252a4a87466b6dbbdf4694ab86488ca36c5c0929de7de9ddbd13a098bd6d15cf7ed89fc5973ae4fbe75d1b03633df7423aa40cf49bc864e3f921e718ba4a4eb6b62c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h486c8c51369fede23221fb2738015ddd918b6712cdf054c2f0111452ca68be6a7d2455d726bac4ae0d9829db539acab297d4b6a0dd7d95be2b34226333a04c7a0ca39c78318d0cee880c84cc23e87a2d9f221de65395f65a1ee29bb0d2586f0246f95db8369c8c25e3b61af5b7f1feed0ae04f2cf795ad2df937034432315073043bdda5a5546cb87b8b2398d3f93fdee660d567869889c5d7b16169258a968f6be4a2ac9b0caa5a700e374788a317ae0fd2dc0a3586615bcce950b117cdc9e315752cfc7083b382798cfd7421fe0f97c71e9f336da0e2f360973c428f869e738c62a6f0a111734a0cd7ae126af3cb1a4bbb3aa9f3b0274df6ff5b0b5729db6f3abd8da1e01b2337585a016241e1d80dfac9c499bcab599b57c0da459538ccea00500675a91423f49b11a2dca9729e6000c3590371f13cc8c5eb9e89ba055664c36b3928dc4ef9a4525fb05a882370062b0457dd3e5cdfb6dd249ab8d6ffb362f327dce107721c6ae957821ea59356aae8e2adffe06017df18b80a12d7f66d37c3de91c63dd37b8e1ac020d548da45cf5ba89be7fc95650e0dea3eca1e0c18aed0fa5acdc13dcce1e384c4bc07cf8df913ccfe326d154a2ab7d090c729dd3cb273223dfb34395a92311e909c318b2540f52172fda6a392716cb7a82746fb52342d747075e0e129d1fda4646d2f5262843a80ddb96b9a4d3b87ab36d7d00228b4dc24dfc88ee378b068634b85057308ecb6bfaa431c5482cd4b11ff807443ca1d88d5cbd855ae51162d060ab9fd0eab6d175bf045ce2981ed92253637cc68cbec879a68c895b33ac19b10874e5a89dc880e244e56213d659c89ae7cdb8f51fee703ef8e0f8170b17527b6ef545b457027138026f6301e244577097c31c7f203e94989718087d44ddd8f0fd1647c60361ade4446245acc04dde52b6107b17828de6954990ef00b55f27a9224550d7751595b518e63551c5ecb62e73f55895b6e302ed39a574f588bcc39daa954d8f0c3847193235c424cfcb8d4d5b0335091b668637a0882dfc3d305402149dbd7707a1f2c8c97ad85c0904323d876793c21b3a8a50220b57261c41e9aa61aa8f9ed1ea16d775121df947a705873a8c64d3091ddd9d1a8f68030df0b3175a443d31f72bdea37c6f6afa34a4d9b694113ea36b6065542d85ec8069c7012cbd18e0a0c9dce83cab650120ff07d695be33398d3c51f94fdba8bad46351936351145c061b1b1aecafb6536fc40610e200b2686b5dba87f6650ea99fab900575f8db8ab890c9388bb78b0a7cb4934e3c28c5811e61717cead9b3761f3bdf992c745d72d16051dda296dee74f4a03bf6ae48c3a75450d14c9984ab73a4ffc65df57f07a9f2203b324d7104060aad3b194532c4f9584e81862316e88a34cd125d27a8fce5ddea6b9b7875bb7271cc0ec7ff413ca1bd6973;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc545da58c901f1d80dc0dd569a6d5eefe53ff6f8cb55e3c44fba801dfe20e041f521e21c40fd17b9e20159939cb251060bfbd56acaf257cc25fb7ec87cf56085108cc2fcbc140b8721b0530a2cb21f25e175ce4afe87a7076a1f060633eb174c0257de312c704bcb08d7c5d7c33ff6ea558a9fd0d2429a71483d2e665626b6ca7787948994b6c9edbe1b61418b3eea4af29b3c4f979d737e31fc93fe7659d93f7ba4bead8b8983d47f5e2b45a73d30b5888d047d407529dfa62abef573edcbc8defda2549b2b3bf788e34f2edafd0d8b8aa95b008664e7a54a882f8d32a0ed47fdf91a2f3b1a2794783e4ba6409d6947a8ea558d102d6a49b2fc219f7473831bbaf094b4f201a91079de91e239e70302956855ae67fcef5a71ba2b611eda07b141eab2b1fb0eb34f3a4e54fa94e5517d2697c9a2793d32b4ff7c41ad0dd6acc24d7db530428e38894497ed9d31879fd1749e45a22305b7ea30f0de3c57b44fcf570509484862d32606e76d9427e94a580378fea3c808d89527322f0c47d70441c3a0b89ed140bab42dc507cc353678b7ff2a406f3094dabd778f09af262cb0ec6ebd281642e3f77ad6e26ab2c94803da740e79945ae2cc32bca6ccb02f2fd0cdb6dbe4ba0539931926c1f9d2d96a602395d68c18848c6ec49f789be007d818e467962dfa6d296b50e31f26d53122deb1aaec01fe3342c2d2be685e7bde84c77085a3301a6753c9e9e19cee5e4129471bcb66885b834f9b5637847bb124acf2af8495c6019775887ae3455a3eb9ed19985f500ce1c3c5c42de8aaa41105411b954ff0ec80d3a6ab886853fe9d6c70a4a63e9007716c0e2a4686dfaa425250773f90f3f158a618eb0bf2f78c796942442565391b247f3a780592a55d14377e850b66cdad662a46b87dbce6d0fa4cff2cf22380ca8bf6ae9233c2fad94a18b0d39cd42e3fdfb73df30b2d81bb816007f5624d49c13285b6348e8773889d852ed6ce92451e2d652b1787857356055b8d0939b43db2592d8e5d33cf4508e5d1389d7af0a9797f1a37f993b4fee58e581c29e4959c9b427b4810b4d1147668d9af0545cd8f8913c1e25cabb6d3dd2739f96c8d4620084c3cd482663e335e7d12f8d6ffc6a3c01d7d93df6e6d26d96a7d63db5a72bae39c7439f83c50cef0fe846e15e316edf0ae4c8d4cf7efd79f0b1c78f2ac89f15f3e06ae461f588ff075ce842fda40577d1f7a26102811b943ae77797323866eb3d6f3d656f029bfce1f2036098450ba692ab73b4023f6ec11c4f511d27313002048a690a8e935bfdc0b6699cd967283425504229ba35b18f6dc2c6188a9dc4ea990b6948df3a7122a7aa83cf866b8a4f29255c4026f2a0eadbe0ef4bbcc60cb0f27de064fbdf8259b69c09e2bb40594a10433872df1aeba5fa7e261d0d0025c32ab955f6873704e77801b474654;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h828fd93984e5c408c43b78cfd73fa5c72b44c9dd878a739939fc6add4d99714553fa67ead4f0218bc7923e941abbcc250f5af5b639dc90449d503631c166ed8613601bc04d695ac74e5fac875e3130e037b3194d9cd96dc86fb539d3bc5ea00cf1da1edea8261b69f73c9b471252d3fd6bf2d0b40569021fd02191b198e0ad9371b1539f30c386c92c722221dc843de14307d267fd198cc220716192d90d931a874a921219d19069427592c8265fc3bf7c4df552be483fbde2269412d56b0685ddd33f03d6ae1a212aa14837dd1eb174d3f26a370c30122b9444503777528c732cb04829b8e80628599563a5930cec3af7f09cc280b72d883ac3b2face0a0274d1bd82567a35848bbaae24c6f8767e0a5f57c3a93c6661426fe71a2eadf9ce8bd48b3b9012da14623a4103144821b2b69e5963adaf5fb8502a66cc93adfe0e9f89565e633fa36250909dba2ce9c9b486de96397499826193ff0a5dc25f2e28f03bc6c53b135a0f1a15dc94cd2829d0ff6252d2cb25866de08c1e80c2ef2b2d9d92d38e95da6a70109018abbbaa25b79352e2abb58d338ba7f2e7da20d87819b2704bdddac7df80b2c66b9dc9a80affcae8e8a8c19a960dac686172e6f7b62689bd26a36c859746159c8e588b4e3859b53aa2e6c3b5928e12ef2fd254b726ef65d32534f2c6178b548e67fa1e4937b19e327915fd0506a78ca4991b5fdfe8eb5c32bb553a90d2ca30cf7e443a6a24aaeb689edf8326c5eaa79bb165b2c8c16f3ea9d2af2ee4d1158bbf21122b02553aea5e4ace1d38ecc21dd7bbd0b4bfa51636c391d795368948f37b2f5913bb0cc2bae6a8a3a38a5d7349c0821086264354e2b20f082e5f9abfd360074187c080fd9099841f5e2aed3338ebfb31917b85522e604478e93bf8d4112ba7640d342ca93418c15cd38b0f9767e4b6ccafa02e00548c716d7af38985361f8ba85bd22bb4883b8bbc2887bd870f0a27c3484657faf6e370edc63477d13aeef97242d5621cf1b2372a705475d3672730f1c8bb8544747b2170fc604228abf15a6d04f9e43c5f4dcf5e36d2d0a94add883cda748a4a6945eb6ac84724d854976d7d50b7dec6316adfcf5d9d2d5a7fee8e89404ed75adf1873ee59799808587b7926a11ddad0ce1fbc1ae0870b4765c14e87fcb2f6a56777a8c36097c206565b77536b5ebc0377bdfb89d9c948f3e27ad9843fe1f423f47aa70439b6f368ff1a995c16d1f5c80bf3f124179fb67bd0e8fa738c3570fab91547359979fe816bec982a1207a360fe702accb7d9c006fb2ee13e365932fce2aa0d4d0018cd75edca56a809c358e8b8072346e037384ab7db3216c1269a434b7402ddf34a5576cc589c7a53cb334a555af2ead8e409ea3ab224dfdc87b7f01286a4f9424fba3b716da03cfb18f6b817a2f836f64d61a9126f217633ca0b67d9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3f075f0ae1494d2e6d5051f4fa3f4ce2856b0fe0b358b0195919eec2952f61b1f5e97acd1eda68f52edc5d5f3ba6678d24a9c4037e8aa34f8c1fc2f0a66d6346df983edc2ad6831555d207782d3b26046e5965f3f432d8accf4ed4be4daaecfd8956dae5595207f6ded7a8a1f55099dbef54f2711f25e6e63b20ff263e1b4bae84e6a91d86fc1f4a1f2060659960218c6a5e23e759f58da06f73dbd49b233d65d58f2fa1b6bda1c714b8168cfb7b48bfad4c003a6145700295fc91616f6bd37e4ba16fb95ea100daf24800ee2ae93fc8f34b92eedb3d7d45670f63f117225244764ffd92b681afb324e5db95a82fd74b4a7b02ed1b2ac56bcc174e50bbf78caf78d3278c8f6048c4a01047b12800ea10ea6a6ac8b7e8d8768da1ba6ea2c58c20e64b266c2cfcada88367fcb88e6236b9aa9b273e1210723eb1c38e30294a860873fa8d81a230aedf70a41b3b138bc53aede92dd15259b74bc3efb8b47cfaf1aa92527f04f42cb42947a4ff1563624ece58279b0f7edbba9341e446b154a4e87cac54f7986b66069ffcd49c0ff94946314f2f6e3099cf35d95827d97098af6a652bf845dda3409a9964bf17f4adc992fc6562f2277112af2e684a14d6f363f9b988b27df445ce994633a1514ec301bb7e011a8d9e326d3ccd8c5cb6f86938448f282c5f73cbb07ffabcc55aafe375c7ed95b9673101792f3a550c51fecb2e78a5f00b4c1d5b19723bd79144a6f7736b52cfa702fd14c7a7c08ea55b76f6d331092f4642d7f01b5b4b773fc0dc4fbfefd4c6fc6715145b5923b2510451300915d28115e4ab84432d6d60c051567cc3aa35a30bf9e4a3d80a690b642858b363926e0b09ef9cdb91c752d680700aa9b668659a94bf098ef18de4368484ec353ed45bc0ed62c515e1fc48286335e1906e3c2dfaa021bf12486cfbace0a934f8fc051c2fed397e9c5e5dd017882983e71f6a8388cf8628d7ffa62bc32530cf8286440863c0f8e55a7b62001a43c143a29ab7c6e7c72c4689a01341c6e405c620900fc00e2c18a897a40e265702fe3be4e294dd7007f8d102cd5df901f7a363fbfd0742ba4e2a28cf3be2b9cbe9efad39506181f17b53bcd24f8c863dfa59aa2f841f0b0bd57c3ebbb01bbf094f9b8f9b4b1bac0cf171ac08b4e21b9df99f998bccbf147732a3bb5b1762d9b436ebd4328ed3aa0628d180c061215a341446ebff030732fc35fd8af9c8e9a225ceadc0b64bee4842abe5e7a9e6e2aedd180fbb0d89bc0af5867d7e6b18d9e5537e31e37096aedd8416e0498c5a68775b6277468587cb9fb1afef2212268a5ff6b9e9cc614a7fa4779fd3c09ad73e785c7b5e43056e6e26073ca9d4d70a246c445619fc91e142dacf13d477cd8af842d6a9ad4301bda71b420d463b3244abac4bfb2e2aed352fa678085cea4c95db698ec79f67462fac8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he00baf389dd6123290062217c9b6691a83cabdd1edca59c45b577d5578d59c76264208a8e1ba4ddba457a7b101b180adc95903e5eb5649fa9a3537636d82485a325c805f0982fef05875f89b230617b8d4785cc1453054028ae1a97bf175b483f4d8b74160ef67e59388545bd5a1e038ddbd8a4ad6ded18807bf1fb436f76c0b66d67f541f4e4b39baaaf34d259745141e36f1f0237b067bf8535b0dbb7cfac4643280b92ee40dc7bea7f08a04a1e2c2717a4cd03e3c9ea46ce5fbe82fefaa7053995e67603bd1fe02fd8dd3410581ef405a053b18375680cd329c50e722c7de652ee687c78e0c5a4d0da98a295637cb0951cedc62a0dbe1fdfcb26c3e270f88e00354be4396f6e89d0c04710f69d56b48ca71bac9c6cdac2827efd296aca292a9834b47fa1988b2c588df985ea340fa7b5905b8b2cc4f05d9b5fc0dc66ae6edf15f9d20465d623ae3c47e66a5dfedc614fb372742a19a2825a77a667a2105745d0155f7e906f565ac93a0144054932e849954eb6306b344ac238d8cdbee4ae5130bff30163fb25834e87094f3bdd4852638dcf44dab4689c025a2938b5d6d625a0c1a181582aff5703bb92e5b1b554ec8210b5ead498069d95c4e16b6c87603d689b75bdebe3473d272aafed4947b688ff232b7790d4684c7883e76722d890b543cb644e47634d8431431453cd8b9f9f5498e30408499e49058e9e7f1be8874dea74a80425c2681f7326f89febb321910af7edb43939880fff233793413be54a74bb4cb673f8594f012342f5a0600b35094cf3152e10780558c2d0573d14952ec2bf887d830bfea6867e28f4c58264b674fbb5604f3117f5aed21ec8da3978c763c6f94b7ac4b1ab1eb672796d896941c66b524bf330616d6c338b3723ffdd175aa10e52e9a7869bdf71a6f512f76f8b63b0fa1e94f4c3d0709e4176545e9baaf143385276699177f6df5a1619cf05af4381944786503fcff0dfdebadbf16dbbc563dac06229342eb4255db90ecbb69f9aa9eda5795c020cebe14f35cc5aa34d8c20ba5708401645142ef9c78fe07502b7690cfefa4a51065a2f52c17c917f19a72e92338ed63007b62636da432684719f617dea4dc5657967e6abbcbad439fdf17f3108935d2353b09788bf1b1124a77138ae266425f238645598eeba4677cbe9f7dbdf6719e8a4dd96fd980f5e2ee44343d5636505a447b3c18c2bd40eec12ff2d3c6db39e97ff84fbf4600ddbf5c1511818b26d6b3a555980a7ceefd0c5529dc716804eee3763408880c2d0d849d1af6b6985ceb17a9c64ddb0cb39d4da14968406d32da856494530f2ba4117faef496c501320baad89d18529a3eeb63a3495849d033162f2c8396c35f0d5131088ce0805c0e57ab0858de61e25ef9d2b9d24824d70408aad5984dc28db80badc64c18c9fc4988ba6516be1f7a5a5d766;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he6c46abc7d00443003e59196fdc5223fc5318188326ff54b81b842015df769039f31fbbea08231aeef5c0742523ba6cbf1c2dfe7476c79376b5ec5be5a07e0162bc77070001eec3cd741055cf9a8106ef286d1f28088dcaa0f88ee70bc4bb2fce38bea6001d95d1dde70d25c6abde732113c7a413d877268af70fc5be71272d7ae74da475d5ef2adad6d64e9e9d226766b77c5da0bb40ef337787196923a8e6a35821d202369e733de59991cf34a9e4dec64c134cacba0e8f07e917616ffaba85df3d55552e388fd32cd64cc9bca31c34a40ae2c5a27cdf094fe081d79bdcf06d887c8af2db9530764ea2feec54707de32de38a54ca9182b957f595cb04c22437714f719c8e2080f19c28683e33d3f429b6abb9b23455c21e32385e12bb7153ae23b47ca304e0c2d73adc23c792ef4becb02cd68ad9a03b33d8e3869f93b8eb62085b7da1da977a45f28911f4f118b053d7e44686d33f723aa069d956d793824dabcdcc8e6cb68467ef29140ad83ff7c9c16601d3f06c8ca5eadfb888196d518af22761ddb9f6b2e05d216b7b8c1d4b8f9f9399f07e36187ddf0d9c80b261a813a406678c882fb58821823e8cb8980c27154203a7228e60531f8bb399282bd4ea848eab0e74a22561f1ac48ad7c62c301596a2d9cfecc867f3b4eda6358814c16cc345326715089deeac77180b6a8688ceef127d44d8f182d0bea804f01c9cbbd68b021fad1105add079f91d1d8b8f19a80ba0e0a01cbb241ef9f0153994fed71f7b8c2052f011cdb57d0c330b18194d9785acfdff6db2c736511c57d5424c05ee1e4da02bda256e6b06624aff45e71473676687e4ca79be3af69c1ab69dbda64943242c3b693cfde1a3bee7b91f1f3d7e38213d66db6be2bf14a97fb230c931b3827e485a75ff52d0172be7226ee9aa89e8dc96f432f716b94dda45ebda9d6d2e50ede4745fec13c2882215ac8fcdc616cc485b6b2468f8eaa99df651fb72383db0bb998d82bb61089a2d9a3a81afc529cea0dacd4cad112bcb7a9c11f0c6edc81c0faf134b015cf341de79b3349d885b2d185be4c4112275e9d95e30ef4022f43dc6bcc4a28e74a95b94d841b073e155e9f6be14a8b6181bbb08a7e797da7a73d11b73e5b56aa2dd5e00ddf709b489bf994db83050b62669c55fe9243eea33c58028a3624109ee2024bb8ac2f605c97c7d90c21d4f97ad55b2aaa23de019902e3607fc19b47574f0b8c5130db0ebff3bd5df1f172a5a3c726cf1930e667168c49992f7e2a48d81cf2ec35fb46be94ba68c7ea0ed57748e9a0b7d68e70eba9025930dfb3dd8ff6392d4e2d2b73d00c78aebcbce938bb5496a3ea3b78c8aed5b2e2bca65f78cc647e0f9a25157200c87b023325c4814503a5c2ee3917641382c6e93b390c2dae149edf38add0690a555eccfc3cd33cf496f60958733335ca122;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h2398de1e0de02e16554870795059d3c6f968829169df388e99da0bcd793b5d910fc1801a41498c2aaff8b76d90147e73a318284f205ef318baee4e1df9388ab374f4a84c2f0f24ca1ae2278a088d6eac9eac80fef0c51a52e14ab607ce39b71aadac584a4db29cf7a9c9deb1dd36105f98f1a09cc3bed4700e98c387b7dcece7cf7f5aecfaa369db8b0c51c669a2234446ab527b75fa12859d34f529689196f110804930b8dfb0548c9ea94e0859f3da138fa59d1ccb0eeae9c3f570a8e99b3c513d0ab2810ecf3c57e6f9917a126c5a33a05e1b5e9d06308a8ad27442a94d4f17828be680ccab41b53cdf1ac296eadd8c574aa27491ae5741efd83681f3b6cc16eaa142d04cc838c4a85e29a4d17bf4ee88f433bbedfbf624169ca90326e56211a8ec7ba0d6a7f7e17105837eac09bb36d6c6236e875bdf03b68d8d4c176b685d8e16b3caeb96050628facaf2f71aeb77815d50ccfe51022da2be1db6d0e5ec92e8fae36c04d1e774c6013fd6b9d42d441e28329d037ddd4f226839cfc1f5cccb8a07514d4dc29d4b6017987263146c7a622114c50ca06ef90e38dde0a3c4630fd453cf4623e0191c88139cd4cfd382ad2f39e547e6b5bb73c7673080695475cb3b11d02f81bbe993685569dec2245c86ce95ea82b2df824985a5ef4d3cae785e39c8fad8b7793fc21962e636999ccb2faa1b8d198a67d62d3e73cd2bffc9488e1b813784b73ad8f67ab5dadcd0ebf8e072c6dc014c8df1465494926d4e4ef5c22430fb54436240a4867fc8af3a0566637e0e608de49348def5c189ae19e4002b21ff470bdb1443d53be7f23540d5b64fb5b0cd53355e92ab27c001178680bbb26a7ca8bb346d0b4ec2abc11589c69c11b3700cc83dc6a3cc33d048bd0529681a2d3c4ef8b9039453ac6a86a5d11ff12daa5c36974ead94fc390e1043054724f0210841fba897844a37c68af6584a1a9f4067ffe56e503fd73777cdd24d2667139321bf56611f022f6da4c6b80dfb4ecef43de50796c4271e43a7a318c2a414c1fa0222fb88aec1c49fcc58d1ebffb0f259f1deaa04938188c8adec951d85ddc6fa40cfa85daf85810bc6dd71aedf18cd25dd2f177eae6c0f329ee59193241f907542a35a10f4f2fd4aff435e161a2f947f885c0c1f93a388d4418e268b5d3245659a14f78d811fad0b18a38d15b53ab168b3a0b7269586fd9a1a9848b53a0521530da729bfe479ad7e34e45bfa1e61d8af51b89d3da3703e8b8e5c121eb2a461c31546eddafab1edc385a2a848552465651e54a0da786a103d8b0e91e1213899eb34259c93563f31faa436edaf7506786c4f4f3cc902f9e1afcd9c3c9ed302ebe13e27d928d50c79be4bf1cc9ddb0c00a249f4066e88be5a6dac8aa099d50e8104552a25717ff407ee789e64459e288709c80504d87465c6c37b948d9ddb3f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hcc36f17f3f82fad02b2f81a37780253bc9bf2da16c00ef6351a72f0f96f06e3f4c283f5e9bbcbc4bedd7b7888cd10d5b6400da762cabc34e212e71f159bcb7769e35d8e74f8a79461de6eff851dabe3cd40831e365d2e15f93d8984e9f869bfd360e485b8d1ef3b453bf7f08fbd5f508b89787f992ac32c071fe5f4197d6cbda0ca0f58f1c6127bb19e73d9662d2644b6dbfccdb82e2a31a31f41fea56b640ef12eb996949158884ffb9d1359248977a65bcfe6789418ad78e4854a52267a05bac77613a254ccb77d939d4a27de34441e97901e4c72a8100bbf2de992832fb5fbf1ee6b2b7c31a9f0324613ea44b4b8811286ed0da6096e73f4747ff50e38f9f261adf0e6b40b3620b97dcb088b63869ca0de59da46dc6fe91ac88a566e96234f3a99fd1cd336026b0cdf532188f1a28e732820fd9e4a22c59c368d989ea4be6c9e66da2a7f17b4bb5422b6022279e1edab6279e4baafd30a91b75295eae6519a90581df1a001ad2fadec604892ff98b552977951db3c876ebc68dc30400f427c4dccea0bc0d0043c548797797fbcb8d624f4b08ce6fa948acb72b55aa01f4de69d3dbe7aa0d5e5613f8d0e8a238ae07a03760585a34474dbd6c4d6c5c73683bbed941998ca4dce38bf2bae60d44fe0e0775a66eda5908df5ac678bfa55b4bd794cb656c3cd60350eca1e3cc1516cbd776e4c43f00f800786a0ccf39f215de0cdf29673eac278b0849d9b17db6052ffee63e4d1564840d810bd7eb36551a944fe8b48a81a018e7769868df9a56e960f433c685281ee10cefefd3f0a813a1ae3e308cda3167bc1e8f09fe25dbd72d8c655ceee873f635244b27b267ef9d16b770cc0f5d48a3b7e42100a0cdf1b0aeef20c3476fa3494dbca33792b45fd78c133d0ed96ab050d210c780e01c4565926a4d4d052b4676a712d2a2bd919b9d0b93596b234e486774693149fc1689c78de3ec556fffe7fa28f2303019fb696f0563b37a6927e85401132214cb595817720eca0859e4b30fe588dee825742bdc1f7a40e305dbba298b1f5a0e1d59c354bb8df0187afd7a98ab8fb7c1cc283af64681ed122afbf825c73710deb89b4f3a59a1535168ec10cb584f18509f7cd806d1cf025f9f65f7a0e5ce49a9f534431d0f2b9a34b791eade9bb126a75322e504b4447957517109fd4b0fdf72165955c3bee60522cee8eeddfb70c8fb40857c78374ca88a0734579f6d7a696b7a614279afa80932d1b88165686116cbec6c686cc223d10800f34bcc532404ff228aab00e89abc52a1dff5e0b964fb23ec386f580dfd1c3ba553eabe64edc4ecd988fff378b40eb5e90232ad43aa3ac81c167d70f94fccd19460089ce1674bc65c70bcffd7550d3d2b845736570e50b7cda668954ac3498335318f9dc6a21115cfedf36dbb563c4b164a06307657cb498647600636115a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc498b187e39427b3c4265f8c436277358a452bead04ebb1c333f0ac27cb3afa111a366299727ddcc324553889fd2d3ffe7159eb2b5c3c5f9d169e0b7e2f826c60997212301ec6b71991b99f76cab3dffa3e342e0299c814584217378b74b270e28c6da6bb45d61be4404f69182b80de739fde8e4536f2bd74711ece2f44f1bf532e1f388695001dc79f887f3d2c97bd6ea7052a9077f5b4b7154b0bb574616e5db022ad2dcc0dc3bc527e412cfdd0a43af4ad74293fc30d7c12b861653cbdc66c966dcc703720a34b605577dc27091dc17f24b19615ba23c94502f87205ea64a7874d5502a8c1c5174244667d33b5d88d6d6aef55fbbe74bcea59fc810882d564bc344ad1cd1dacb4da470a79268941c26256e9a02a0326d8c53f068756994b7ab25033a859d6e56c9e3582b40ae61cbcb6bf075b1cf07ce84df2b3c325a7816d8861d04ef4787ce41340a73c0dbc4044e88458ea5622e8486ba20eb79bd12fa225d7079076045962aa209868e371d2d423a341baee2f457fee38765ad12f1dea096c26b4e37a19de57bb541817bae143b7d416fc6c48b8f05c181fd834e958d28a5becf2b20acf532f5fe231b3e99ea6f7c42b4febb152f60f44669e25a9d2847362d6b3828f0aba2d69f1e8e8c07621fb8bceb970669d39476fc981cabf9be1bb9163a270b75c25f4672e70e9b7053e6dc87818e5792966b807b0195b9a2cd714e825346f958f6eaa32e61ce6debae76523dcfcea477f112f719fb80fb05055aeb3a37aba78061b0d607bd5461d3e432fcfddc0390ef7878cfdfc012ec8b1b6fdacd85a9b67b20ec12a1d25bbb99de0aa22c990a417f3aefaf03abbbbdfe0e39b848d98bb3ebec6b7db1baf988b5b6e896fcf5f2b085d1a9d4492aa3f4c160b2d1d946c3a3ba431539e50b88117382830ca1def6ea2791da78d07d1858ee1a575c782c2544eaf7f42b3a39e8967b811333ed5ec0149c772f18257cf1f7d28cf23cf22a8230dc2f2a5f7f28bd62c023956432ec9b95d91680593120f50598c6489c9e83c24350af48a11dbb8397d875549a689f726eebda307f52c1ffdb8b9b52b60b9f6be4bdfb0a75effb34b51c87c284e1b0917314955d8da5cb193782d31573b381bec0dd3c557b10c03542fcbae07fa400bb79de7149371e9f46d91c9ca186d5024935f27f75735ff0c47fded4cbdfab56585cbb90f7a8314dac8af51b6798ff847c85a2316f4083c91c2be38173c2f7cf56a352af8178dc8ea198847cde68f81ec366e1388fb26b3a8814354cecc5c9c78753cca68f32902ea82a0e7c9b11089bb1ef5a80ed68e5bbd296b5ba372b9ac17cac7369b766be21030791f64ed74a0c1f8bb7b0c56bcb98d1609f8ddb91412f81aee6887122e785618877898d0afd420ad5daea2a6f9a6e32a527eb6606766b854285936eee2a4bcdd7ef0f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf3951a589a75645582dd543aec5de41f9dfac703dd00313c259986a2570442047011dc9c1665cfd23d514228dc4ca30d8354493757a70c8eb8b8a47b9321cb4914fb5d7e5a4b9fcc760c7d24d1515a1d85aab8281b2a2f8c6d521bbad7a783ae3753425b0d7b7920fa24c7f44f8e0643d57e2f0a92b80fa1ed6bdd325f8c18405bba89724d567f8f5c0a4390fa1e7d7c1427ba34113b5859d96292271c8d880b4fc7257d78c3d55b2098421ede11ff1bf2679c157dd39395a5674b89400c1b88d810a1a0ef3e5e187945dbf5b6ed2911464f70ed4061d70e310b6eb314445cb30e8f1620eae91d4f9bb846a9a232b67059c1b0ec73a72903e7e3eec4bc6b6810ca3944ee128edff80184b6e4d66f449ff7bb49204fafe61cf7e441b7c2c940abc1b751798af05d828afab236c674a752f15b56c3a738a7bd8c717ad44b5756817e508dca78e42fbe366f776d6ab17017eb1da848bfcd71aa023c297e6fafabf0b795bd97d48071380453cfc2ee6f39e1ffb0851469b7ebbdadc3f8555a6c304749492b49f560151c8a3acbe433d0bf041a9aa626177a49d85fdc1c93d067f3e53de33388fcada9edf6810e3cd1fdfe3191177cf571f58f227985d2df2a828fdb9a713c4d4e02c0bb4a8bedcc863fc72020efa02dce7c58230ff96c13e333e9871c3129e7e63e801a77a484429ce22e3c58e165f4cf7093f97bc7bb304e32e1970df1e02d7185693f5d29f86b098ce8b3f7845e071db7159a9a448233e1324316fbce27ffb733943c6fb9bc89aa7f69d1552bf1780a3f49b9b01c0b7767ba892045b5d4997a5ea09f479df8de0710253ca602955db56acf6269fc3fcf81c5fe7f4e7759209d8da1751d73fa95feebdccc332f95c7f90c2fa549c1082d8995d92cf1109ab6b9e97a00fa8c728afe55231b7c88858dfb642478ec89b8571b995d6b9a11321214f57601144533a9305326e4ff96a78666957a550b26013a23ad0b1dea923de45041d4c1d29cd64196871f9cd65c0d8509eca44b8ea8cc0e25d90149e9128dfcfc9e535a803061dafdb810d087476f71ae2c8f58ad12096de702090f3e2a05866adecc5230d061d1d398d7b17fa6e3ae770568dcb320e9dcddbb4ef6c724439d82dc408432de08afe60eb947f0d1cc5586d1c587069d1d1ab970432e67a3bb0d7641fc048039b8c9cb0d640197ba70df0b17a60a39f88ad919d41ff7ac4e33fe414d01ffb7989e9fea76f8b65113f4d6e9c7c8097cc02bc399c8fc942c93f5d1d1a71d6265050fc169f57c89e6104166dc2d7cd9933dcc14b0636e3cde34f7ad71f7919931e3677f57d322ac2ac5ed78bc83b8163532f171f7dc3f5caf4698e41f40693f7c20a2122828ea0bcdbbd280cc98d890b9540f1c0cc46ed7b5db9e14b0d438c8bf52bd7e4a156b263ec3aaedc5853641685098b2d937d95c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'haa90899a9e126e489c05eae262b930d5a0ce56b00cb452b51bce5605ba3142a350bac1d1218cf47a45d87fa8c6ba7d7795a5c0a83116a044826d84701aed500ccb459d3a8b122cbcb2b93bfda88170bbe1bb8c8637f7dbadaa07669cff7011c9463205cea0320a0494ac4d109909e7d9be02755ff2e2e13f916d8feae8ec9b0b4dbba26eb9f883e8d48afbab10aa809c22c882b31c9013ea9fefd54d74657ec6dec5bee317dad875cd1fc088f2cfab0adbb4391c0e7b648ff2bfa466a0c0a6989a0e6ed70c16cacda74bbabd062ba9d43f2f8cc313876669410a1f2494bae15747597cb7e81734415bda6365dd979d2c622b12b82d09755297e2281e6e3c4e73ca9b551b9af098f507402cf0754150736a5452b06fe2cbe40137d5714e3f561ebc7808e061e34b52038907d075dab9392458d4ae18ba48860baf5cdb02c7a94bfab0c41847480d8cc2ed7f8feaf47a9aa7f1814934c1540ebdb5ebe470d19ab790bca0f5c77cd50f1efa42e78b07720620e159fd5263223e5f64eb5ab5e54a5faadaa0c749e3e71cee5f8485d9120e4e9454913811d65e531eefb1144ad7d92583cfeb3983dd16b4193159bb7d238b155d9e145e625024ab33e5cc3d25bf69b7cf7f4680cf0ffb100caf4742a1c59c769365e0d49c57ac5de8cb48e4d8de864d59d3911989df5cd627d1d88fddb9604380f823a9d24ec8b94436f2baf1673cd29e00edde209dc2196c47dcc0e3eca3748dc877f0d7612d876dbb3f6babe8394a4444f838f742ba20d3eace8ae1501944b4f19c8cb84a749ce3970887ee0821742e8fcbc8b8821e2b6ac2eee3f3d8761e26e7e12aa0adf365bff37e0f0544c2579b02db07abc26f4c7661f0a5aef7dcbf759e2be68d3bbb0139f9cbb7f49bee1b74af4ead03e38b4c81911b3856917d7bf709a3ae71fca65afdc1fd42a9fbbeedf6a58e51d33bedd221ee07469695e8963d2d2880a41e8ba39c4cfe3e3b788affbe9c8bf7c38ee48a0dccf6a137a04905c978c602d102a1d1725d031d8de3dfda833527a5a21034bb89d6e0c7caa65ab3933aa0cfb829897c081552448d7038ec0ef7dd7257bab5ee3dfa395add1a480f523be90b86535561bea55b46dc93f20515f07da63f7e286da49a0103c0ee5d01ee6035711eee8d28b5be6fa2b8a746264a0558dced887c4399fe21520132fe424933c062b9fb9cda827c9dc0cd9b6328a2777c997d7e61e4a819b5c864402ba24d58207d2fd7dcc10fa7ef318cb1c1cea2775733544e806c7bcebd0af067d020842bca911093842826eba1c21193755db12a51fa3aeb5e70707fc4e49d765331faeca2b089116f747e7779d91db6bbd5d4d11ebfef055f25df21cd8921391b6026131fb1f2c596b9e9795ba6ff26ddcd1a70b90d3070b3bb023b578a080194a198520e7d1b6294e68bc757979ce6854a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h23625c7e3af78bf8124aa173c78d6c43ce20548b19c1d741a51aa305045611d74e7a0649f8b7a75df1a59f17a01572acf31a9815dc23fa483e2214c7e2b6531e1c6975bbdda69e04cccf1402c2c6d63123b80a7ae69a7d06bc24e61fca569b2530906db2cad1a9e19e38b3ba6e24dccade257ecdc7f006d126bed3aa3a2ab9eaf7098d2d950b9cdf03a05ba6deda9e87d2adc4c81beeb2ad899f2e0f5278c49095917ce9686d1d0bf8c4d7aa56fb5b3abc208eec2b6b3e7f5b758fcc75ec34e540e95a839a7d87aec240f61436b488f7fc87ec4e8bf0db6d3a44a9cbf6f6425a3d6c24ebbe87bbfcd5f4468437cac2ab5084756a6514e46afbd24cc5598bc973f173d10d06415f52b374b66cc72c82bf0d654097237cc48017414485f0bfb21825498e3c13056e77dc973d700e9e3711db4e44518a4b54a6ed2daa96bbed520e120cfd13ecbcf861c22b89d733bb0928c3b3c80c9990b9866b4421738719efa836532baa12ee228c2efc4367019970133acb81ab7b37fc6a6321bc8bbbdf27f22810a499e911aaf7df6d8760d81b7a2099744d0ea2d400d6169a18f32e2de12863105556d4e835e43101ceed1ea5a443b24f6c5d0be8824c3e8b654db5c38c3cc369ce01f134d28f75885b54fbfe04b898a17ccbe34e325cb48081fd439e8540b32a3c82a4d95d62730801071d374ffd50539a756111cc5ef0c2c47a9aadf2ad65114f436b9bfab29654cfa4e08cecd4b0baf357a5b7a67b5b9c220155dfd84a80b6360d8747a9446d56e46e29007e55e585dfc4e4f658fab8be4d211719b9a5eefe23ea24bc789e193b936d73001002900465f5e6e01c84061bfa151d8e110ca3dbe13b812128813e029e777aba7e8073d890fb49c56bcfef1d6bd23e54ccc59214b8cc8c9715730dc1bfa3dbd47c693bac2a1b0337ab6282d194356f060c11e7e4f79983735de3cb76781785fd11c208f71db2834f261c8047921794c8b7597af6b065728ab33d222c42aeb819542e48dc13cf42cb7ac1cb5d93d537a016454cc2273d7b82bbeba0ba87110ffe5ab9fb7c2ce012695fe188ea537e92d98851b4d57607f9cf190644a6232ee032326ad4f20d93ce5a8e87367f9f217adb869a866edf922cc66c2e2269dcc610d51e8862a5b8483b49d890b6204c0e62dcdafa21e74351d40064c10ce6330841d2c21bdfa4bf7e03672d494520ff8b7d7f018338be51c0cdedb69259690a27c05bdfa5be0f3503a5592d0bc7b44f331b50a1da56ed86a491f57c24ff1c4c57efb5d1b93c37583d2a1e521bb8e120ca2f071d8b5b0f1bbf1d69fe5288ddb3674fd63db9720ebff58633fa2e32b3a4db3bc769aa2411451136740eda980de0d6f3ceb5cb620e9665fa774d1d0f2912f80361fa71d0b6ed1b2daa6cdfa7f8e8552a06bed55eb85994fd722b24dffa1064f30b3b59;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h549f9cd04ef7a54101835ebbf4bee9f22020d6f6080018e47393676c06657f04a1fd3c2382fd140d565e2b84f7f3f9ce4babdec34bf465405cf2e8d3ff61ef9126cced7dd43840743a1df954280fbf94828a78a1ef7e4e1248dd3e2f515e9dee9f90e70852caa9674a2d9f61224630ba79e9310e5d103b69dc292a10a1a0c73092176fea050566502d615bf1a1cfb5eef1a3a81a7e6b4488436b3f5950401538e102d200dcad209e19e394556e323e2d795a2cef1927b86377819406d242c3f9b2331294aa9cf9171ffb179dbaad96615e9a8873834400a3e6d37676f2d1f960c562686d5002fccf51c707b51e2cf1a96baf7d8a4b022ec9b319791df73c7ca1f24752a0d87468d887bc650fa9ced58d082389d3bd26c0dfb36abda79b2caf6bc0050860b22d5d7669f986ec21f36074197ec081f7e28f5eaa061eb38e55c84deda9481397b004898db145a7452b613dd97a9ec8b89f6572b74132940f9016e79f29f4b4ac80802abc149eb46394485c9550417790d932d6ffdeb7c094d4fa8a5cc674cb7b9da21a7c2989df1885c3b2ee88d656f3800799a9dc8d082ee012f53a78ca849c87e57c05ad802eb185edcf4262bbadc43c86a3eb06ee2a96ebb2e8f695f11970be89a3c00550a13f5ef8d707e666dbb6a3778211087721dfb6ae71cf84819cfdd41518e64ff0a447957da8308dd47b7627c8c0797009eb06f829873045c219e754a99839097f81ce351e37b27121010ea0fe692e4d250ef988565d3b4e3a19a51835a5f3d109bc9c741e8d203eec4ccbc292a4d2d02c9599cc7f2025428df2b0405f578f9f57762feeb7b6a4dd1e0de5ac01ff7760f5bdab60a233371d1d0294064d6d45234f61335d3c213de2580425c2c3e8b299f3c12e78ce093d7c5157e4e23d7ad21d14238044f04a6e298d4826f49028fb3ad3f33d4d9075acb88d793ef3e665c0c276a15a51b44214fe009992b3707129a76a5e7d3332d5d869dd21c986ed17468068d65aa5028c1116275479d54206be9037c738a1ca43b31710207de8e3f72aff2e1f62b8d5130a1c628436f7c35420cf839172a6c484b1d98c5f5580072af53e427e656500e72a949e300596ae6f789e5b947238bbfcf54187dc22999ce32f61fed643017008ce44503da1e2aa6fcc16590cd8958d2c93294b53305a5326e7db1ca46066f4c95e321be65364367a672d6cd23decaa4c392456c686c66c87e51aac014b4bab352e967b3913f1297a5e49dde7ad3bdd3e9ecbc1b48dca6a82059c9756a31131b3eb660f08405f330118934377c91be7ed80ae5ce3c77c6c607d9aa79c4a745c051a901b0a9750d377bb22db9521ab7d6ee463a8e385126e1d34c8eaa86659ed849204c50aab03a54cfb539476cf060724693182c69c492c3967d4e87b033b03037aaf24fc5cfea73a33552223f3bb34d8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h655a7dced14e1d65cb5fc64c37f43546f63be035f8242c69cb73b5f32ae5738eda6da5c5517f1c277a4de71f28a5e5de6eb0dfc4e8f19bfc5855b53731e67f512bb0d4ff34cfa7f05adc4c14d2f9dad9f3d88cb458bbccd6812c0889796bee374c84cd32c5c98f002dabdea3d6004f669f02287cf5fc94c4c5fcc6a1d7a3cebd646244e9bd8dd06c48da0df7eb458faae9e678697c87251dfa47415467d5af9410ff74a6f5d321955032fd7fa29cb3956c69d9c1232db96c2e3365b5630e5a5ec2ec8311468b6c1ae49d07305048f5c80241a09b0884d4184b86890c5673d0589811cc7b67877f4e65c49e25466fe20e87ccc4cfc5c71839fea7b3e01f152be1d645fa85b9d2ec7ee6dfa094685844338f7b0ec21e1aa3fd231c7f743a3201bc78757bbcc386bd2c3fc4a98d11e4d55a7c34d22440bcce7b83751f0dcc7249bad80417b53fa2051a493a773cc34d886e6733b1b69f53196a167ec13bfbf5c374ce0f9968d91e67e07b871c58121e16d9b759418d12c760cae64c860cc3f70f80076f2e08edb0a6e7c66cc27cd24f8a706dc17556f4421a8fd8f12538d806a365d1b0cef24e03aca78389f3bfd88959f6d7755e794e9103e0ba11f53dc603999e7b4ddd9bb950e7ac0a55107611fd145a978a0023f2cf8ae69b192d1ef6c5e7fa3aaa19cc8b34d7784e332ad45e93acbf8be772e912e370b4d8744e0a456d94ce4cf332a41c5af0cb1061ba443c5c06879c51b2dd8b796fbc714d4f796c4daa6001d789648a22d237427f77c54d8a5afb135a4568e5baff09f068b865b9fe5227480431725493faf46c215b0e99d4957b4632fa4279ddd8483bbe2ce9611651811bd000fdd1dbfb3ec76c3ff837220c75272ccb8b1dfffaf775a426e9a2d7aef4afdd7b2dc4741a05231e24657199e40d1edee9097902ac3d5ef299b31a51eade7eb29447fa5767aaebcb6e97b1638902cb6b28d0dd48a94efea74951b3d14cc0e4acf3a66d8d44a1271cad8e3f40eacad5ae5af9240d8b203e9cc89e906da371235434dbf3e55e931bb5c7e4616e6f362db3e04a8c92da56e674de5066c29baeb605f664cc5ab8df0a3902786cad62c8b329191ca231db1582174f9319c82bfe863669570b341ab94d6e40458621b1c031471f315e695443b9169875c829fff92d42448e212485d7af77b817e09a2040ed72381c58f552483df9d2428b53bae6e8e87b39a629678d8d43ab874522a993bac7325a7f0108e03f3ae3d962414c5bc3f0232ad3c5aeac40c1fb125a62ebc73c66367c82c25f3b3cf02e8605ef0e6c13855ec29c1cb69105f710b22d6ad386f791b7a82619e831b53dbc764cb0dc997286320e80240d38a669ea1ff420c2d03a75da18d23a51d9fd7eac94b3eb36dd9e18ac2707a88774b67e63534c6e06842c4cc8ecc782539155d22ae9ddb5922b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8c6d12c98ca931fdba9ce38e014d9885ba8ad1b44b8776df61bc5c5313ede4784130d572d052bc2d3d3bda0b01ff085b9657ea2a46ba0ed6cd22f5b568e2e16cb2d98f68141bf63b98181738e18f58513a127dd56a8193dd42223fc2e801827b1c1705e9e7fad11a184b9969b11487e7fc5c7920477dc0196b1bb36dcac3f326c006d2b4d7860746e30dcd3e05fcc56403b4b66efe2fadb96cfd5095944d296e34ba37ce1730148559de46b00f4ae6fbf95e6d25101c249def10be1e092deaa665c630566934a415894f93715c8c51a0ba9c351e5f2b6aea6f29030652f6b5e1c8fd394c96332bf0aec0095f9faca03b01075a9a91f554c7021c873fc5608d0397943a10f5080de61402986f4e87f22e6393cac12cffa32d1ec97864b091b6fc1522f1335931271747157f94aa06e33a4a6a4a40698c134626f9cfda51b97549f5ec6e8101d87aa4cb917bd4fd539ea101f5655998e8a6eac9d4b0ec14b8a3e4a5ec0ed9898c6a0ef733fe9b29b8db41e0c6c0ca6a1ab2ffa45383f6c22fa00f952b80eee9d170cd1915b33a250056551356c48db1dbf0a13b7cc9683138dde23d71a69200c9a4704ffce7569fa0c05bcc8ad815c13fd9d2f94cd8b0b5927bf47576a4f06d5e4f7f30dd30f3927ea8e70324384f6bd99d83ae45df50fa15b48e3fb2fd238b54f3587e17dc025c0af1d1478a9093a4f29400b9c048c49884db98671e7aaab89926775d54272a9efae46a89541f26ead070aa89e2bd79067b58340455cf9483686ca4b5e8498faf88dae1ff476233eca3acb720be95164f0c748b99aade317b796d61e891e017e990579e82e26a8c817c73194ec20b617499b327ada5280d0bcf1bfa3cc41aa0ceb1c37bf15322fced35462d7a111479a89c3ce556050334a09da9cf9437314fdbbfd16e99a5e9f7ae25199cef964e09e6e22aab2697be6c9741a7bceb7541173992d1f92163075dbb033ff5a5509907fda8e8e32acd37fbfaa7de24ec2e028c3f5ec413497b285efd14cfc022c274d8841c97cdecf2b27df5b7d915fbe73eb133d362140624c4e65d54ea0fabd00bfe565b998db692c2b4c2286f2c896539f1ddaa7d6ae7bbf52f18a5ec74119d85e56a82f36da17e71bde2e3a136aaf303e3ad3591a5e3b92ce6bf410107e56c26aa188ef0a77487df3de390fb585f791c1c68f83d2fe54ef3d6e848e66ea61b9af0fcdd5b4f2068c1da0bf9bd337add599fda5bce839846a4b7ff1019d0c069d0689ba951b71c737f903804b8fdb60c9951a3450557053156336bddf94d90d0634e373a5852cafc942176b78cb602d7a649c2b9d5b6664ae9ccf81d47f6475f6ff3f0df34b734e5baa3e91b9e48803ab3239929867e9d2f035645687c3afe6d44fb3e310b967b9fb6384f686b06e62e43e35fbb34dd8b71ace24dbab557a125c2dcac056344;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h592dccc5a22c93d3516f59f424c52d9bcdd613ff463b9577d52fa95291238df5a79b3a4c72768a733b29b0883c34c020b98062d44b695ac99e71263bd72a1d65fe9b49d192f8bd822887c1d7f4e65ad10b6d4c587fa1eb75bc09a001d407678b2b50f56a61b259814ee3b3d210c41b12cc7a22434aafd18dfd40204cb8a49fd33ccf9bcc4f1b344f77e0d5315ea1b210d500f8f992916738b25922cb717a6d76410588c4f91e12041e36c81e298d968af2c3b2f8bdce1d0a4f45e9d1dd29178fa51a5b8434f5f650d32b8ccebcb67da05989ef5ea24afa53e6077c27aa94c9ec9bfe10c4a13f4dc827e703d5f388ccf9c82503cacde62390d962511ada463879309fe4daf5215fc0855ab68c7ceb9ff2d250a417aa826a505df6426145fd79b7edf37c4ffc2f540215b36008a27142069305de274823b25a03ef8f8dddd3ce6af2c2cd7ae8c84f3027ddb4ac41ff305e639b649a1e33efa2a52145ea4c2c8c3ae84c57bfd262dcf979e301edba1f8039d27ed6c61e68b30a2d6050709fe26da3c0a0d465f382c3678327618a269fd86d79427791c36b16d4a0ce17abfbdee8577b71abf830ca966a837e50916bda70943989fb93debfae1eb5dd41a54ffab748d5a93e8c05956f20fc43516cb701e4cf216e41ed613d2a5e95cdce5297b8e109c4367fa95d46d67560aacb159a9fcf64219d25ea6e68049d3465315eb3811b831979a2c86ce382e0a55abdeecdf676b7a3514ea387148535fa1b25ac64adcd716af020f53cc4550193fd7780212f2950fa639976ebf1df77ae2e895055adcc9eafc0d41aaa62537dc643696a6c0202ae76ac1ab2a4da2e174945c9610bb8cd2da4ef2ae98fe40f90e66c7d9074f2d6c24cf2a073909e9dd13bc1e839426281440cc16405f75135e78f430e7807f7b0bd42e12cf01ab0bccba8b8e8ce1f62f2ecd5cc7d34fc319248693d2131bf9d9d2d21d3f4fa906671a5a60a9a5277115a3b317f42b8944c739594babe41384e58c382fb191683ac9c8a3cf488ff1e940edc2cd9679f38ff7939f0ad17ca300cca02cfc699de0b6e2a96beecd18c42dbe9efd672a689c72b08cf7cd0b1d427a445adf8388603d203ef002d119ace5da48cb433d597283f1dfc116754bbe1970907a73e8f7106e4441453254f7b7a58b296d83068efe9281e5a14fce8d6c0939d779fdb564708a39c225fbec7ff8bebecb9f2772972e8e9508077f4a306052ca90f683c75278d242ab5abbd2fc70de86cee5626cfb8720a9ff09f357f5ee3aeba95e7f14d39f3f19dabc937fd3cc3037ed708e0f9c6ec43b6d6c88acab6cc6c42b6408cd38ab3c3596b51e43c9e8574a4ad5295b3cd7cb0a84a2460c4d92f56457078d63db2e9714430728d77d90a5e37e966c756e0b70bf19915dc6cd2a11867d928a866917dc5ab801c86f4d99e03992a04;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h14f09518e68210f300bdb029d5991386bec800eb04cefae3d9a9b2fd0ec63ad4bc17b632558f17403317643cc885a85c7748949e52f5c10a7e87f08bf0728e1c80878b073cbe1257b2b9c6c1f94b7e84166fcdc1857b2cd51cb36be6fc5f9f83e4120d3ee559fcd21320430500ed600f33c7ddeefe6bd10d9148959ce9c8d2b5af72e67026f2f3b2f39dd1dc7764640b9dd1b59d6f164118487e50657afd47444e22126fc7f3a019389bab0621fb8d2ccf52869e4672ce69f7b177e98a95f11fc60821d3979d5c0521ecde86c2b679b4e3e6a60a35e8bd93cd5befe081b80b88338b253dea39a7bfc86f7693ff33d8269bbdd211a7244d70b159496d31805a62c495759677b0f0c7a89496fb24a740ec77d47eced57e3b3398daaaf00c880030a4e248c527a99e0fffb2ead05922714a87122e136e1eea141a88f48b220cf8f70a893cf30190c20dbe4298b1bc8915eec1659f23d08f0dc6aa1fa31945bb21cd5d41daea7a753e9888dea772c2bf9c25134c5f8d39b1b761fccb4c669e59df7b67dd7ec6c7046713c6c905502e4f339f32ecc67045aa93540a062809f90ffe3a11b6d56bb494b5d6871b44d7669475cd706bdc3634cb2248dfe5caab8bd9aa69e346c929d0f229f357c5d94c3475c884b5ce29bad27758d8cd810003cc9ba8b96802ddaed2a6dfe3a18392c23c22536443f4072d2ebb58bd408510a9b803bc184fc2b5b0095f3ecba16e1efefb5093139efed9fbd7fac65d0012b97b768e841a395c6619e314db9742f400cb4cd44123bc9bfc541340257a986f0ab610ba0ad9485a8933e6db6cc9d5f90a2251de23c9f0873b690f815bacac5a6b666d28f6ccb887125ce3816ebc0756034642512a5b21881b3af189b61401d2ea497c970befdfae094cf8b2fd1348550a5c96d2a9ee822a9fcfed9aaeabcbb15dbad3dfd25e40efdbe5785886f3852f14c9998f23150003cfe44944539f618481bfccb27798bf2879eb76fd9d72c5747f18737e9eb520d3af1eb99af136357ca933097668f9fcfe20b50e010de7b571860f3f30d80df22eff325c7d2b6ec340bb0f5d5c05b0e0afb5f3e9126a80f4a2e24465aa9b725e1f7d7d54417e41941c2818550f9b867bcab159d105a5524a7c5377b12fa91042b58f4d8e182b0e9fe1b4e15811a223e750ce5f2ed8c9bb4f7ed0e2cff5303833860cd040b6fd4fce236856b765ebd8ef5a052cba95382d8d5a965b4f38c2ef5d067ac2b580ed1da3fe38824d61d709b99c4d23f3791d4899e2b10eb801f99a2f8bcf15f4b97a535d9cb16bdbae9dceb620a167d36962d7a6f6c75dc3d7ab1bdac13fc8c57facdd0f83a131753499401f5d8e90a426120df0327569e9850cd2b2549234cf3a19dba34935c6cedfc35e4d238900af93d40d6c01c8c221286074fd5ba73e84f7e298a1be3ef32d1bc667;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc59ad0195c4cbccd4308beaee7401dfea7478d730cb806d5b56a2dc64a1f6c75e5f7516c381959d335ea200fae3ae7eb5a31c9f26675c36a5e91bec6629eb05de7b2be31ad020ad8e80eccb82fa9f3a8616b515b22fbe5777790e223eb7eaa1676c862c06a4f75aa50f995e514e57d25ae74c19a0f5603ec522ca5abfc6abc3ef28aebe8924247ddc69e7a0d99f30f903923ef6d899e5eb6faedc2dbf05a8cb055ea16538e191863a75142f0a9760a83d4f0212b8104908438ae683b693e2f50ce29f89e4f2c6570dac3c304af16f89408d2136eafdba0ff2ad66366922b6f2a1b0325fea22ec486ac5c18dbe059162b34e4ee1cc68ecc129e73d69c564fe5130d0ba9a7ac62aa6b0f246f1feb5adeb857315d755e537a180da91de552aba4d27b7fdd8f92d992852906c7f7882c43eab8884b6d787ed55cf3b9bab69112f43809572487ab30e4475eb2d4faea6ca6b8475530a1c255a14a46ddda035e1ef7f082ece9f3207492fbf6f704a4d7c9c9e5770521d8a190f735719725ed9cd3a9442ef4f142f888e6b3fd87f4694581e77ca1867d27fe2de1ad5138800f00202f0a394af232be22795e40d43e269647fe5a8dcd71c234c60993969d8957eb039da80d4a372a0a7a08b8fd72cb4018ff6233b3ec50796ba1ee958aa68077e7e3f32d78d6ec6e5fd3bba993b994d2201cafaa702ef044384e7408665a7c0fecaef8fa921efc66589ec827f055476a2e52aceb490b0a4dd58f055cb633c37736e30f78db7cb8569a5f575d243dfbdf8407eb03761f75615ba3802a734cbbbab462346551fd5df905f2457d2178a16681837086639612c528f6f843c286933e9146b8f1bb946df8edc464f745886905a3465ee96afd656e480c354b380ebe3d71e7821037a433e5bfb394c690e350de766f56e42fc524d20fefd2679901571a524dfd050987c5082ccdb6ae01a04c53270541125aa19ddf8e6fdc6ff677c524f799884c455964f8c00cf7a29b2d92dd56ed0d9caa97729ee49ce799c3e9ac7958fa2a5bd761a9ad2b1a5b76f8f85ce4f020abea3926f6a635761373b61ff53153c4495934f1ddd81d3a224df56fbcf3ac9c21b5755e3c2f114c316aac2401ad1f41a3db14bb354a85572a1a533d3ab5b117d85b1ebe48c4d8e238a091e6d4395965f529a54e996250fcb55f7e1e950ff86b0c91b227c2cb789bf424432885b3d47740a586f0fdcbbc35132e99cba8608625176b971e4b793a7d6da9987119000159676314b1331d185d012aac78dcc620d4bc9b285bf6682a28db3d34efd566b18e0ea3f20e93469a81a37bd2d8d65664ea192ae44a265eb66f7b5d4e8ad195edb418c8dd523cb58f93fbeef3e496cc9f421b071bfc5dcd2f09cb416f401459051325e075c296e5298ba7c03a9310969ec9e3f18b1f5da2f8db41400d108375f600f69f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha23f54a4c249d3b077993cc61ebd0338ea667e62893be3349984f8b388fab80aca0ef27c8492518547e1a52cb0630f93f6512613a614dfa627e8b4c2f35d53de19469bfd6fceabad1456a8d7111e0de1f9c7e7bae01093bfdd11297dccdb85f5260f55792cb081385a9747dd784343fe969c77926d8968b1797722652ed11a071d7f811c00d504b249341ab1207a798ceaa9eef070e0f883b5a350717a59357cf65a520cac9831802bc18654bceb9417b402b6679ccefbe399dda94416b8da92759198c5d080deb937c19ea1b17e063578123b385040cab51c7dd7952a66609c6be57ad8d61200d416a5bfd50fccb10a553aa676a630ea282b3937562f31bff43452c32c11c343b55c9a58d4f2974c1e4f30ce2ea296170551c20c7ca99976f30e786db9d1f904fb335c9bad6566b9c4f47893affda462fdbed2b8a3eafca0030372c377298f36e22ecbdf7a8a002be3d9585b294c6cc3e9d859cd54a49c4195526a7cf6058615bf7db2b217546304fd4671c46ad87882a9e23c2caa2fb6748b518e0754f490473821ca079eb6f3d0e2de35954379a1d1b75f7d4742a0086c92d5ff6939229cdf6a46a27258ce7e4b429e14c1d0dac9bc53281f89da499f0879f76da2f9625c6e284c85a10d08dfe6d9641ad7c2fff61e347d6454f1fdaa93b0b36c798bceec1b858f26a153a4a750df5fb62924c4e6ce0c67ca84cdb3021c88f09d702e70323929017225e16b2e4ba6497e652ef4bd9e38f7e1ebaea7ae20937ce4b7d663063ff64fb8f703760e6e84b6b5fc037c636e266cc8033500a7bad327319bbd1a97c065e7b292e340500eee1f13f6b69fb1f4ac006db2cb34dfcfb238cbe8dd022bd06a5b35d29aed28f4664a723b37c6663ace7d7f480fbb9fda42035fee215dfc929ad115c921fb4f95402db2215264c8fa0e3e1ea5650a49183446486780235ca47d1e26c903e66119340d3de07aad8776692a6dfc815fef2272dcd746e815eda928e8e64dd08fb71ad7a3fd95c1a4b6c9d3f021564adc6cfc0e0783a60b26cf730ac8492505d44564ae987a15b0048943fd957dce0a6b19833f01be73f84c0eb6b0df73a76562146c2f077c3ce7b20e087c585c74720177dc5745c8109aab4759e6fc96d1f1aa50a118c46630d1377501c0e4f550173ebba331e3d5597e7c904a41953796083fb445bfb40a77044ad3b6d7494f178b7c36aa486ff6414928ab8014d3119932dbaf6efb9ad5ed0673533283d448b0dec55261740ac456aaf8147579d000eaf13b8d9fd557c7115d1582df0c85d292b1a504e482508171275e126da838c4ec8b4c2fb08a1508ef8bc18d06177815235bca404b67e9089d84e799adb84c9b825cce2ae66e2fa447e4a8e79d7881b7fe5ddf6f4a8cbfb0573db0d355ffc931d8fcee5b2e0f7932fb19668c1edb938689490a6116f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h32dd9e9b51804cca305bad3ba789096ee75bf493c5b334b552a680c023c2c289a9c2c388c839c89e4ba2527581313a4f68fc5aa3210088d469d5d3669de6bf33d03baa5d971634873268dfd93410352be683dadef9c59b209b5436883bf33f2bc91a4adaba17a55576d56f3f546148fc9a1ecf756da9557b75fdfd1a7b308bf147a1a65a1aa38b369bee893d33c8f88f796b6cf24a8d8fe04ca617c88be173f7ae43f68caddfa3a05fb1a110bb343193da9588b7faf996c69e46dc2dc02a53c4de19ad00ad8616bfb0195d3878c2f890c51bf81a2cb6332bacc5aecee0673a5ce9303b74aa081ca537fb350b5520549d8de4da75e20e938b7ecb0f715bc9ae0c36e2659268b1dac1c52c4342412741e96b4015723cc7c511910db6d624bbc539e792cfbc1d61db36ae8075962bcb812fcc3e99e35e2beecb420f44d3e4334adfae3b6aff22db9b36bd19a5b7735bc514938bfa2bb0e49f4868f279e148dd6e524615ae7615022037ed80365ee221d48d1cf7bf7066a8291f8d1e7e483c8135ee9991e8c663b7ef3a3961b5d498563b7dd4e56fddf9508d3d14429573814e2f68d8cd777040765b98e5a9066b2f341c546dbe3db7644ba0e47963f923b96493a671eb7400f72c083f898e8cfe4cc2791b2240adb0e50b17e12968f347c032c861886794e69499aad1bf91efbdd76b4e9ed4075b6a51155fee2dff80ec6f0824cc5c39cfdd0182e361df15d0bff05bb21912a47b01d015082771395f59711c74590f5aab59759ac38473a95681e0152c3b43ec40194cd9864af1b2c82d736912924b93528a9f7e9d3e7254757619bb1cc2ac61a7942a3c5164100e5a29ea981afb8489a7da8372057eaaf3501ea9a7d6638496fdf7ed09d2ec9cf46d4eadbd6e4ffdef5e563bdf1f5a1222a28789daa8bac7221a03f9d047660b1d33d41a01451b4d539493908f69b76d6fad2bb46e9b6538f6f48434346c3789d4763656cce4d1bbb591d7273a287d67cf0e74d9f0ee9344bbc1265fed87356521e27340ffa18e7d14279b523c4f1c5be3ca520a920fc27cbabb8f3101def1588e1c5e0399e957d3346cd0883795964318056d42913c914b55b5b87b4eace417880559968527cad2d8e53ae5ae57ec634eb6c98267b09932ea2bc45f42b7ce9fd2300f11fa91ac3bd551593dbd9b2de52193522cecb9749693267b0703d908658518f47caf7a7ef9b5fa49f0597f8241a7d09d6cb14b3d37c387a4b3a16aae005fd075a1e68a92dc6d983e3e6b9cf8808f08dc6c1c9076c6da60798b4ae5dea1f080493767e17287f94fe0ed5d7f8923b01563110ac831a0034a36551d1234a647560cf9d50da12fc7ce896a1565c83c396a6a1762f4a630b980cc3606f794b31119a2e97758f0e62348747e40d1cba796f67734f0a591265bebfa413ec6ef0007b3c0df70e64e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hab8bd23134877f420449c43a9be48b42161f196da7a2381877aacb0be3e36475553b69866ae35665da0fd324dbbe70378ff1a6e5032f3e82e9d53149dd5c537ea2892bbb20a25f1b44673ce8213afb49da02357c1eca78e5c26a86647a53a0b479a222c3ff5d5f13f0daf8f27ecc481d7216bdbf94f96d6d439c1cf1b220b95e4523987c8fd0a14274fb3f2cbee5808becfef81a5442e59a9d6f9f5cdc02d84fe3459c70c187329cfc011f18da1885ed4ae372c37740aa80735f81d45774e9ae15505538fac76233029c067f3930120aae1b104007cfd8b02c9d236bf474c675c0ae19f038f998eed4372403ca2dd3c6e26be142102b942a9237bcd01768f42ec5489fe7aa2d4970c67d20c0255ce2acf3dea8fc136131926de2b772976bea746f5b0c09d28db57e397d0402c08b119acb497e3eb08b0363f745b7b33909e34a00cddfd3a81c415c9ce582e5f6c56d5acf2adf606310d3ead6f63f268f20607806bfc8dcc72bc6ba8593834c806f325d5a6c919b5ebbea60f2d64f9d65a30ca8fc3268c83e96418566bf4f1ec1098e38a8b6aa3fdc891680e0ff737919494e78bfed4186eace2e59582acaf9503a59e5e0c0d31f3cb610c548e97b2591f4588389c708a503336169973c69e0d2c04b78a5823a1801c129cdf2942d0bb1051b176ea10924fcd4e154aac37c4e32e90b9ba302d3411dc717f7972a578b65da904682cd0ff22d2cd5ab27156e7bbe9387af101dbb37399da449f80f78df582c1da0b450fed27b31094dc8df81252128eba9565d3082569bd6f196018991dd24642ef1ac8b5d0007ca1e52088de51555e3297566984766ab4c1dae6b4b43724bb385490eeaa0be7e649d488c9333ea9b69822fae8fae114382ce614ab122a029fd34b68df9ded26a0b6e85727647453ce73aa01a3cfdc2c565a8e1cd71b8c1a27f98792fcf7391f85d9537d2e9913c0d692712a68dbc8d4c6aec5f7bfe7c322d5cfaa62e1c1bb9ac11e480c517170588ce0c47b783ce5070e40cb0ed011b9cb45f4adfb9bec1a42941ef4eeb4c9c5495617bc47e9b493bfea8b6237b872d6a67e37a6d94616e317b988770a69df639e660d4de77bbd5eded95cc6476575100170f558ee33fb370837565bbd446035267602fdefcd2c29ca767fa04c06fb1fcd17f88e54734381adb4723f4d85e504d7a15a0b8061b55f75e1779ef1e801d06d2f8bdaba62b48b5f7ac6f2523c671c2e8b4f9e68110d0a713e642c7ebfdf37ff5738e6c49bf9051f67326a906f4f2a0def9319a755c43e71bbfa6d5b882e4aad7f0ce7999088568eb5832f14d07ac4d5673618295330d47d6668ff0cc7f9771591a05840b280cce0192f2f5d16298b14c433856e4704fb40cd842f73bdfbf246f79ff9244012535c7987a1ddd5e2c7d2bf1830ce821e2b146e334d4d5fb79aa3515e9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3b3015178a5adbb3e2f0460e57862f9da2e7ef7c86e01e2c6efc502bc22ac125d35762422990382966d03f92e04654934f339bea19d282380b59a7b4e7fbc701e3e11728f7d1614ecc0c263138ce37d250bbb02a04f2c05e26e8507d87a6732512f97ac52ad0584b83d13dc19ad10ed2059f7ac22388c31352cecb64a87263acc2c0159bc13ddfc556a3ec530afa7f0f6c8ce4577fa66fec33ff3eb99e15ddb36e36e43d82ffc270c82920acbb1fcb0dde20b1a4439e4823563082cd6e205ab6628c3dd631b23d1e7ae1a70340b24cf05a03124a8ab286b0748b1ebba2d0e7fc89442e1d265202ede9b23f8aa7272051e45313293a9dbf781dba277f8f55a4730db01d3bc3d6db72c9d32cb69971317aa6c10042907b392f0a80ecaee975eddf328b19b247529a4aa3747f0bf1ce99a6b480aea8218a771db7b46ed40b11960d4b16723f48b7317e40832234c4a32f65a58e9e691588067f36bfa798639fc927dff66a976db593debd65ed8a9e18c4aac424b55d25762498a8e1b3970d4f855f006b6d382bf59637ea2508cb940a2eaf44d5dd7cf56b091ae443626182ec9fb7bcf0d7819e614db61fd435a07701d3b383f540b1e38100262183af984fdf6d188a7d8abc89665842b76e2f6ad658fa167ca46da027dd02fa8e34cfa6658d4ed9fa64a564da518f5b3336ae4f54e1572946e0bb3a520aac970292dc965891e98a74da479f7de4b12be2041787c779b9a818c1b4c2b756a4c8307ad693ba4da3c25d9025d8af11946216d0c88f4b4efca6a47767bf5d6d0118d0bffc69ee9f2ea23deecd1dcef5daaae71d28ac95429374079bdf975334a7fd5582d382d41df536b8092e9bb01e107030f65b68d8d771b1454e1ec98508cb0ae6ac23df5466e679070cb152a73e583ee3b94b8fd3a3f20d1d68f1864328679bb7c3ba23f366e5c9e55979a54ecefe22909563eb93fb287792e8defd0b097c24566fbc3b3246f182757150f2087298b250c970f3297d2325d0c906401dae0a3fd09956e7a0493d8d653c769a8882294b0de53f3327c86fc00187830159a40b0ef921a3e2e94a720dc26dd8f3cf5a087a571840a57010f53f7f25b221b4adadd4096e66565d6356fe9d7707ccf4122c4ebff5ae67815860d63f985e3750daf7bea74d99775e4f8202abe75fe52570c17f9291f8cc022ca958a515ab7074a9ab4cdaf46ae2a1414be682040ee74faa5b0665425b2ae04e92586b54d3351b1c2f430c2ed8e7aee405a43bb007a8c9b7722a4ae4ac23d24f1b612e437456e81fb2b69cdd3e368a34b7e653c97cc9b35f8ad28f412ecd14b4cdf58d09cf10a910670c1e1ce49b98b397a49557de556fa92e706b222d4cf15b90cd7d342a8f8f34eeb8dbdee64ac4cae56f7ce8880d9d087b6730e60f4e28ea6a8f1f81f2ec60609921f3f17799b54616;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9a6da3e4f6b695b8f548c2ad63bb1aab06f8e19c1d7b61d313baab0d8a79deecbba3f6d547cab2d4e5b9b1c15243c8006d3db9f9bb5fedd89ffe9990f54bfa8cd9436667c9b810c7aa3ced7ef9efe778b59ab30cc3f507066a46a93c403d8661937e5aefa3e6e368426884892f1e35f0f5e2c3695790fe016878177ee544c4eee09e15504a3408fcbd4bf5409ee6e3399ba7b9eda389d183e771432262136f1830e2ef11d254645ebe893e686e569c56e5c2da2e93432480f13c8f1a457af4909ba1cea12a00b30a286cd076b8119129aad30ebbb90507bb9229ffc9851b1499b0a761c7bf3f8c92b1a71160cab6619998e8a55d1f1a39edce02965b780b871e06bc8b447a76cdb2a8122258dcbf614e55f51e49abc26c96796a5234371f51074d48270a900a762e7aee6ca59cbb2c7dab60453e1ed2176069d9f56aa5a116b406f4c688b68a6d617923a6e15306e345b981b14b4e00699e0656610c7d0317ac6b75208c13c1837d40206caaf7416e84cf3c10054ca587443b48b49d37c40c2ec206efc2d696696278384cdb23d0abb99537f0c5dfb2e009d7a0f786be221c69d3cf767f11a5974050659061ebffa52d58141318d430df5a38957fd4642406fde723f998fddc6e5db47e2507d7319055ffeb08d0cb889487f43557a70d44a3683b3079bf5efb4e50be8641b2f75ad8b892ade1d23d1b330a63a5e6bd5156a86c4949548c5b3f7b8bd2c6058155e0f731192a19825dd056fca358227a86796844b4d63a4dfaf48d37f5f38f7739947ba6b31036d3daff8c04309aa82779721c1aed27ea5cbe5ffc607962a03df560df6da2057fb38b4b7d2925a4ef0bb408177f260617e1e78f4e33802f89d66b38913cd1ad70f16412538201eb585244385cf00a6cf62d90b81f71341c3b2db22aae989b112c3a1fba2bf730f2011a370a905ff84d4b0f03bbeb49f99a02f5bfed214557f4d0af8b6a9db058eeee0c083e9cfde3655ffcef8b11b7f66a6e79bc96b1cbe0a5c3ff74ecbb190b2773b76f5439f6fd62e81514371038e282326b41e8e5c1ada74c888ac8875ed15ca6f771133fe53f3554737171c9513d4143b3a56268332323459416e070d298266dd17084de09fe6d4e62eda376caf1abacb71f099943c34df7cdb003f64433e5a13f8bac1103ebbac86391ada60dfdb8c2487f221035ecee9293692be7732491dbea8419a28377c739ab61bf7099cc92b109c0e64813b15d0b70ca7dc4b86e1c925aa477235037afa88a265bf2fe6d0ee61bb23a234da6dd6d719c9079e4c15467c4dc75fa4bb6cad4feaa1895826213c88f2bc79dc04d91793dcf59a99b5fd5238189e6a8d3d4067ebf6714fe6bc8b56d4fef79b0bcef9c07c07065bc17d30c70642ccaf826d8e71f75223707047b7f91e8d0320c318990f918f93eefba8564e3b7235028da;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hced5023a79e765c661653a18da2c4bb24a317e231f84573bd1c92119f33d922dddba0fec15fc97727fd810cf0f74b57dc730e39ca2ee7c9b2fc87db7990e0f8d9bc8faeeb7ca37de4a1d9bdedb38e98ba60d8095a90c93b9089b7a8e81fa11007d5cd1009a7c6882058c5411612eda48799e1bcaca5e2460a130409506a5eecda31c1758166dfc398823920db98be8ea09912e9f4afdd944409c62781181fb44ad942286897d99ca7e6030211764495353dbfd97f4289ad38d76cc7e76135c0a5178dd92baaa5f0b52688ded343c02983731e2c2bb49a6afc872ad9df144dc6bb6b873ec0fca3b44db2d56247a9ecb7eec92fe876ed6cb1e45cc6b7a07d11dbcff5e34ee6e3fd76cd284a6639d0c7d056d23480cc4ffa0cd34ef744805154d26d7a4ff1b04ea2ef07ddbd69fc1dfd2d79d03809a448d6132bd045abc9806f9c86699ec61b1701c2e0dec6340728c99280949d38c9acd0e67d910da73825e1497cf8d075a03134c159838bf0073295dfa42b01b0df5b4f4a1bea64c07c3fe4f4ff182d1aee9ca5f224337c34612bde1f016924bcb80d048846399f34563b43ab17a6ef3537df5fa21d9e213d265dec9115eb36b7d8cb337805edd66971eca0f80b94b366c3ca21b7c2007d5a32a90ea4e1361fb9cf77fb1c450fb5a7638dfe7de9eba4a33ed57d229ec105891b1e9ffce7e5d5d773cf3a0e5feb8e65b356dd57bd540c9353eb8a7169fa6553f4d8e30a0c25ba17b23b06905a95366463a8a48663523ba6b883c8e3bf349e4dcf6721baf74e104190f2f9a847bb9da17742657553f833194802e2422f97d79f1eb303a139a9205331c49e0e6fcb9d45b94399f03019d47b7366644fb62051cf2ff17b6ea76e7407a27173bd5587bf5a44ed1103b8602d7d201686e2c23f31a16ca81ff89899d2068ade78cf1e0e849399eacae6e24f33bb39b2af6a3b04f74ff93165eec1643918f7024c562ede62c68a77cc8b2fd0c2ace827fb08bebc8e521ba0d075be2f8ce4ee606ad23d7e0111e18846f0669403df4801a7a512d54f21e194d35b653a6c3fdcc688480fda616af69d091a8fe78c4d69762514ea7b837c2557e3c695f7f618d46dc05896c4cecbcf3e891b62f285e7f8ceaa651b44a3ee967e496d8980d05d65a4a39b7cbab6ed36360549395c41bca61be93c0ab4ba9c2c56a28f9f1f994fef41ffa985b2d816a2cef0327b17df193c7fd4c38ad24e26483e96632839c1257194ed45aea56efb78326ed14d7dc21375e6ddf104df41d553abc02ad70856d1ceee3861d2cc39cbe2af85a4aa1370cf223712c389d778c484edcc28a67eb6a7663233c0fa668ba4c731444a65c0198a9de71d06e196d95ff4381611d1673086e47e0a2f5c914692c179fd1948605f607779ae9b378c3912b5f6c0617b01673948357b7f08004565f53e9a729;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h240f469cf18ad77c70dc5c251ef60caa11851aae24587fb27e8a7f568b873ca8793f6fb082367623cab7d51504b350208091496f1b91a1fc710ccf655b99cb39ce7b5130ad8e90d457e7fcf720bcec5617d6a719bd19f450544953a5d140dbc4415c364d0f207459f0a8f8deec6376a986868f3e6d343009f15d4a37c8c9e6850554df929856e54b3f629740e3864a3eabc52c58c943ec61e0b87ae2262282354c75cbbc85363157271978019380d3fb91901a36d4c034937ff08c3e095b5ed68ec039b27db4412171c0ae7fb8c2148b7529ab4f0976d5349d05e34983c7aa8880668da98ea0eefeac6c270f86c28992a71e6c7458bd9af8b24c5c0a7fac13f84682665d15c5d2968c0a4a75a1e9551d8893d6b6ba1574f2527f81515736ccf52c42ef026aad13af791949dca85bf7f89b692819091455661c34ee13204dbb00639b7e887a024f0d50a39b892e7c160f505fda19aa0d138777126463361a9206980c547c4536fa2b576832c3a98c28989d156024fe7ab69f67eb1e94ee89eedec10e54cdf426e0e790c413730d65492b359d49f302fbb51f8fde044c90a69ff58a5e0154f3b7e32463bd1c380d9d221030de408340944af94f7afbc74d099d0a3a49ca0b70a4206c46f3d536a8cff18f8ed346ff7735b77e452b446b3a431607446f79a88f918b9864f12e7d39bc5c857150779c34203381b1ba7313e3f9da72b73bd2d892bd141f55352f34ed77d6cef9253741e81d603e2871b73f13652ba2bea782ea106c4379905ee2b6d27899f144f4d724a1517e45a270e74b0cd0cb0d9f2c97fdd9e1eed3332473a8ac3d92e2f067825d3d910c8e0546e3a1fd5b9e59f4716f79973fe328ad77d870c38b769bcec914c471b4e0109b0eb5b48abf31635f05d541c3a1bde3166577512ba4dba47daad3e3416bfaec9677c3c5007e6cecc140fe03dc2db36acec7b3715a841c5bf262cf1ee613b8e9ea65ef97ac7b121cd189c99e9b0ffddd6f94d782ef5435b0cabfa4b13bc4baaee51034c1603cbdbd4c9017b064ffe3d87e2a150d9143c05e490333d2026916dfb2e34f05c24ebee28b726cf684008ff289010843803deae24fa527f2d6087cef5e1ff06252337695327115722667bef5651a1508278d2fa3e0ac5809c0ac88f9c267ac8177f1cb9e4612916a361924355f6c690d8f36f3c92d31cc7cf1f73023cf4f90a79be4e6c2320441727d0007c6e6a02e053c066d422a3f8baeec5f40ee25179f6dcc1bf165c0c79479992be4003912f12db67b0f43f8ae1fae48c784677fd5e283ed8f0c702314729abd5167727799742afe0382d7f10e3a56de657ef6d643e0bd6d6bb9388cc3ecafc0b29a843194509095fc59887804f7d8fe879003aff41fcbb26c4667a28d8470358eb2f1faa4487b44b227ba3e1fa2824c61d938bf7d3d3ce4dda041;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbda3956ed4cf172d8c259558f67a049b8dea6ef38d82c59d006c236b3914c82cad5fd10fa5b5f9d8116702f9c9bb9dc9adbe663f781363a628cad03959048d01384af04d871f75dc581a5e97f86bafb16b7d71e5c2fbe462bce0201cc4205e9c54c35f69bc28267d5b358f36d34fe8312355482ca4eb6ec2fa477349193017514ed2bfe0fcf10739a58b84185756df2a1c9dd19649071af4edb2aaacf73d6229a99447db95ddacd793f4139cd164b74f87ad339b694ce775abf49d3e7de6705723757779de74bf114bf9e6b52962b05731e56c39f9799ec3dc20c5740a2ba1d6bf5f9c92ca377d2f375762f4e52f136dd457cd185361553fee8089432aececcbd5005a5b94caa208d05c59d703ea8ddcd66a32b1053b9705b498027050f1cb8b08655cceae63fd586c200a404305b6c5ae162da6c9f2955d3fc90b06de566dd783fa1561309deef0b2912b0bec6a09746f7a6bc65c706f532c7046808eaee21f19e8e27606cc454202beda06a141c9db0b41ad42227d6e5d6956d2eaed23d064b9cafb8a12a3118b22b26ab9d19a9060437fcba5b8f88d2535186773bea9969b2b68ecba739f9bd6f69c58cc5fb5e297da3d2235d66756988bd32852e522c70081251ab4204482d5ee93ed40f6cfc8257518ce6ed710915bee9d450e4a4a29e213c02805ab45ce340afb875c3724c3d7642da7b15e487fdb9040321e7fed70a82f9098747ccf859c420116e2e628cd00b0674818fbf17ed1f4d1e2bd2f8f72f11423960b8350c4bd5f8446389c8dd8d03db9ba1c240a2c4751e8aeeadd27507f9f79ea5ea4d556bb0788d6111b0d5ea3bb490930fc7fd34fc19ed390cde7de108c5e66d01354fc52c8f1ba99ae381942009bdcf7d3b3206a123d8485a3d7f26b4ba3024fa794aa906ea3310d3c9551d233f60b36338ff6c5865658643300aa8cb9cf57422046af6c9ebc25427367522f8208e743eb471daba21646b1f27da3d74a1f3a40927b39df18743e9bb079394b8e9730d3d112b30760f363df6b212e3933da9b8e47d64ca10e45027fbf2fa5eec19eb84a874a8c41d537ca147d1191f1dc52f03eab46ef7ce67e7597117450dafa125bcd9247e14b97ac5cd827d005b3ebad2396c0de52422046198de920033e0e69c17e68f914b89644000b1399b0419cab5d0cbf71a72a8e520ec7a08f8e242c9cb8cc8ee3967623cc05a0bdc938949c80b9a2624b1ee54bf929e753d0d98582e8d4595626398b5e406520d5dfa7a084bd2533485e4fff73cea727f05b6e888e87e76439475ef7ada12079ea46ba455368d6823d7896e05d80f38176df52c6453bcd372b34a8d7aae9c0d5d5500064892c1a3d9117892fa57ab3fb9e6cb849bf0f3bc3b8578059133fae5c3dcd244e0ab961a64852b499ca8a49e31f54ca50f5c2734d953163e7efc161484535ccfc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h524d82829cf4d7c427db10c2ca966f7a55fd4f352017666303a9c87fdc21bd67f6fbd8552a0369470353a127f347a27cde0f2795350ed0c75070ec8c373069e8bf5f5fb49d0b356cf39517239164c94a0b51cb45792ef2c32877967174c3e908b8eed1d2ca336d79863341cb9eaa7f86ea35a7c6df2922d99a7b66a67099797418813f39581d1d29353bddd2cf7980b87cc6d8d4508495b8f2dd96100f2d1d5cce48190e1e94e57aece2c72f8e2ace5a6e843b19671e12513c94bb4fa8a1654133e70716e68e493a28044c9492eee46ef94a97331d3ae1be85a7a79f3af0b486ded0a3dda057c69275947725f5b2fc34a3fe4a1e37c3ec8dfaeeab127f093f84c3acf12e3e82bb11f762376805cc8a38ed55d7d35e9417b0bab2a829f66f7ab45a634e1628501bc9b270d5fca7ae26ce8b5871a66f87a5055cba4e44be9e862bd2dc7a9e73398f1674ebd34b7a12918c4b7e8b5a47f107618cc5b90b5b2e32ed20503ac3ebb1ba785c5daf1fd8bd57f63385e9fd2c352f93c5cedd48f9c481daa2542dbcb37f6bf55b7d370c037c3a2aee6d199d17b705f8d84701c40ccf7a6b8b14a0226d98e4912780431e021108d5d6321cbb5c2f0fdff2a6dd9ebea5b0e77100fa53ba41dfea2f087762922c4ba9bb1592fce68dffe37defaa10053a143d45a7c02238d44c85e8cdbfa126b06781f4a55805b0cc02f9a33c565c1526e369985c4c3c9f1a00161bbdc16d0c4e02078fd3349512cb5bf031e1c9a392145651730dc6f969952dcd2ebbc2232df07f9dafc21a1f63833c088516f03a51f829788f9118109c8e964dbf196dd525bf0456247ae5aee3f5c07e5708679e50ebc687a33d28bb5a2668e0a23f8c3f421e3a2a46d40ff9446b8b2f72ba05ffba09731a01487d99181efc2a72f6cdeb53946ac896b8aebba81a4e3fb2cf5e6cdbfca71c54ec70a13b8ad06f0af6f73dbeed1e4cc285382b8b081aca55ae5ab41abb3f57ba7e383d9301397053ff8a72b00e3d5139b194e55ec6cdd3a30641ba06908437d07b4518863f1aa4be3666ae34f8303e557d11b484453c15bc462f82f9768f97b6446388cecc651bcba179e9ee8fc388ae95dd2b5b3c3f0a00d89db086bc735409eb5dfe7b58cd7d1acd6e47e3227eff608000f489f1e6b7b782ff7db659431cdd1073978e4278ec47472c8b616e9f73e8dc5f28bbb5faa76a4b10c460379a37b491b6b35a739f35d68c3aeb8f8c9adaff37c2817c9c8e5c5427bda8e58261c41aa1de94c1777f7d2597b900fb20b0b7097877a275ea0623383160966bbc6fc796a6890adcdeaa357a8056aaafb8c2d5c081447edb9d1e9f0f8e25d7637f14bef56e0b3fbc59133a852dd5c281f29a5279515e849d68dcda0f9181b565acb1eb10a249dc201a266397c4c00499e658cc9de61b9444484f612103f60df1c40f42;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h36d548f95c4959b9c6b0b0bc8185704b9269e99b344e845b6012c9b345d9886c97a3996c57bd74994c05c549077f39fabcc4578be5ffb0eda504e826f737a471627daa46df4c24c556c896dfec6fc6652933fecb5cb0d1d61a2577e5fd10da1c3fa93f29440d824e5ad209bda0641b8698f31b5a923e365542caf0d366446f5169d0b5eb17ebf424c2bb94ffa6361462943fe694f3b181badbf8b26c17d78d433dd24caff05d8e8125c942d9724f677d078984f1944b8c2443e59db56c4f265c362a58c65e123a1235ead96d881e4f1ce81f4fd826a6b4ca56448d8ac5bfe8f6bb906f79ef3703597694c2c895df35f57ee5717f23e6759d874a57793701354e0ecbc95a787242297cda477719f7d70ebce5ae3737fbfbe3ec61ee6ef2120a6056040fbe4fa11b094930b4cc7dc0d61333e0c338c1f28662e8c3dd8d87fa3c31c26f6407cdd3784d285abc24ee7c233358026e298a5dbea93b8c644096495cb8827bdcb3422a818bd7d2b5bf6f020b43dd0cae900b974f6deee46e0e25b765ae3efa76846492e4227ad021a1f5855cae16caaf85f807ce0e3f4a70d60c5e13ff92d076b33089a427ffc59ef2f295ed807742fa41dfebb2f368859bb9da82128069a517d0cf16a99590cbb45545aa80f96dd702f27ac9c7374f90adfca5635aee151f3c9ce973ba4d893bb23872229873c5ba2943111cd1dcc92a39d2c94ca705c48b457cacf40876c05691c26df1cf9b0db96fc71df93a3450e378fff7974812ee08b75aadd727e4c95c36f7e663d0c8e1915e1cae62f9368ab1e33dfeb811c3e2e0ef8d8d7d1868810eebab86a50df834808f0dff9fcfd2c602110b7fe7e84b45fbdf022ab576d2f7d280eb7a958f0bfb5ea57bee4b0a2ceb141a7beadaf4e02fb7080a2aaa9c324024277b6bc72bd58b357fc14283a726b105437c1170a8c1e7c1980b7e9c1604290c407e8ebbc0c5c36323637e545d1b035fb110db016d361d0ac29749b18ebe6153829d2d53c1054bf91e0188a211f30685bcd0ef1069024b62e8359f8e1b5f433ecbac5d6a50b84092ed6578564f0032bd9847962515a045e71ecfa50bca374718a3b2078a3ed262e567e740a26aa4b7753080ad0de453c2c4ea3ad6f617be5c37fd832dc21f4d879481ab580bc999bc4f3abbcb8273c1e38cc8777e880812043c72c32146f0faa3f22739cbbcd006e5b901134b1f3bd6082c40a833bda114109bbbaa22f7e06c5a04b5d214bca42e933370d1dab5223b8d77fffde5da5745e16f2a93746e899760c42f005c042c7caca72e74b0c7401bb519a33520b846d20c6dbb956766f2d2d556367e5cae80db8bb011f380e866fb485a21f5d77e437e187f6c7e75cc7e877abad276f3efa9b6b52428b65097243577f840b59eeed95ba8a35d300158b9c3cc770fd4895c101eb21a6311da7b418c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h55f3eb3b59db497f7ab07e7970968e39495e94dec62f2410b0f54af60fa8c77f2a30fea4091213d6bd912604397a03bba4a1568c456fa2deee435e8cc6c5ac7d188a7fb865a7d9280d22665186946a99943769d4c8d36a8dcec27eef60f650c40269ee622513804408e1b51c2a897deaca19dc152dcb1ae14e8aa19754decfe2da56c8b8437c80c3c7d6a3f704b9689c4cb4c3ad308ec5b9a2ea7ee2e499d741e7a513203bee1af03fb34601bb643a715995d0768723936524467297672514f99bd5908bfaacbb3d12193acdac6e83c40d892658d70138facb68144f6a6ea91cebcceeef91616e21e4dac1280024449ee503626e98b74a2de95485b8e7db6cedb1a24174db81ac695753c3ba297e94d8e54e5f197ba35858ca192d744418bbdd42502e8e520a271136858ebb2a388ff22f2073d14596607b955c2e9b025362fe41c30be5af46970a72744127c0155b636702828f55650900d735a085cca30432d3be7b694e7ff917b5c7760a2c2f6de4f321be3fd6d75108950834389105411e1fe57854c3a38d95073cc24d9307e47501dfa5bf607fe4d6a88ceec1178a5a4c0a925e81d52a6c82c3173298d46ade46a37843f7792981682c9f6f677b6c2f0dc4f7663be47228e96f6066a36ba5b28079ad9b583fac42fa339c8a3537b3db13ad2e07a5fd7cbc11d2c2dff76099de76f06967ac76328083d34055b7558f47ca6a8f78c3b9c751a44570d052ebae1d9f3f6de7c986d0cb588aca2422120d38ee76ec743181fed17b5b8685303e15d176bd1380aedaeae869ffe1005b00469d77813e7698c7806e156e617746fa30b765a0359fdf695e28276ca618d3d5421dcafd7cc9adb17ec69a081f82db292951ec1833e4b81c83776c8b88fdeccf7d5bce148003163c120db267a9edcfa1c6ddd234b6fe4c9c430963fd2446d0c8b56be017b4f850d893001a88e20ad2e75db9b390c9a1864ffb44e8ceaba1eb848f19acb2078e1caf7cd872089a87aeac856393b6cc4e12601b87bfcf47a2d99cc923f23c885525b02ee1f6c98044657bb6f92092b15f4d3ab1b963175d65c04fea54208ef681f735120b73471892a2d3abfd7ba2034426c1ce2ce183554bcb8e4183bd8e711cc8c195d3497e4668149aece09bed49227718f8929916bccae3c97ae756ba4cbc55800dc628acf96670247f80b5d64bdbae6c0693936ff172b8eb980949d9d38642ac984268c5065b626779ead06af034ff5b94fdac58f7412f09a8331d2d5c47bb59c31290f334fce961535f7927fa9ee5701637be2ced1ba7099df59ada8935693f26c35a1d1c318e024607994515a2a22947a0015fde573ea9e75885905d31db2718728c868647fb39098574c0d01eb51c01190979679df99199da1e5cd2198543ffcd63db8f8deae6d6286c7c28f56ebe51419378ee5da7bc7ce711;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfb39567036c6fb6894d5c296360161493d4a65ebeeba16c8aa4403f1b2e55f4486d159656d44e91ac52ffd7c4737372e0de00bdb4fe6bbcf55cf3a858cdc24dda8582461c052af6ca8774c9203c972cedf992ba58c324333ab681576b7ee9b692f1b6db0fc0c96721b3c3c1ea82638d191d6b3c6e7f60b4e129ca9c7813c4fbce33c91fe6cc4e290cfd399472684bcfe20df3eaaf7857efc4d54f81ef6cedf7867c0f8d1fa86c53334aa0e61a88442a3387edfac8396443ce08b4dfb22eb63f550e47a8e512ee1fcda047b91a092d93431f550183afa5658d3771e45eeda470d1df258f2f4d2b68eb26632f6ce3e4677e6f8f1cec013398d2c50276dfda3a6260dae90d680081f6a51b81f79652b1425f8448d8ee3be63eff748bc781f52b66d9e82998806b915d8e8026e83f04b431ba611caf7c55acf83cab8804e0709929142b4a4f826021cc12c8dab140eac9887105715a426a8a2d75f32ba2351ee263e102046152b0db22b2328daf16168007b8c8f39a401b32fef1e4c2b0f25680c19bef1b99d98643bc6e4fe6a434ac55911e2cc18c7e8524287877c5c03ff8a73ac7e3e74ff64e22a013c9b17e9b0c334a3930079a1510e82e4abe53436cf024e8aa8f46ffe5caa1f424bc1dde4bcdd12b5d941deed6fe7d2bd5d0039ceb81f6b7a8656802ebacc8278fb24165b162f55721304f9430684d1abe82304efc62acdea8e95195e343726d33da026757cafd3b99268d679bfc76d6d963f92f331b13f6eee231c1d9bdbd7a9273e6b02d94ae1e6aec98e889bd2d7cb0cd532e3732694d30d4ea114f11177cacdc40d2eb078c7ce20fc0a107b572c10fda600643aecea66701973eda6a0a2489daf0974f075f9c1ef697b39075338c7165adf8126ae00029e9fa192749b0097b560c3d9a9ac8c22cafc3a05c285a247d404b44c255d1e0b9cff2b9d8d83bdda36f61a729b15ce33a0e8ee17f14bce2c5abaf83cef08adafb969461abb63a1d6684b3bf8b54041ba15e3fa03f3679c9eea105f47c0b91ffaa0fee2c7f4790284cad24a6691dcaa6faaf7b1c9729c59af8f24825965f920f66deb0d69329344414a7c035822228e5c19d1f03b8d4b661d312070da70c1c6cae279af6da609f275d0cf91a0cba1f5b8968c42504ff5051df268f8d786703bb405859c4cd02e87e06e3a0664e76bb5d9bf83c9285f1d7e6b7a0ab88c9070ef4f3d92650d63bde92ffcd6674e5545eed47dd4b71e9cec6e1c345fb62ec9a36eb870f16f41319276253c5fc16eda500c727311483dce16b94d493c41cc9f41cd9a05dbbb2458acd33fd3d83c1bad09115bd741653b952b1fc2c45b380277a8d02739fb7762bdb7f7b3bf183d3ef5ba1c5ecbb3e4e70008c799671ec2cb33c5fa18b564b928bd3a5e58242e4f1084efde727dd5914cd521a8efd6ada67f020f7bfb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc96cccbe447140d3b81ed1a42a0afabc048f561718fdbe6dc1f54fa8915c00ece9ce7c688173557b3367591d7df9dae545f4ef4c607a0ab77908b3fd28717c6bd388bdc0b0473e50455dcea7a8b3e8145dc826f8c917a14aca5f4a67d5230f06b5736427b2cbd83f4248293daa1ea8c0bbbd43b83b120eb9967046a5511c25e27f6cde9c0e1bbc40343dfc1e9390064db465b6657be513349ba95027c069921cd462aa6aa2a625f0d1c9e2450cbdb8e8c8e9fed0b76615c07658df1d9fae461752908bee417dbbeb1fa0978a83c3b284dc46316666c4f96a11f6f77462f59ff5ac5526709e86abcdb40520b028e9802c1bc43743fddad9ebc0a3865aa09df84d9b6f54628ba12bc92476559c8ad1843473f8e3c8a587f86059cba93f7385d768cb4c8d33f066bea154b803cb6b73f51f1eee957798bb7bb238f64384b732e53f6355ab531d451f1b71fcd5b550d40e4b8627ecac161e819f6ca3fda5f58a58c643e6b97f773b1d6481369653b54238b085b160369a68e9573327c9b8d2dcd685b430c01d682a031f61fffd69ef2500718f82c4a5d2adc22ca5a79ccce5b68087543f89a9c222190a5736e15fedcb2b6936f2c53b8fd37496d3268f1969b7c269940d5aa33f8aeb33a7c71572751e62b044a973f47f25bfe1f9b9e89074b148ccb31a6ff07c7033860fffd9c80b56e4dc15e01e97f4d72d63b89667d726aa36a2ef1dafb749909b6c198973dc8d5f16a4ab1b3ec5e740ad4a6ebdab95c033e6fda1c16a8606e11c00ca0053129f53fec7f89fd5670dca8ce8607c5027d705a770b0297415036cb390f8b72cd4fd76022f4e8d26874eef4c4bf933baddc222d04d639ca63887dcbf032199830881459751e00374f3c8c8775241c823708121542406d3fe7bcd0eb21a744bcd36c9211a7b7094f314205d3e3c69a1be781311484cd80433a96b956d4d1df824623217c586e17017bf3e9ad6758f88c67ed145947b1f011f5ffaeecc2b3593ae584fa7590623b1b4fef7e04162fa8dcd80cf9a605f026ab38c09f4c7ec8f1789436074effd0a3588f7ab89098e91628a92291135a1b051d01533bc7ab018ab879a2f8e86d4f51caffc57c9f0ac91a1872f9e73f8899b76ef0f2e4cfc31b7ee2895d3220bfc17f651281121de10c1fb21b1bc0c8786948635951b1e09640442f8dd234e66d9b6c9eeb685e416e03c39e20860056918043a8f30d236e084b28d44aefe49ee7eb24a968f76107905d0c5a72fc8aa657185e228f33c3cf4d402d35754752d24f83066b801e2a4a8fe12b2044b8ecfc13e49bd8b9b829a88d3d33ec9984460d8f5b954ac5b44520b310a3f9b9646c808ee0fe7c2a86e2afdde984394e5db454d5bcccb63aad3165c6827d3b795112ced989aa9dc3570e8099b1e4d2040b1ca2302609da44c4f9c13d365780b047f10452b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h741e2342dc82bffac5b40f6493d71f71769982fbf28f860304cbff291f0f477d2bf1c106348506328f6efb554257888ccb04fd66be867f161d5be86ae7536c26c94c84a1c996f40320f91b47bfed1ecc1fe5785a932d2f5252266ac74eae3230324d2f36fd4f240b3d374ad043eeb2fe19129a0dc4520ba912873e608a8a40d5929054220d7c03eacbbe32d056219e8f60221d1349e34f3731096aee83271d96050dcf7cb09b0b739a5bf2e4d81149f4fd90ab8b13fd39eb0d9445b24ca5157f709b59372399187667c9c4ae3a07518b9a3a10e2bbd61958ac8231d8b4635c5fec19d67bc5c74ecef2168a68ef9c28cf9dc6e9e8190ca97ec1e7e50a77261334de97fdc37c8e059b2a46628cf176abbdddc16d833b3a0c384b462d324567c023263c8eae15f0e4dcf9de401664416222ea0de2b9d4904d70c8e090b22295b4974f2a44c0af19ff8fdbb1a8d9aefee2a1828b160ee64c468ce943a65193ca0067e1fb0aa7d18a87c97cc9862fd9e852370ac3abbc98a8949ed96ecc317b56b16f06ae535ca70c047db2d5b95f4c54851eaaa0d828b328fd3311bf3c62b2cee0f713679ae000684811d3b24d48dd47b4adff074e6caacaaafbd99e30701ed56134603ccdf32f701215a93de39ff90fa66c253e898ecead7a69254ada76ed2609253c532c085b283785c015207a2eaf74bbbe62de1dd98b07d82abd461d63428b2b3352be7693ec3e37358849ed8d771abba0f3a67bbfb9249820525e728253301fc0351b5223d187d16d49a3d1c143ef8bb1be5154ea050013eda30ffe9a91123d5abf0b70fcf61ba66135b44157ae854ed7ab885e24c93ec6c9874d9d0175c89cd4dc25e29d70cd2512bc426ec4be9788a2b4fd27e6e88ac10ffdd32491e889258c3442ca9b3fdb864e68378e76f61ea0487b08792fe58391fbbfc6ededd9b4bbc774ace8bd7172d31c39cae2c85ad86e0ad505e94485a77084d42e757a653331c71df8bf7209855644ed8d04e34865b3e4d5857467dfb81855d5c117318a8968687924ebf61224d1b6117bd7106d34dd567f952ff2393fe18dc1ec9017510a2cc69569618b35ed6267618298c7e68dfc3d86715c5730f0dc20b11886cacdda4c01885bdd5a71d231ea44a8e3c13c849ef502a543138570ef4fac88412f3c58f1ee723643365f84835cdfb365133802606853c72f66c704fdf682d23f0226e14c675b0ec8dfa4e07883b94e000673740a15c791b4432ae290e12404e9c1ef6f5a5b440864321af1f01f873298634951f4137bca86404403635ed070d84286a849082ae24c589771cd7eec73b3761a72bd9218dbc2c8e3c13463703df8ebff062162e952fbfafc9ef8beb2c2aa33e5d1c0f8d53274e3fd8db22f57024b23cb538184b440e1a94866917fb64d9a4e691c59451ab2c894303a96729347e73c3e47e5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h51e0bf02456d61c39a387932d610773becf957f906fb0a971a2be450b45a52271569e4acb48cb5687b0f791f56786490127e18db9a3a61bb7a00bc534ff0a6fa0bbeb79f43600c1cf35de675c33a6ed49eef154c257c77af5cc890d07f43b0800b70d1b682849907e720b1cf64f8c6645060dc326d8359e00dfc2d3af409b9bfedb56c66e5544aacfc05e9d32c81296b3130639fea1b5bf185448a9a072e67a0fbff7cc8ab2b798bd5bf1c0e92f4623b5805b2b2ec0cdc5d65fb5435ce5463c0e42ff1f42f3d337cdc70e5f7494ca4de8d2fd2cc70a4480e8be56dc01b3d6b51f55d135adbd4afd1a0c825b3fc0d543ac88b1d250ebbd73215783f3c19acae8565603830257c224debeea9d1360b7b79919bc650c7a584bcb38bc33420cd931a32a7525fec1dc3c0cd00ef28e92da2503301975ccb5c474362911cb9a931403c47186fbe96fb81c3bf0442e7e29b698b28edb98a9cc271de2959d077c559385bcb00968fea8be30e33c0050b64caa066bec51b2984487d2538ab78f7c5e0b00eff32cf01f6f1a13200dbb98db9dc8cddc46a206ebdfe383390c6a569df3888f523cdc16f0a16f6b344e9268318c1ebc356946bb8d6c56b70e6b270cfc4e909888eed109c3894d0557418ca87112a56bde2b2aa371b7afcea0eb062cbc8c4dcae90ab10555428be9f1fc881292c6f05d78cb0700a216ce2d2193ebcb043b94b3faaeb8a72ea921680aa6e024fb06f44e340d782c3071bea81a241dc33d535c856d1b0c87f17a8d6e297ca5cfe368adb5c0822feed00dd895d74017c64288edb15fcd1d42a5e75fae2b22e0a885202f5c4cf43d7c6f9a2237d34a3d6f93e15ffda265bdeccad54a17e192f41b226edfefe7b823c9772cfe6daae9706f615568e9f6feeef7f6dddb0d1ab8efdac286a4c1e167a4110ea263992b4af3894ccb4529438e70485c66a56b5e283aa94cdbe0be12bf691e9d8ee9bf972f7012b4a27c32247ee7cae4b909e0cc8f90b1c4e582def460d260109e43152ebeef756c2a4ef81e4e946b277b566cdb8551e42c6f30576b4eff07721870dd0b0f4ab1891428d7a393453be3242c1d1ff1b9bc748ce3c8e04f2e90fadd732aca056d4cb1e6f0b1afe262db583d2e8e20938fa703a220d5c0c3af24d6a07e914c76ab2b38c210b27cc47565c449156a989b23773d1f08b5b6a6262001e93621e1d134219c0b8a4cdd8aca89d04f12803b51eeb59b5a97af3ff2acb891f6f48191f499d5f07189d7fbae79737f0051e63b5512cca92b0c8f27d074f18600a410e4c75a3df195121f081f0f67e77ffb1760d46ddf15ffac075a0c4bc396f7e954eca1231118b4060f201cfd8e8b98ca9d88425afb3cc9299644951033a6b0df875fccc5dbc75fd310c398af6f9e542ba716cb804965973ab0c3c4cbaeaf118398ce8e563b32542e452;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h295d9bcdc44b433724db42a64f4b49b4221c5b9fe888a9c5a5600256170d3bce0b1e49c92448150291dccf80a83f8dbf8dc035e65fb2b6f3caa5b271aee28438b7bd9149cb42298ebf75bc020f4681ff77e318d83695f7beab4c66d5a450ca95f7d7801345d97a6a21506edb52dc7f53b658852a21c9840849970232207c2ada3744eba4c2a31895fc95cdeeaadc2ff894230416737c61a1e93f9aaba2c60320095e8371951496b54ad6fad181eeaf2dce010d6649969443f020d3eb8ae5e1717555e28aa40f5efd5cfbd3ef821f3f54e4f5303b7eed72a88696960107fdd9e32ff05fcfbb42d8424c8f4daf0291b4b76137d90fd21e2fcc0f263dfee0a44837e1ecd488d2e14153ddaf7325cc3c3f8dc75723f48eb873531bcec77db5ec4513fc0e4a1c8bf943802728af7cdd1f5223b7651978778707142d606a444396c40e76aae27f0a31feb85426ca3b59cddf36d7bb0189d7a7c5d7328288a61e908cdef16c075207b21f49fab2f814509775ef11c6004c4d7d3b4192fa4bfedc0f70d03c7d27b2e2876b0ff250babd9a7bc0e45c0b795ee5d1b1bd54d5b45d044daec081e823b406247ed4d7838fde35a363ba2c5720802c86efa638c4af02ed069157896522d20a3b65f3d00f952b334f5827bf34039e92911e1c9bff6fa36f883162d639bc05562413228e147369d6ac083f88d74a55f18c8b113ef9a42ef0515b71b58cf9178cf20f4d48f57defb91f7922fac9de0903055db0a38eb6ea10f99321852ebd14120add77d4204f258a21e8e66964659b9a60df98c2bbd4a8df570cab8a7e9e5313a18b7e7547933f586b408ee9ac078eec3e64507bf7fe4cbe698176b6e0eae9dfb19f110062a802a8fb119eb75fc36389e9b6d61a998999e92d6bc417c565b30484ebd84dafd3c44dd98da0549117ec0130d83b5f193a4411aee08b24bf146d64949de756e7935f4905fe4dc879c1c413787219c2434edc9a94b97e5e6c9c99ba633293cc348ea9fe3cf89e0f345ad3b624c881ece60dcae341d2e76c89521c42c273dd6a87db4fd0ad2a99dece5f40d6d6cc7d7d1c23d95fab187fe7b888f03e65a899777d29d4285a842c5fceb71020f18474a9e00ee0126da59346f55514f0477d277aca62084f068bfd229ecc9b3d2f959dab4dd4fd8264fffb98a3c8dbd320c75607478c4d35855b315b77fdf1381951b5e132582a15fa6973795b3578c6923c59a14d31f7bbca744da1b7cf68507b4f5bd275c747dea38094e6445f1fcc8604a1ff096f716380f91e93cea554c8161fdcedc7a3a0df86385dd410360bda1cf85e9e1249a9c62aaee5aac3c37ba7cec232330caab43992acdc0f7ac27799fb8867f1d57f3edc1baab4d87aa7991f87544a1e3ff47089b1ce636b28c356779b61dad34df4f839dbbee267b6950b99061d029199afedae14f8a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd7634fbbdd730465fc669847cdb55ca0035ba70b0043e71b7085391ed487073b1fc8adab53a458ba47708eb88a6a141c28cf063188726da22178644a6277adbdc5f0758a7a9e5b7f0fb5fce1a5899063291b83f8c2be55cad4c7fa3f0ddcc34ba9eba68a849aeb64a2e69089397af358b603e7eaeca364995feff957a3a1782052f612204d49f608276c8497c962a813f0b04108824ba018fc740b7852d1636df775fbbf06e949c6b30b368b6e8286654d8280a9002be4c22b47e747d9300b2c7aac6ffd26faffc94f1d6bf4237c2a6b06999b7344e7225033ee3cd5940bca5c4abda805a4011c3703ed092f50f88980f97ebe5db67f20a782e188176a7d5bae14c75aea34d220bf9e9869593e23fbc0dc21d15bb539b22feaf9a0f105908df2ea3000461f88caef62e3d980b6d726db597992e73da2e424940c12f58f0133543164a6e03a9ca887139385adea637ba269d956415f1007b644a69d986efe1de8afb6c196f2d60cf5b6890683dabb566246dc7c06c1031f691b5998c696492a961f876062d6c45afe52e9ab91f9df0855d0e3ab25924076d204cb3144c965f9b80b70c2039f1de6ee26e5a654ae314a70cbd5df81badd516b89b10f4f4a2a5351f987409ef1ff02e70b0ae042cdfb50a3cbee4098c9dab5618b129d7fc277f465fedca00ca1b9536effae90c7b47f72c757558887b026d8c23540af8b85eb8e29c1e01633a4ca216ce2bfd30f53392dffb2a45fd441675745e0dea011c985f65199ab641f04a397fd357c91870e9d97e08c4881843fb87983ffe761c8cd09fc280c79a53ef132af317de6fb330ab3af08f1e229ec429d45fe5597192929258a6ba3c8246acfd3a11741d34614c7d3576868795f736afc9021e8466b37601598e7e32fb4ff364bcbd6c5711a5b785943c09fd4a61c63250aaa4d8a9067f324b2868376ffb42b39f5955c8a7e2e69b60e5a8a5044dd36a7ad4b002c4bb7cee23607ac8a6b0d827d750ee29d1fa30a32c4d77f25ac3498a7790d12de92d169735714dfe2fe562621ec59e2e05b13b8931e964bb30896fde039e1246d729c817923dff36da0dc37c1e230efa71caa4ae0396813faa6a55631d5a0cdba05fca196eeee20d3db7ef721eddff0f6424146f6ee67c0ed722381ae3b1137331b662657dd1f1fe04e88e0ad4023faee9878f4c36908f5f955a698c6c2b2ce916f0e5a25530ab84857b2abc201f765b0ccf97d5386eea09f3d22673545186e66c92248481c503c77cb6710371b301f74bd9229dd9cb5b1c73fa3f0c9d7e0accce6a22d651bca473b560541453707bc2c4443995072491c1b61deff9b977c68fb4d2b681088f86a0bc2446589e15ce4ef418858798ce24827bc48a2173ea989de4bddb482b88a5ca407cbcfc327e71404487463116f3b3c941e5a391b2bf25aeec97f9a9473ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc316ae50192555f4c3eb497d010196fb594e0be4ca3640b3edbc52abd736e7ceb1dad9a1437a7d76ab106124f891c61904ff92ab42b46d40e142e50c34c5b9c3efb037cb787696b2ed1c99db1f0fc073360f0fb4f7ab420883b366b4639665594a97e15bbc2f4b1d9879fe4b78ea88dd0e46e33ea0318760e540cbd95bbf4479e277df1b93993707e0ae820f74685434aa650218261a8cbcaa2c1952eb4eee24a6a1dd9b3dea87268d703270712d934b594c9ffdb153df2403c381e6e734cbe2dc93f1451ed0d6c34ea96241941f67096a67ff0d8af1961ba3acfb59df0e8995a8f4df17b30d8e34daba0de30ec4db8a350b6b1d6c3ef708e00d795ee0886ccd655089ce780e808f68ff4b710af041a2f1e0f00ebc86b2c09b99335e5e96f270bf45d624e0bc309749bcf379a149be64506b2df70b5fc42754a72071eb4f7ccaa9680caeda6a942d6e76ddff6d87b2165521d0cd2f5daafa2c055d9468601a2b8dd2f51eb39fdacbefbce2adecb8dc57cfd9e568fecd9e299bdf58062e1ed103865b6bae41dd183f905d3a04561e40b55e6b7c5ebf7d3f0c08392820a07d84df48fc538d92d2a3c2be3da67d89173ca1c40a8cea335e70392287e2ac2bb8487178178ba91ec1989d837acae33277836d362416a2a8b86f79b2ba1bf07ca0b9f0a23f75b5d353cc67a24640f72b32999c6cfd67ae26509fbe608ce8396e1bda0a0e6ebbf600aa4665270276f73f9debcfb69f1c3b68e882df67d8fcafe3d645f68d027132118532e600ab179467fb8754a39236841ddff8bf69c8c82564e00721b681415f72014f2003e6a625950d4d937bcfcc8162fd8f6e714bb0393c5a1835e090b9b57ff35595c1c69877b6046a6bda5f12ced034d1447280ac2f2bd53d07722774d124e37aca6fc7979631cff56d7e528da2b7770c228306ffcd5c30c328428418c228ba26a170478ef352de7a412de24370de11b8d5a40c9985c300d3c6dd4f9cd93f03553201d64ac2b0a519db515e8ec1ee06d4bb6eb929cd0be900d5aa1719c94be436eb2852d8127702b6d216d52218181873a4ce5039a23b53cb9bbf8f642996cfd3efcf2b4cbe7ee766c61fcba48c12473b6e04417082e8a4d6c191b7fa00fedae1d6f97bf2449aa39c9e886ffea41f51edc861bdc328a399131b03639c1e28e3d875411d21cf768784d069aa90b8bbbed4c02ace9efa96264f9a591ee035b1438d2be996710828a807b1765b554b2d6944de26de2f9249b9531b27c03d6a24cb9442a232e34373ec10618025808bc8c49c71a4ff76da0cb5a3ea2a4debdd46e1d7a4d263fd8b0a1561be269fca466d58c40c52360b5b5642149093fdde85e65af6fff775a7961c03a823a767318329c411d7931b34bfb819ecf0f1d313ab1788416e2b49fdd2b7acbfdc4d0d040d8967ba974723be68b277b2f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf48d9ed8588c8e5187b761ba3a4e2f25e87ccaf413f13fc355be0695e0f4c496b9eb46cfca088e7855f3ad3f16d6b6cbf3f738500fb93d47147ac4f37b504cb1560f54a797531b29a45efa85b373ab30c2c0633b24754035ed44aacc803c9025d08d007d10c853f47497894519c7a4bd0f4360298f64680d58a0a424e89a5a08aa2826102421c179d2f9574f0e94980d3f2f9d8bf6c84126591075d589f5e3aeda3c8a713532a6ae40f27ecbbd9ade51f0918fd50e89f587f8e9a8879cb1037be35bd98e4800d0232e3db4ecb3b52fdcd367a151a7be7593ba4d3bdc82301b30c9a95ee3d0b0793950c553419c99a4c4839f521662afce2c30b67d27d080d08e3d19cb65df75e7305dfeaf0f6c401ef39f77fc218b2a08331b7c75aa75a91aba276fbc8ae66ac7ca6459686511a91e4717dd5c5e8904ccd2cd52e00eafb657d8ff3997594c637a3258f8e46a76cf9460400ed6b84fcf8debf80f96d8809e1a3d9463716f8cfb92a631ea3bea648e3d0c1f3165e8affad9f66a9398ea46b1f3c353f1562553b4d12ab9cd339c85fc0da0991b88b7965c04f8dadaa4b93437741ec35b1b0b5f2946c0271a3fb1eed8027c4dec18f7c010f9715347203b9dc828512964e88f975d91a8139f8d4fa9069cf2ffeeecc8ac510d60648c3cfc6baf0dd8915866ac85fc57a6a27cb0e392ac261413a8791352bbaf6778a0c30640d99c04acd116aa4b848dd3a974c361d636a70d193746502aa67f98c763c8578816aa4b16076f772c482d4e2edc9657678cb25fb9f2ab931628f77f8f703a4ffc30fc885bb0ec661b0633c8c75153284c7e7e1bc0804d13d7a5cb702e405594b7b6dbf3b82ff2b25b61d7229c2f608e5b02e124eeb3caff877769596ddde31b8d2a8271094c4e214df2415a41b62d9f78f845be68dd6149d90fd5f0edc95b59b57b0666335eef7c10a203c5da2bd54b67f9b8cc0b165e673761922b9000b4b6285a714e46d5a55e2fcbfc7fdd83e07913372bdf77abbe6bcdad1485a2b5d3ca3e1462cc60859a0247bd3f6381f127c4f2c88b43997c2dc113b1d64dac7525a3e1e90b0174c613564d207b31674aa4d02ab277002d2d7a9505f75712811ef756b6c81fdc2b7a686bad9278125a9ee9cc375635ab5d479141d85d1a334611bc67bcba8b06dbbd8eec4855ab20a1f0168f06a61b74e8358d83de9df0566e10e3ba61ff820469ead8e3057bd9d6b311749a0cbd1ecd74f385f89efd76812ca5fc1d5f4dd5410c4e34343aef57c4235283fc00567150d46c792fd31e501f4c434439adb8a81a2274beb51e847aea5abc8f516b65f04eb490dff146281bec0880860ac188c456d841250a6947c614d710dda9aad8fd4ef9617c288a4da58e9960118ba3cbbcd7083b197daeb24025db51ae792bfa6b92420841a815291a228192b7115ce8ee40;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h841e92cb3c4e9c9e6a3de109991d7347bd642593461f4051c5bc8f0596f4a2dc83ba8d75e8f2903349051113d7efffb879148de994a2c2dde8cf540e87b3aeeb35fe5a8836fa3b185adeaecc81a00c47c98857d7669e14abe831e194dc564a300b2f60d33b09f246d8d7d9494aa2da7348bf89cb70482258674758df909ce38dbe9ecd770186de45ebcfdedbe38b792923abfad7d390467d0242d673f112538ca31f888cefd6022f7dd839dc23171781bf100b3a2e9299e9ae90748244ddfcd6183be30b4a60b3fa61db02f4463db912730ff9a97cbd292cc6cdae261eefe911acb7767592372cc520910d45d9c8daa9725c22458b7c18d2ea59cb1290fcac60b68dddf3a2826fc3998cc99abc290e1aab8443ad18efbc47d9afd8f60df6608f5ca39b81c920b17f12de88baf0f645cbb0255dc9ea2c8e0d3850ac8d2a0011beb2bdc2d5b1e0c39bf3a1ae1f644d0afad0449d1bca20d70ff3c6729c08548fac2757a75992c01905e92a8450053b713a38ce59325b6e73259d2f9b9c9d25730fcc5009d7b5cce0a93148abcaeec5289b14870fd5996595579a95fcd61be9ac1cb792f118fc0c9be408a2c802086c3a57dd475af50eab46b65bc94e236b0517902d2f833034814927f14fca879024c114c7d3010b261b762610fd582a9932608883f47dcbf209a0f291a8f94c1205ad2b2075f4422dfdaff05f20d87614045602dc17d9c9bf1551cea185d058f6edc84c55b55abea2b46a97ce93830ef411214bfec732b854cc6a78fcc2a298049f12a00bb5a363d746d55fb48f5e03db48a7f2c774cef081c324406f4a40aa17d3fe169394f269617ca28a6db340b739240b4a2ef986e2bd48e5231bf8b1bcf55d758ede0d355ccba87903856000b1bb010aee1349aa2f1ed58e3dcedee0f374a703c63d838109c989e6f8ee846f5652f9f4d5feb6929e32c9621020e363552175705260bd570c122abec9c9d9183ae04979fe9fa86316b4b7fe80ff9675876100db277bfd98f41313eba16e11825a9c4447c0b73962da56d2e5602282c95d24c30ef4587f4f78fe218fa1831320aa004551433525c1a55786dbf49463a180749bcffc704a6890aadac7568c3ccee5fa22a0cda1322f473b2937cc442ac098fa489c3a70a785c0ba63c6f1cc13ad537bfaea6084d59e0793faa6a24b172e659f13d0cb00282fd027439c7cb3fdac25f8a0fd26142763b0ceaef1c072aba95c71d5391177183a1a9a3245e6e1a757386f92c5ffa763bb2d7884a0d4e5d855eedc5519f7cfd78542a366c49987ee234bd1e8d3ea610f61dcfcd48c0315ec7449562e830ab13baeb36a41a746c110db007f521b3de9dad4e0bf7d2d3e20b776efac3466a67d0d354165c3167855c52bfcfe0dbd69fcedb174dadcc46d48802ef1bee0cfe3dab3cceb1e0288c3db17101497fd6907;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'heaecf314bc27dbd37ec80cfa72e8559df1368b95e3cc75cdb1a82ea7535a30072f9b9849909a6a623647a15ef638d6c14394549a8c1c94c2df974f669d17386b2f2781ff3e05148a2f7796bda0e387a92e5828fe6b22a57ad5fabab9da615aacd47e3fd7670f16268e7435846ce4463fdb6a174e626df242cd28cc13388515f40d3ba550e976c16d005113066c5aeef6ef89cff20942659e58e14da3c3746df42b86b21124014fcd61e16c8fa2d5f02f7d624741a420c6c853190170b1ab15d38da5f60f21913e14c0539cab96b77021ef4cf218e4c45ed39e80294688d5c4ee241244e32a979845c21793b5283cacaed38dd465599a2d0122240b4c264807ccf924a172e7cd58745de315e83b895df010f3a3b69a19210a3b3781dd0a601db4dba6003066ef7e7651da1da16285e67fe26dfde48513986f2a565a5eb66e38c27420470c5b28d71231923375bb687d23e9023f15e12bb8a573e5371d985c8f7ed5c99193b9ce3fc1a94df355209e2bef6510356f8941ad4eae2e97050cb2820110ec27636b4ae173800699b750143018cd1533c66110bcdc80c06455e50b1883454ccf1b4c31f814205dcc8d657d1ba516c6b3ce8942c8866ad74c6e02a247414947dfe65aad7ed44cd49e425d80ae80960e9bbbab614fa2a6e0a4bd5892c81e27193917ed72f069f82efa92f92a449b089256f2e49c0db62f88b379ee84d8c501f8531dcb7a920fb5ec1129d6c75b8306ee3f3d1529e7ee407aff4cb65edd13a02f7dd3fa18d9122af16032b2d004f2b75edf9fd3422bd9f77ea605bd9aa0114d923a65610b689cb5ba23dc64af58dcf43263fd787f3ad9590ba41d24a716a1bc69036ddbcc652e94aba338c12747aa49c379ca7b83cc248b0298502d0e4bd79d1d3c884a38449f5d749be849cdeb66d801dfcaf323f480a92e5424bff4d47b9f66b5558f1e9f9431f92aeb35935cbffd9067de3b50a0d9002d0f287c9ca2877a7aeb5ba0e93f4f6e753b2e9a8d4f91db2cd560787f53628533d66f90e02779ed2304d8254ba32b2c894a94bb9cb5c1fb3ea3282255345631721fab3e6041ccbc6bc6fea734ef7f718c0bd4c3859d77e25f68129bc433e85b8abac0cbc5306abdb9d5c492c39c0b6961a57cf02aa5bcc2f0a0147885967259dcc4c19c14bfc961981b78013dd703f43943342f274cabe63a910e01fdb6c78a06481519256d274483f5d888e645d2699efde79eb3ab42d3811d4b1eaea593ed602727ad438ff3ac0fba8070ff1f023c787b98982408284af55e4f6554f8f5af819a3a45a0f03a08e6816d3908ce0809c97655d73471b2607c08580ce868de559d9d338d2960440d2c46d42dc7cfa776dd1c3fcd07bfb9f5d22c20a8a22b404b6b7b2d2e90b70964ce76dda546d4e4e05272401578220ba30902bbbe2f86751c8269abaad9910e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h52903c56c500b504d18ee1fd56edecb88f700e1934973134092f7bccaa1b455b51a76550e9ebde03b1fb7b603bc91431a11feeffab7c10c3851ff5de3638c9bafcb177ab74fd87d98f5c3db3fa92f3cfa5f7c4504ea94ffc50a39580107a5a9657fb2964d913d2119458ef379c287ab962f6ebcb5028e6d1c68d1b6eee03b3b16c18679e7d08897640c494b5beeae15a5c1b2c5c9c65383f2260b7b16bbbc2d8d3180dfb9ac09e5a63895a59c2e5a345dea8be59c42a1f7c2608c2971eeee94c815af578d4578db1125773315f9682d33a88b26c20dea1c0f9d517ddab348e88c07c2a98437aad8d2b13b8b34129cace236d5292635760774ccbf1df417b341f79f1005347f4e72efbc85911fccd892f80fec6f523cc9328e93ef4e74ab58fa953f0ad9acd23c14abeb0063e801cbc5c88f89898a596a55c42e2daddd2b8baa9ddc9f8941dd88f17654a572d7ce68611d4a94b3937aa7f43713fce2a912fb72dabc75e8eabe06ba80fe13f7a4d38d1e38346f078c021ca2ce211d1f4161bee41085a4cd2aeb7564d85947891e122d494f58fed1cb7bcef70b9912527204ddb184997d987fbabc693c050000c87ba2f5c35cf230a9263387e03b79c1bd57c88ab144bca1c84bef9706dbd04ff1519889c69beb47f75b239341c5eceab949e52cdbf00108ebe932302a1a4f73fd8e95d372e5877644982cf4490076939c6cd39e09f4387867e5c43609c2786a33e4618f284487337ff72f3f0caa1943e21749e9f65d6efa708e48891ddaaecd7965f9f9de312898d602c63213438b856c14307e61c7f039db1083c4444e34b6c178a5a362ee97b10d8a335dd3a4ca20150ec358e5179306b8f57512657b9d3c494de2a566c0464de78995ccc0e3e85c514f8a547c7e8f8373c034f8807997077770359275def5b5be3dafaa12629e9e6b493f56724001c141883bca9a3405354ab7db74dee7d154929155a70c446b2aeb413f83eab7e909fc8c97c60d9d75cca6eeee161bd570d2b4e40bf43bba12dc2c5f19284e644be9465db53992aa5c7eb63a08dc862ea9786c184cdd16a813aba8fa77e1369166c466ba24ed2c48d6bb365577fada50511a5d23b127090eece3f4f90abf0f88eb2833c02305378f9cc0e577ab14fd177149b8292dc697ebdc5d3585b63ceafbaf5fd3cb78f1092015ee917e1ec230941195b81f6ad04bc64ee7c175b7b27f2cfcdeae2446389a4e9939a954a54e8b73625674012a7421c285ce1533f464ff4213716d55536490fe4d339121c84c8ab3db819246f24b1de241998745aa1507c21b429396ba4ef0e0f58149da1a5a7f973cfe53a5bc5c0a174a587573d67b98dd6168f747d1502c0fd865d543e1814af444ce44412bd4eb133ff78b15b5fe17b624122d6fff41f04a5f97ba896b1a7f82e710a860cce9384330853a5c2276b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h79a4fd440b5dc6bf8ad66f94d76c24e859e9b575e4ec18c98f2423b7b59c05cb910e6a75956b62116ddf2c2aae9f288e8781fba69403fcb96f359a1113e26c81d591ccb0f2d7e5bb245143ee2e827d6e04505f0a86207adb9fc76618aa08eccd8b1558dfbf5a8b753b0c422eb7f45c0e0ac79393035fa6bae0a576cbcb9436f199912e3fef46b54e0f70532033815dfe0825862bec089497cdf717981cff098327108086d4c5f7b255d0df3641e0aeaf591908ced251f023042aa262c6c07f7a9584a1fa251e9c2a68c60d60c1eaa58252654626b2c842ecbdaf6967821d5dd2b4bebb20a7b448075175052381add13676e738a5b0949d87395d1e44b1c54ef40352477907bd9068ed25bc75a22521ada53f16e413c7be66d4135d5d5ed76d26a49042f1e218b53d6fb7cb6ffa921fdb93cc33f2c5dac4ecd7732403a15f96eac6861e57fdd7fec031198592ab13f1de85a077ecf131d53429e36e4899cdd84579a75fa39fc6c96e9784e9862c98ae04a4f2c2e0877187642666ad5373ec9ca9610aafa7f7a0f9525588925dab41f0ff7ee633c3820c2408b300c0e18e6ece736d120ce23e1ec3cb869f75bf4f9b69ef905c49ef8e6d795cb25681cddb340e5c6c4f9fd42b065bf1c734defce0578f8d7dd9a77d8181b918ab0d52d6abc5520fbb260f5852c58a8ea4aa54f959ca19716301ffaefcf394f91e6540347cdc8c25a53502caf336043def52eb6172778130ea050cd1e82daab1799ba2e5f117ee8e55da054216e8362c103151470aa0cc12d6b48d6cdc568bc8c6200faaa403115ef3f0abf6b4a336ef857de9600d19c4e429ea6c428c23364c7ab0b613f39b1f7561721679d3d9642e261080770f28a8bfe5163d202a91adcc96bc2247b023c0d00352fa1aa25087a6ab199fa6accc0ba21b692a96bf08b21d9490db382e0f7f821ca837f1253fbdce6eb5a2e20ae5347d35f844b7e69f437fd653ac37b9142e50ab53959b0502ccdf536799a40941463de0d3ab1033f89c90bab94f54823f6f8dc83cc25c112dd9f8c64958b6178bf6bfead2e33ef598bbea3d3ee0288a3695b9b7f09581d8dad867f440ca90c59fb17b5a652975a27be4c197897654fde6b8a52d4f96d5ec52ee0baed197da6ac98fbe664bf1d2f3fbfbe5006df63c9b4ed06bb383dd0659f6d497c3874cfdcac400ec01b0cae93d52637dfb74698cf595af969fb02df830d406a337fba1a9a0a6a8f2652bab7e76cc2d055ee23390c8693ddc6f4f29c62c586f57eb059b5cc3f1b16b105933857ee8a4287bb2a9d80051faf4240cc33939f6bc6e7372b231a85b620c165c9e4bbbe78f98edc3a337cf3b465b4231265757dd95a4ab3f9506fa74359275ddfbac65fe36254d59757ae70954678c741552793c2cd72a25cc94b21f398bbec0a891e4ee0e37d4d30b2eb73004f3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5ac0f6e6dc834a470a0a3232eb1f14f7bc8b08aa83e94eea15ae92fb7d73d35f762bd68fd115c16f2a5aa253096e9785ac1167558aa1e3e27eda0750ad7584fdd1730f9f10aaab92f7958ebb316b564e99b0a3c7f7f1a0f6b26babea68203ed63734214d153f4d1da11f271647d7771907374809aa1c8d30b80e1fcc87cf1c5e5148dc477be4aa29f372ebfe7a8cda246c26b666f0245e7946ec5599590a94d1f3bdda2dd76c7083b5de1a4fc0e35822b86bed53d535d6e3a3ebf100d185109931a4d11f70e7b88d59a4e462a981ce5ab25065117cc81c83e8338a9911779224248a143333ffc5be8110c61872aac5752e1f0546d2850651cbb03389fbdfa3db474dbea81263b6857c7ac821e8e78db93c2778a9c78d0a5eeb4c53bfe4e585dec820c1cbeef07e25ecc4d2dcad203c354374f1faa177e495efcbfd8637a3025301a98ee7b052a7f7b1298261bd73e6d1b4b3f98f0bb26e8f65c0d77e3a4a1f71eb12713340f39e5e2e78cbfbd0f7037b049650862a2ed2e4718a39a5a55db1f40913b83a9bc923abc371a8f87b1ce7f749c04082faaba9b14b138d583a03d4b9455d0d7acac8a1e82bc8bf5eaeb218cd6c38c5922973a4114c2d57d86ede40d9703b59cfdb1acd84966d4a692dd01117b73654a85082af75c107a7497909e37a887dae91c10a994d83dffdde7b40a5c4c7a3575edaf8f724beeccc500c112c9514a969a46b48c34d2db1e56ae11148fd6f0290d21109e7da7bd335f94c7a361ab3f8107e0ce09acfbbc5baa402b52b597e2555f405a111e4aa98be6bb85d56d670cde99594026b179309434c75f7cdf4cb0bd1599765c734014cc9a7c14b71747d22b8e27055147dc93fb8fd58d13545d3bc43b07d0577379f1e1bdb972864b851ef474101dcb6fa45f4bb2cd6bd15960f291b68d98b4dccb7cf147b7f5ae46e6aa492e860849abbe01dd99a4b77bf095494f3aff47b95fa662a5fd3caf11cff09c29b7a42b91dd89df49579dd3e28c7ac6883c44d0df26e38ed5215c8c3b753c9828594d45b8a366a524f6495f32c5f2781fe1f4fa50b0334368e13cb7469e07ce4245a8c611026f18e1d38fdcf3bfbdc781c3673e61682e91c728452de873a26dd7c36a2c5a028c8f12a9f5a9f558b00a82b9f80f3f00943872992c4c406793964c55596cc61969c0158e9936512648e12c8afbd42a929e30e9e5808f49bb46066db81ed4499982a6e1a9210c4446a5db5b2715a2c4bfca705dc51aedd86c2ca302d9a0602419f4df9d14f05855d947606624a0521fcb9ec6613c3da9475b5985553dd4d193b1aa17acdd1e252b6649e9c4bc7d248c8e16f51da82a89b51e101957e4f9b728c322f840e76ce818cc1573e85a844087a1c650d421db29d8974ec52164daed32b521826adffede9266eceaf70311344f2258320967762362d02;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6d94085995c08a3e4116f328ca0ad497c35c05a5a650ac97d4807d4a7249bc5b27338859b398ff9b52793afa428a1379591552885f7858baa213d6a5f8bc0e30d5b119591bb2205c1f52e21c11984fa54cf72f26b71b12e3395e757a01c01db713032b4b050764bcfaee473ad9a9271600798f928eebd263ded20155d2666d9a812b12ce06b39bd279b6d94b2a03f9c730bcbde894388a197c3903d2eaa933fc7b8e5339c3a19860c9f6d40b02391abbed3693febc6f7f8a210c3497cfd1ac8d1ae4dd2b1fc661158d137c38228c2fca918050231e0ebe99d49fc6272222aa9e0fca4c493efbeda0a75fe6117451815318433b81ce4117aa17ff05f3cb16fbe05ec41d488231aaafee07dae4e18d1d032285e7baea01d1dadb297f947fc7f64e6c062e8d15a43f8db90749e0f20dcb9dad0a6e297c236d59df757a6e200e8549c87d5491fd0335b4728eb249a175ac45c07f28a83353d6480a1c235a8b77aa655aee1411f40b19b0dfb1bf1ec10ee364d42f029718efc24baa041cb62ead66cd5b30d15de28c955926bade3b00f8f4c124b6a2c3d8808898e3b9308107bc3ebb5e87d42a0ab361515dc8a7c4510fd58008c82ade8f60b8da6c9c24e0e328eaa12386ea636877fc60afcd147122c8062df1f5ddfb0d18afd3f59dd61d8d5f22bed3bae9a43496a753752cfd146e8ae1640189c9cd3c116922bd522c3d7e458ed85543487b2f79141f165f24daa3135e7fd60d8fd8f07be60cd0b3baa56e2cdaf7ad8ab561ac24f886d6aa758798436968ece6be8299ec73496369586e4087b495c0e63a63eaf8984ba6e389b9a64f23a0eeb025ecbe600f552763f9fd948f3a3b93c5a4ae74fd5cd50b912c891ef742f66db82131bc125e9fd43f4593c5a4b6389d893ab6ed6436aab5e8ca73d723cdf17bb14ae80d47049f87e63fcd21ca44f643ed66c2a32be03e9770d2f90b166698beead641c1dde504b6defe91fb1e7489cdc116bb587b87c00b1349d3a95268cdd20516c1a3d8efc4e35b83cace9ecffd7ebf65180112b951b9fadc984b0b4e5419f291ac7e3414a801d6303d64a0839ec232656c66f8ff851dad4dda3fad4498ad0269be7813f6457c92b43b9764b5babda83016944dc5cf87e121a9f778312a41ff0a63a20ce862cd301b6870ce2fa430c96eeca36f55ed83ccfa55d022ea0cf60dcd5bbd831e451a0bf0039cb02ff7cda110bbaf49b8f404fbc62cfb40f0b6d6d258ee69520bebd1a403b11c9248108238b8883f3b1d84f2a1a98fd1ed8aedafeeaf664f188febaaddb7b3b68ecd5af445a648c885b8d896b4cc3a21b5a315efc6a3f4edb64d9bbffd71629b0d7ea169f0c04bf07f91ad222584fa1d33183bd3e713756ba5d6bb5f7dc055ff418e2cf556e4d28cb4053d9d018e6cafb1ffafd93b3395f4a67036facf09394d5ab035;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc4d8891c4124a86077ce27d7be4ce5926be4caec76fc2e77b37a3f0b801bf3d95e5ee5da10c923ef945252b519798338bc4341f4364b85f004ac835d59d52017c81034cf542198d1d66869f4e1dbbc7d24a367f67bb6c883b6f9b2fff9ec3737d55232e7320d14a33eb6be443da04104165b58ef7b8f35d954fcb93b68ff4bd2bab34f35c279fd960d11eabf25c22d94eb09cbfdce19431b3bbb4c90adfda0532e94dbcf18e13b4bcbf3a355fdb252e39ec2977470bff6d03f1195eefdd4d2da68b343e2585a1420dc6def60a60b4aa97183de90eaa6c46c916237012fb37dda89d6871e24bbbe5df4d75df4cd5c15879942cf07be54f66964e136fae4f8ec640c148cae4ba7398da5645d7310b7d9f62f46a4b5f92a7fce2e96213c3bfa6d716cb860581c18b60cc6570753ad4fb62d1b59874f29d75729a6f32516c1e1ff87628c9675cb96de381b24bf37ed2b16e70e92536c18ea11c61c4e6c9294e78d0d80290f2d14c97355ed04561797e8a4e89d77ad67d1c964fad7237d352c13d7e6e4f64f589e5030c629e840020d8f674793250e13c70d0cefe0ecc0d5660145857dbc39f4e742cb735744352c09605d455fcb59174f18e5339530bd81be6309547ec70b5d90cfbf80d98445e2b8cbe3800af58944ef262bd9cebe6c14338a0992953a4fd22d913fa0137a13517ce35d7145406a83ce0b3c67423961121beb5f25ae9166a34d99f61bdbc769925def3f4c596ede93df54a0c6e68a5c168be6d5e842e55dbfd0b98a89e35a2e839b0ddd4f857f1e653ac0c9962a9ceb656ed80597608e72945beae723d713e1838e603b6d2584350da0307f279fd28e1aa56dda63e1906e5c02e02e1096ad0baaa8fd90ff7a4ef98762f402a86e8678ca78ec00b72d538ff1578f143c03482e3324839db9e9a99f46fa0ffccd307dbf049dba097aab51fba168e97070c301d3e0639f3aecf6f3aac3ef1fd750b52fdcb985637b728dae857997fa950a0a912aa2e0951387e0a1aa01b227aa8538c28b4e84206132a7f31eb225c7ebf774a30abd89edbb63d7d713586d419006d2728ccdf3e78d937e026ea57cd46b15f35a02fb86840f3d9e83b9045b9e767969cb0287c563caac5e4544a07b0e67cb26ad6cb197e26759df54664a728e07feb86fc02375150d91367f24b9da399e7bddd65a8296c4c2665f6fd320c36ee14bca8edb2f80dd34c4d6de49ce390b024c1557e28e4cf555613f02f056e4db5d3dc59b591e5c34c1898289613723e1cdad3bf6823202839d7f6e0524e62fcab2f8a56e14564e863805f80f09e9bfd905bbece2f6358c6ab50b96827dac7d6676a752cd8106735c7f9edd578d9741fc86b143f6f5e94f79aeb407b20372535d48fea7718fc18aa31de9a6625528609379471ae715a5765bae3ca15cc0ecb7ad53c222f4ab1cf06232a6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hef6f9be1a880b7b09dae7f254e71a98ab2d5198b99799af3736a6918ddd46b9f6e9fddc98a997a2c8f5bebb430cad6cec4b4d4dfafb0dc915ee285baaa1590bc6a6ff7ebc75a74a9f57f0c0492ec39dd0e9d795167bc81dea266c3d54154c79d5a273ddb977a0839abba41f1d9e58a24b0e1da38825975323f39f91b0f777aa93c6c9fce95a98ce4d39eb8c1de6589daec4b04996d8f42c75fad8116f76aed40e69dbb6cd0e1d35a673a61d4f2291d3fc48216e436a8fd2aec8c57eaa0022be414c3e0f76a63b1680e6d1d2897029c848d18ceef9776726ac75ba2461581eeac93ae300606c06b86555297cc227425b9d241d2a372bcc642a57bc4a69d51d670ad62f79cc88d4176fcf7100ec0e1442e6a58f1312498a4587aec40240d96634c76afaf8c3acfb94855f663e340a9975024810d4d6a5671291245ac7ea023ab5b9a1d3ad3c855a2b0dba9a6ee3127925aed880bd404655124489963e67206b6a5743752f92f372691254f299e43409637e9a82019c2d82b8e634d9b08828b495a651a7179a087b4cc617b8f6cf84fa867939a18ba6ef7ccd5005c988c7944c0a486d7225db344b63a65baf97ea39e528e6a089a49bad7610f5394c32bb8b98a23a9291aa4d74431d87af6cd32f8b5d1c09393cf1c91780d3c9a6dcc5c0ab3f240208f8d8027abfd6e633a8eb08d7c7451f5682ded509a65c32df3682e20f6e5f27398a6f642d7870d8858ba70802eeab64122aa92af5461395b4e82bb4669866221cb1f12f5ee53409f6a91ca2bff7051e849d74f41408767e602a17dc4a2debd4f076b8ea2ef6b544c4a1ea07e3853ff8cd8670dc7a7d3eee006efbeb592a0f76ad96fc04f120da8de7d9aebb73a00038a818dba1fe96914de762065ddefac7cdaddceb34ca2c524c43971a033f14286bb354177cdf2d9083c5e0aee8fbf57df8644a50e337621f9d5d53b2fcfd402c5c61c288f6780bbc051d55839ac85c8680418d0019b4cb660a03cd9c265c32297968a02c9aee6f9718a4b5b29d0fd2e7dcd160544ecb9ef3324818c63d08e397968bc797da83a12724bc9698d39c8a95760c2314afd9fb83be3a836242986395e4793ee72909b75b40bf42de8b2d8bd259f7498bc9c8197661847fc117883a898b207abbb0f466c056ad2890cf5411c5a21792418ed56759e12b8472503c34347c1df424d1a1c79b0652448b1cebc0877f38c166878b940c50ad21886571b0cc88dc5261e6fa23b2fc91ae5debe36eb3c66cac7b236544592171ea66d0cfec53f868c345c8326dae139ab070a1a7cb2b8dec3f21ce256124771a0d93e1888cc44f2afd2757c1289de72f8d60c7ada856f3d73676fad1b2820fdc3ec60ca56d41e73fc51074675d9e934e7d71ce1eb183b5c028d092cd98ce84cfe45da04f90525700dbb7707e5752e18c45d6f7d69ea80;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb007a72cd63afd47211c0086debacf980b6447999a95743353a125a9b262461e64169c91e33e3751ecade5be07ff272c3310c0fb6c6d5244c2e3ae721321445c5292cdc7f26fd0b26361bd9e88740bae0beb24389dff4b95d5cf5599768533d760e5c787d558d30ca52bec6c270d0255d8bbeceb38af57e4d0f764b0838893c1bdc1839d182d2d457e563889cdb67b49836803d5203ec67cb6e00d71a9d20f751401485895790d09439b3aade28012365b7f0dbefc08391f3ec62690990714d546fb995de6c0aebc253207e6016347b455a04655e936ff023c1f9ec63541ba97831bf56db1b2b993334fa741606399d9369d951bfe923e3b3c542258ec21eb789c5738e0588e0f2fcb5a32febc07ad4dad14d9907d89b8b4881a2ede470249c3c5f3c36e2a03857e76c6eec507212fd7e1686b17f8d3164fc04ce4100b074bf75dd22c5937f6522a9879d9b3cff1bc5be09f9841d1089168ddfe340f55f3f785999cf48972a523bbc15fc9fd796d9023fbabc6e080aa9b4baafe98c8dc37910e795c4e64086b23b181cc385d67bb105621424f2f7981115fccce9961021de7b260e0d255f83b9a26e9fce8ec210a8af88b19b115f03d22ce0012bdc9f9f064befe81a021fef73d91632c14ef374fae2d97239a1a5d616e972c3f1049ea2a7fc6aeda32fd9761064e560cb4b7542fee40202f96b9acf9d2d736bc06e4127e2e5a358fbf19b9213c1eab2fc6795d1cd924a47d35e9c5656e6772255d964864eaa4a0f2a837f701694a500e4ccf16eccddb8da8ffc6015bc3d0fbecc4b128ec128c75ba6ea1e3118bc724561cedb113d86e66b87c823138c7c85e3b0c94438758313e5dfcd563a2b64f8e7a76d7b42d31ac2751ba9f728c3e2fb9e222e8c9dfae5bb4ded8ec6e927b68819c467ac69370ea22eaf466ce0cb2584ac01fc96f3a9424fd4270a4edd1bae34908ad0c2bdf23e52d01619a531978024d471ce58b3bebc55761f5a96ae658efc8d2c1a33feca0792eb0789f69c16b0b29024a6df4202ce2c0be6609b0bb60108891187f83cdc771144631cdc5e9b206433b4d5601f6c454dc93abef6ee4e37de4848f48c43f67322e4d0274fc8be101b8387cba32c09f3df0731aa068b8bf9333168286e840f1a23c66ec864b38855515cb03938d6b9ee71e53996bb79d18eff1f2a8489791bf285948282e93a39f7ad6bfa8773a3a79105898a93302d95da9ace81a4f0a9a118365dc39a5aa4a9894010939d12d710d6f197636e90f2ecad2c8f8f29c834d9a0a2e575476a1b3d72e1b1a672e8288093aa391da3dd4bf714069af31c599aa0a843957d0ef96c9da2df3badeaec59a49d89e5a86f3a07c572dc66295441d7b9b3d2d6673f0747b069e96e29eca3e7cd00d03e8fd065010291d46fa0ca8fa18c6d6fa8dbff6fd87b9ff3da3a81ac74fc9d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h46b54a3e56328ca9425ddb87b9cd11b67c809c82c5217eaf97496adb55d56e56e9ebaceb8b57a78fb6df56d7cf8426067c17fbc9d2dd5b69e5200b512cdf21b27ec6b696e84ac9f8687e44e6e5ab003142d5c179fe7d1921aabedba2e0b20e620dd714ab8d33b445cacea743ff08a5fa62b4b6711f458a70b39095d79bb5c5796027a9bd4bdea09b71bdf3aee360b86867c273ed8660afb2bc45a13f729c5a8eb022838a4d7829f475741260feae0a3c88bb1f5f7611af71d81f409d3ed2c6f0252fa19f2c6f0cd74d02aaefc2592d9c00a8ba671109adb5b48cb5223b854471a4265662301f28a89419ba4c80f8c0ccee7d1305ab27adb0d770ff006cd44452ed95773618f3ef6b3f52e5302913d8171cbfc396ab1db7b616c2a9c09e53582d069b3887d5b99be80170e7570e0686d1c4789e4a3046001be40d63b97bd62a25e93a93df31b634443eeb789f87189dd878606b31346b9b5f9bd215d01f36939d582f9377eb621eb0c9a01ac1bc739769a7c341cc9846ae932d5d7eecb3b694899dc4114f249d1aee533424bcd4ea1ba53b801425d1a4b8596515114fc6136483de473f240efb5db4c23d642ab5b27ba396d73ea6943a2eef8499a590301cab5c72d53339ad0f97bbe3b1b5088f068dace808363d50b08bc13cc8c9b812ca2c4f68349a4f6dd9f0a7305f01fa6b20793d01d43749fa72543c8f579b90be57b894fa15013acb940e332d4299149d0d5ffc6b361a08de2970bc6e0789e137490ef5e65722845cf30519165544e14390b17015a07f50cfd0f63e4c1d4284542bed7901fde7b6ea44dd35d0bb5ff2e662eaf0987230a31d43a0f694f2f502547cba313ca70331c182d265c9c1fab3edcd29778e890bc1cf97835db67cbfbfd18d31d979db4df31f3dc2cbef3a303bad308e0cfd61a1556d1c41fe1dd75f5bcf59200b282e6b3d2b767856eb7db40c77b21b7d1f088e6dbb9480eb2ca5e9ea8e44556d9b4d80788dd07b0c6d1a8f7114bad3788d3253cbbcda99b098b36351cad84501bb0f083d9034ba00e0225b09b57a4646d71b6632891eb230eee4f249b02e8dcb1b920de1b69acf7127ecdfa92cf3f129968ac752ca52ae2f012c29184f0b05c43dc1e83c0625a0d90fc8f860d9a20a34884c4851d2414fc82bdbd233d08417060938ae1c754666ceb21d3c54ae2f052c21300765a5c8892e2245cf006b3727942e5012a2dc29346ed1cc35357e35b5f7ea32a8bd889854b8f7eabf694f4972b1c76dcc04adee9e1b7bbdc547b7628c4ef8921cb660727b80c2bd354fe8c8b626201acb273dc53118d2e8ca87ad46661983ebbe9a8f352c036424e4cd64561f9fcd4388678346cfb1c4db16f9222032830260454e37c07e334fd754bde8f7127d3afd3b6563cea18f108110a5b97ac459b4f926cb04de0cb5f41f95f663313e88;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6b5878c109eed4806300b3c8803de7264301071fd11d0aed0701ab7e31b40362dd8fac39ac5807b51c042abd77d6b5f78b2527359068c3ab778f654babad8f3730c11c6f3f5f7e118e380b206ec226f5e6b213ec16dff77af12776b62809b20b12e8ee73906d161d990f92c2b9f0e984ddfbcb7e037ebbcd093614e8a3bf41044f45d8b44678b0127387f834056fdb40c4a4d9b41fcb8c2fcedc35347aa1246ba6bfd64c322a3cb96ca7f1264fd2bc68d3e8759136e8624c98b545b145f7f1797143edf8d26a81ca40b89735cf9872ed44bd59018e9c4946a459eebf4323e261d03abebae81288cad17c000b3777f066502d200970cf0f24dfec515ff93d6580ff30c218389fc060d12166c7794013d6442be4dd3722770aa0cd257c9777c08f90f86015ea656d6196c1fd6fb6591046d5d436a7b9b93677a8e565047f8c315619b2ebfa60a7ec936afc7d22501abadc04c10a3c162d1a9dc7081d7c75e8805164de797ba755beafadd70bd39f8bbb388efb6c56c90e443ccd5af648f5ffb45b939ff90c3201244c407528563e77300c3a0060c829e166d77026f73c0b738570dfb8aef11ebdaaf4a299d01c12ed50914772b7a40189c2ab4e62284f315f90117c92087e6ca271084e9331b8546725ea72dc5fd257c4fdcd4dc6f2a82bea194e8c758490edb5bef4f9a28413f76452f21f96fd3bb52637ae5889646d028d1d6cbbb22a652948965d46e67c92aa697f0d1cacd92d7dc1682406a56d4b1b89b306c2b3db8b949aa953755111b2edb17757b0628a9b2109516d426187ac6d33552922a818f92169481c83655c330e4a0003adf810b18db6ee75588142e1210869becb4a5c027b4945feca337b4f81e2a437875b6def30d499fe76d9c3d1feebcf7a82603d5a0043d057b189cd1aef9ba98828ac6ff9ea2a0435b77367afeef940673498cdc3ed38660cb78b1544d428f2fb5680f1c73852d0464f8a35163cb83f85060f238d9ec31741b5af3b0bb5c9924852c7ac24ebb0f1385c0a4a583baaf641fd1c76310bf9f76f36b57dd7e332a12fcd32a2d4673c2385e6460a5cc8d68b82f2a6139ca3e90aa3fe1f9a76ff1943f511ae00309282480edb4df7d64b80048d42960f3b146d2af6e738098b17c1962bae17a3722b6d1881870130f8633f319a43ff3d0543881a72f097e6ed1a5473efa9ab80e7825f90bb3e600021a4f2e94e71a50ecfbfc43e92acf7233a469e0bcc07140a9cd7525a4e71015dc7fe333b26f550cc0c9363a1c4fdd7e5b936fc5c213f0994d69a8fa948e337c57813b05081e566c8db6ea82cb2791d6523dbeacb2808573405fe7114b47c2c64b54c2cea8d5a96280da8e3c55c730c07d6024416cbb3e773b12f162d29eb0d248501c5f87a459bdedde528ac32f51543c45449ae1054f14c19d65e171786d6900629d3f8f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h45ad78891ce59579aaad4b75bde66bbdc7d172cd254ca62d4576ab491aa180e6c02c1c0cedcb20c4b4ded526d0ed49b5b1aae2f9cf629baee2ee26abaf1ee18e7e05cf8851797436d47892a3a60cbb4e31dbfc2605ffb5c1816ad30d3bbf9b3f270db9ee08e21d8ecd4494b37e04ad56b87fa9e9448c4e88e1aa112e3b70a4339a0b705c34b1ffaf8f2e91a9d6c6f1ccd2a83263946c1b0399171c39d1bd833bc7cb8f080c538e59c703cf77722ad3cf170c1ff961f74fa2db9467afd41e26709f80bc55843bf0c869730f1e414f6034d88fa1f5aac2351e050d07d06710895542055dcb6c04fdf6bedef1c6cbcdd26fceac5539a4f9cd1e230f4e18328591819b16177166d3e2151a3fa8ba0b2ad2d822a1635764e95c2321f8dcf3e4a0622fa13ae480491a40fb066ce20c70d2583d39c393d37f16971c360b0fcebd58e16f35d1b7ebe73a32611a5b9ee22c606923fc9acf0a536710435738aeb1f442d2e369b7b6f57bf883d3361b259b589499a3bdaecfabb00b90fadf908cd7aebf55c1c17bc26f136cce97da747a4484fff31a3915da411157dbe219b079718e73e15ef97735d6ef054ad41d1f94a9dde7e752ef89c3116b4af725959e734ed9d7fcc9f428bcb95bc1b75c72df2b682cc948a58c0ed77ab3c323091ba7169bf775827a24b5cfa3d72bc3fabb8260cd73c9f29b835992eee3335bfecae9064ac56d4e9fe9cf18b2a663aea08db4fbb8e282a379337e04874608dda04f2a5e6a1e0d248f59679b767096b05e3831ab83e8b2306ce2209e12f361c89915bb286ddf185e6d099a53242793d1cc745f0968ed41a8abc04d5abd1cb984081339b6a38a3686a0724fb50867d82c9ca41f584d2568c2e36eead864cdfa3774f0594ecdae72ea71c8f0201f5fccfeb197934b9511fb1b796180f79d86e1291d1b552ce3308eee4a963338f204bf3616271bcf75964cffc1dc6f90c718430bdd66b6cbc9805dc8833e3d6dccf938b2394859f8a949a71e039033145aa9227d556967d43549a8af810b4ac39becc4380b4e6d8011ea43d3c0ccb444724ca9c05d29d7ee060b3945e6eff0089638eaec98f534c6b3c99c4cc14612f2e27b6d2770f6534dd1e1b80ac2781f8f63a17681370f51df20a820f49f3002c2e5231393dd358e5d1593c44953588c01faaf4b40235f43a8e0d6f6253358e3a815f25e8d20a05f72f577e9f9ee0580ff1ce47cb6ad95256cab873a14a398400487ae09611c0a4ef7f8392e418a3d552e8876ebfabeacacc4b0d725d3b7b4059669c4f272a71104f879f64e59658975720d06705cea3f93f45c2c6298e47f0d382c487c79e147c9a665ce80e7b297adb6fbf839abb3a814dd37be4b3e0aa98a48b81dc19cc429ad2dc52a0b84692c84a926170d7bf7b89c29d6f3912d79e25ef428321bae58aca591e116f4476;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd43d31d9fa3f84614b167e1805f87d971e3707840d09c4579f4681aaac90e6e3b6db27313b02b19cb0dac54b25494abd993b0a4e10a5eb39916e7ec7ebc766a884258f93e3af533d3ba257633c30cbde969d755d17002729f7ce17b65469f13531dda1376a10c23941770d9f9b48638ed7b4ea40e0a4986aa6c475f23fa0f4043c6d3851325c2f08316fb21af3cb2ba5b02517423fed6023b51467443c43c28cc0b738698f765625122424d7d66aed3cf19101130c85e2ed7ee0095fbeabc6b965f2446b70f8daa8cce07c5df48a754112d67663b84b4ff30a5c3522ab23a0137fb1aa44df083c5feec53262061d994fbb4b072e23818f9df9a8b8bf84fd90aded2d97c45283a7d4cc1e93feb4807246cecb1d64cc445f541efe034d6521d896c6a73aa8996e39cb58e04a47ec59c619e8c61ce47047659bbb34e60e35d15dedcad4fb0dcf0161294324e8af4f605cf864b054298ef2a40d32eadeb70c5c82dc684ff02366335e47eaac27fdcaf3e2b1cd2d31900e3a8677018a2f1d673e2e8720c6ae36403e51921722d29d4ad0a5d182ed80bbcd83e7b42ff22844b4588972d57fd339f81361d8b38688cb24c5182661d2e82153ead093dfc025ac16eff8ed3a7d351cba37c1ad2dbfd7f1043da0a3b5f8f80ec0b313fc1b883d64d58bf573797beaa31012062f159c2154727b9310b5a951550ae1d8a53cbb6b2d1206be64b89dab7e9f3e9ab229c46272e5ec77d4925185d74376403b4866904598999693fa7c289e9a8434499be7b8faac38ff85c6e9d664e3ba160ccc0c0219e0581697e3b2cad114f47054ec2fed07ad641e30ac01424731dd5e5f275bdc3601bf7dae1d3ff7b56040998c6b0cbf6d16040baa6040a91ead8e97fbc7611a44f0c55f710cc65893ecb625b65224380928a40ee93ff5433d2605f2c4dc1f40e9b702b76ab8e895848bc0b08b994bd0b4d8ae2bc83f45676e4247dc861c62a0f40344b9066500ba69e7748e724ebad95d098befd33422d6bd317aff63277f81af33d9c3f88db8217dc704c6ef3ba76043df06599c6ac6aadd48beeaadadb591d8b14681ce38bade3138126fce0e6c63e06eb40a8593bda3268b86322149b6cbe47125293fa616e188183883d947b283d1ee60960cb1b2323f1ce366266f1a8b8eddabc354d05aeb3997221bbbf62b87a80a248cc2fa1ac489c193fb98660128af8c36479eb825352d271c81aa960c28ced55d53fcfa428007153c7ffe832728ba8f298348dc405a057578d0316709b229dfe9c20878e9ecff8b5a91a812752759496bfa0ae1cd6b688c0ed488b8ffbb0a9006579851ea5ac3019a8dc1f1e5385959edbcf7ee82b54d7f09cf4221cb1cc43cc26050e43d0f7779184da3b441ebc628d5e041252ea0beea102a83b4db72d3d5bfa3cc6f284d86043d6a7605fad871124ea044;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h727a56eb1ae3b90243938c93fe0af3cc5be43e0716f51ab1a0f4ecb779dde2d1989c70d3a3f8d2d3a3ad59dce56a28dbec78def1bfc5a19f3b3c3fc1cc205d597908f3f56b276cfd9a3e30cd6138c199d2664385d7572d73547a50f5f2fc79f0437cb8598f29641bbacf5d448efa5dd6b33c3edf5dc6a3c3d6c38e34ddbca8f533043abe43c993733d9bf2a287606b472f9f8e94e65365307079b28f284ae09bc7d10210f2a43e1cd1babbcf64be5a7a1daa0c94d2451b0ba2c0d6b766650f1132f2485e0314bb886a29c3ff7c87f7d9563d63802423b8ddd059e2e78dec263067b836e938e2f0f5924983acddf24e14ed9833155de80663a4cc3beb4587a5c91a929b8b7b25ec8d49aa016ca3afa321ff816d0bd5dcf837fc8cf9cd7c649423aafb70183fc2daa5210b0f5a306769969557fc2274f317fa8c18b35298183e6a6a7072a28787fd6191fe59593ffbae04b17b487ed07544d949b73ab04877811bd8d036aa4039870d11a6a6804c34297b51d9d121ee798e62e8591d64c8e565f326bfa687b945787416a6e3dbacaf5c9088cb645f62284b24941f0bcb0ac6ab190a14c5b7bf8d94f2675c9f2bd895d8d5cfc11b8e469d54f1290251d354d16889bc5e9b65adda8b34d263f3aa2c88c194e9f3bb49563a263059aa3fe0aff6226d3617bc8fd80b9f2e8ef67181a96fbb29b6c31aada9390f5208e51028d024dc62bbbc0f25074750016b1c136e7d9acf6a2f58534aefc397a46d241aaa6d642ad39e06d3b65e747b37dad1a9165794ee9c14222865f3441278edf7e032c6e8ff766c1423cd4164306af9ce62555c7ee542666936d737376f285a4e22a31eb35b1acd79c942858f1938ae7eaf7f7368a080470d39a4c94096248fa8dd6dbc3fc6f32ef44909e95b9e28e2340d9a582a344b89531de776df6461e11b139024e1a17b53ab5a808959cbb20912886cff84ed47536a40e4cfb050a7f2b51490b10046d5cf601bd4923d08ef3d3b641bbb6f458fd445a94a0d924f6367610e085f868af978de1fdef56ea3debad94970bd23cb38887b7bfa1f938534637e97ba1f57fec9d69041517a28857827154482f7d8e2f81d3ee075960464cac35f796de1db3f0190d1aa0ce145ddcb22e61edb2e4e369023e8c74c9e0b23fbe024414343111576abec7a8942391174c2f5f15a5a00ccd3bde0ace2b17d35b26251b20060485d36bb6fef5a877d4263fb6cac991a668d7b6089a842ba5054f76f853251fa9f60cc4ff206ee3476b47958578e4b94f8faadeaa8f068f12d0aa9d5c25eba64e3ff02f5d16bcfb9a69cbf4c49369e6afa88bca17b4c790afab4f48d4045ac4231d412b76b9d4540f14dc1c7dd39be8bc7649f7e8b4df18105e1b475d27ffc908977c72581f640dfd6eec9befe89f23714dda2ce8c129fe5013baf454aac9a84c99b81;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf92ffdcfe9850ed4e951713c39380433b1946ce7aaad66bb2b82063d0cb4c511ec1a751a83041e4dde3286f41ce2c5b30abe73db6d45a4a99f400f5d6d433d5301345b6be6356fa14d73e34235015d3bb5fbd77eb6af5bec45f5b9b26d7407d8b312812546b6da8c8f4b45b467ff827c8a2822bee98200ded82651717028d9d3942cd948ad9cbdc3bd0160986a2789b6dfc3872980ad7182f0b2eabc1b4297193a6f189ac6aa34aa177a78d359bf0ac36aa468af75a72043e5c61e249d184d6da4cc4952994ea3693d564949a87f06a1dc6801f9332dfee134a4b57bfd7e7fe1376bbb67b8ab396211b2ef803b1043ca4ebea69a811886abaa43892fa447060fb56747387767540e98432e4a55fbc3b00684d3f1298ec946cfc69f2d746d4f65d8141a9c74cc3d267745e67ebebb5aa056bebba7db742bbd7604e5712ce32a058bb017272b27f479332abd5b56403428a0155b18eab4c4ce4d58f4664e8195a3d0abf97c6955b4d1852afdd614c710d29d4b004e553524d03a1de8ffa1302bcf0162cad470332d11e27be6d836ae57bb99308db6dc9a9325b5ee3a40cf052c19c774675ea2908997506038b7c97b53e22cc788a6e2fdf0f4d41cb9337e9128cd218bb48aec9b66cefffbe00877a0cc2f6504e4b3f1f62fc63fda5a8602461652ef4b5a282496b4a04e37ffc6b301a4fa31d8a54be56ba01a6c731edb762d31205fa39b53b82e92bb59b65fcbf42d690a5c0efde6dabde8a397e4bd542b1a7b34e41ac692c8fbe3dd2a3562000c38a425c617a6c2ec19cd95015bbf149519dd3b38cc53a76322a831fdfac6ad2d058d46c7a29dc54702a290c908784960bd7eb2839df376f00685ec4f81932bbf0d1732b26f4020e0b6f10fb4a716a3de82ba4991fb2d915c6a4a898d03a4ba2d59e08135ac132125b9b645b1f8659bb060ca238be994ad7ca762e0073f89cf2d90bc6e44c7ac76505da72229cce21e528a3e7c3047326322be9d0a70f991f0658f7cb1a69a5fe8cd829b09fe80e030252a02f75b750e6778be5e4eebb4bfc28a00f55adeb337c180ff29b98ff1dd0e0ccb3c8100a9969764e77e6bca37e248edad6c69f7c46802908ab37f2e1a1b8cff7f6732bae73705b4cef041212adb78727140cacf22606d20c5d648670eb29d9806bd9f166f918f2fb11dd456c30ebdc4f2c22424bcfab47b81fb60930e512866b24d0b4956e9d13d745e45f8d76faaa60d245e99daea9786277876e6dca425e6332e6b1f0622230fa01902d7d1f7160e431751787a4413e79d914a4e3c7dc0c81d1ec4fe06ee0cbb05e8ff5700ef04b1e48e11946e946d85f15d3094b0cee13c2ab63482f5f03a3c9797b000d315ccaa1b8da87fa3dcdf917e869dca832186d47f36a70c279e7f015550b292d37093be386cdfcf00d9690017d135a0e58c544495fc95;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4d2baf2aa9134252f9e6dfc55b91cb04fca97f7da9616fd0159991d9328de416ad74d033d101eada6eb5f28383ff23b7fbda69d807f53a9a91498e69e6267e4306d9b91c02150b0a24c244be64cc94c1416a0eb496475ccd81124d332e3c5331289f8a0ef96569b4e91621f276178a3a9a9230a55fab01d1ac524fb0d4291a485c384259f05e3c85e0cc0af64bbd02f9f1d11b95170dd38bfcebdd98abf0825bbf51e96ab697d1d2115f763a1ce559319f74d6493ecbf0f4baa9e031042880bcc162f1e0fcfacf832811428397703c07cb03144e12f7dfd94259c85cad2c3c0d8f747f519d835be2556051389a15758a2aff21cf9867445986a1c187b5a5e6e5dc2f16436c13b601b0b2a453e4e6cdddd0f655b8abb774128ef3608e796965631e5fe4912f22994b11cb1825ec9c60f9fcc64d4c3ef2b9868ba7c81d59588175c5c2c50c1af74d374250a03d5f984d433ca432a6ceb8b7f83cb0817807dafc131d1e2b7488696f14377e4795c1801a6ada9b2d8ffa0e7bf7d460f89e97dcb3b1d1f25e7e3151c9cff184fe13d5e4ee29f20a427189722ad42a954149bbec692ab9035b0ab19e30557fe005b80082f38666ec4710841916f2f3fbb78929343d9d190d06fdda7719fdd7d71bddf86a5cf9da0c72d7fb06f113e986223a3a1db269f57b508f9505e034285b7fc2fbfa8f0a1dc6d58bf2662e7f7d78129cb925402a8ee4dc12ab175f99a6f3f95fc5e74b73adff50e4314b649f57d31223550931519a472cff8a6022d995960aaa9a592899df6d2c977a44633319f357201ea465a8f55f1776ab1e841fa4047e767b94369b298f48b02ae58e33dad53be2b989639e2272dfb34d780ed64502b7c85fc0d07a307e2e2bf232bb384b9d28f8eaf2ec874f59e8d042891a7655befab7a887082e0188c227c8c05ea430791fe1a63cf8c08d930000ef0ccd9428f82070363d4864abf21e344e16ae34426dbff76b3e18d005a1b417d189bde0de16629944c8ebc85b10b1c5c7e12f84cb80564716f7d79d2423d77c3604962000f07687babbfce21592b192471521d463d2aad101bce691fbacd6380f9099d4dde785cb9aa3583e9390da8614d95c6cdb957c08ebc37baf4b776bc3623bf7c38667a780a7dea4bef60f1a6d858b3fde415a11cffda2eb1fa5e7aa82b0faca51386b965edad0531b6997e1d6f34a3f1b86ea6b2c263c3db2bed69af41da3cfce03ba83d9ed5890e3f55ff3da71a7972c982eef43973069937f83f864d42f86aee6166e3061e4543d20cee2aae543dfa89ac818c79e129a9fc00c179f04c5343c8ead0307505584980a1329113f15dd4982f6030dad5c2280a3e9edced7b65ca3320aabcf709c0178184aba599f29b6536d236f76d86628e72e53cd40455521f9294920d23d6b76ec42baee06ca5bc1f977113259bd120829;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h21e73292a4875fc474f941413bed98101fbe17914e94bd69d774fb65df0ae475ea95e748b5b7afac249143a113cef4ece643be656afa679cf3dc6ef5cc22994eab7d6befd41a50c2a1d67cf1f3c24801b0247b78f01486969e489bedc7b4f573040405ac5b23523acb9e481e32cc6311b1f47250bbc18b6cc4eb29be4297dc57ce3b97b6d6c24e646ddfb4d4737dea4f9e4d5d9809c0dd958e216a730aca7447e128ca480e6427f52aa35ec11971cec679679a5c955da5d9f26e5683059b8e3f5a0e631bee9ec01b3091b7cad4ac1d8cb49a343793221419686ccdc62e3a0f1c1a5e91fe03775540971bb136e33c1e2e02a4c9779d4124cb36d0e9b4fc974780411056bcadaa7ed778593f13609caa8d1f866f44e7fdf7bde12d48794a16f2813a467d8f4a9ebfdbd20a7a1f2b97baf96271259ee1476b97d8107af4e3eefafe7e37a39f5b01c2f920dd94ffece9bc50f51d891471417488510e226a75f545886bfcab0e504485be9108ae64a3efefffe626f13d0bde9f03271d6c75d58e8274de1992d62276cca9c09e53a547e89307cf79acb7b1952797d9aa862d26213818a943c2fe46954ef5c07dd1aac1cf653b5aa3d0e7bb1a4b562da96b7dd06ddd76b4e06c4d0a9cfe3038b6f768aa79837119642146733ca5a774ee85de01292acce9d66b4ffed09e5017c7edaaf76870c8543b742b4acbb33a85ddb3728828064b4e3e474a2175313960e68d3c13523cb10b92b94997037de1ad850bd0e5a3bb2f33f6d19f7301d4ee12c5b036a6fd50b03fe74c34aa817f1389e6b2b41be8f40bb19843adf36c0072a0952c3b0804cb01cb81043125a70a72b99e91c6e3562c46715d811ed8432da3a86ecf65ed388f7439b20f546ead3004fdda569ee40ea7708ea5fcb60ae5404e9d4565f8ba482c7ecfb16deb673efef9215c5b303a517c957d28513d267327b0330626eb140dbe0250164fe39c8badcfd98bc328ad1c2fd31351d7421438ef848452c5e28e8bf5aa0db00d5e9e35b08d57a706a4647b70bdb603b77998b9321d766d0d542c88a9f95d2aad8522ae2830a9656fca3a2780b7a380aea9782d9921a5144622cb4b8890c3892f07681a3378dae7901dd8afdc11bf3600023496841a8d60fe0cdd21b26ec62d3501b519c2ec0121a4cb67fc050669e8d067c2652617abe89d95f7fd6a2b781c8222fd4d9c39ba621d24502500a7e008aa13ad618a7ff8208944b47f30f8ec9ea0e9c17779d810e742b43b635fa268d82cc00b0aafb977e1d3eda94123089c1a3cd16bc0fc2e1b81e89d8007ffcffaf50f65852613096b19fe5b39d8c0f20caab906eec496c358cd04842b7bc798887290d42eb47c55580de9b85bb7672ebb4be83e6b0ec1b68de2609c95329d93012a9f2137610c222ebd363c0a12a30fe0b07fbc93d93d8fa02cdb1e6cd47578;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hcf908cf28ae3b4c88a4e2611598d393692c102b5af767ce95bd4f077f005aac4501b4cd753c12e47e29ae3edb5956fdce3a98dd2b5e556fa29f709b80c5589d65fe90f1da1a0f489c73bb4ae09e1d93b3169d6d238304cc65cde1a90e18ad90cd2ba4106d1e218e424ac37f1b3a520b6113df79fd4b97cea6a6463037688845aabb695d68cb4da7f021353032add2056b5e5add7ab56ee6ad2e3cf2ab2c058ef781fbfbd1953ea3667619b6c49361f7b6f00f84eef6daf0795b5bb62bcb1763b33c630f16f4e8e6cb7380b6ebbcd3112f1c36680b5f7a1465285a32cd6ee407762954a847fa744955415b0bef0fc6b3ff989c3dc730ac134176c4becc62a439446eb2665de108f7c9cd84f4e6257dc664d67c31b565b4d89efbb967446cede9ce693811cc6b78930b3ae56ab01530aa967cf0d89581ecbcaf885805acba816f285e2f749f41c965aec04541c13c089a61c4e57106f7454daca5a13c543f567677bad786c446be9acb2387388907a3f90ecca77c99f0deae7b519d1caf464eaabae33001ca9811b370979d64b91337279a526a699c086e566fa3c222119accead55a9813aa438bddf1b34cd2fe136c18045a0cefdfd16362ae186cef4d24b5b9eaa7c2ce26a23d592254dc2cd9cb253d868315f7423e16159ef31711aef67116ad51e4135dcff9ae0f2f9d3d03c23e7e7b9b4172d6aa07b7490a56b21605e010cccd2ff9d65b8764201a32fe61124346e70dae06f8d2b61e1a47a2743e027f41b768c606b87f605aabb8af93b7089629010215e97c10af7dc4e808b9e045a9c5175edcce9218baab190cd0975ca3d925ba29fa5c9b3edc6bd975deca619eafa0d53d80a38e6d44b586283894385f0ab172478f1641d9a1ba39f29ce759374a817b98844aece6717109fb6b9091454470e3c5601eb94e534952a38ee9cfe34102f29ff611cc34c072ab56f82885e925eb4dfddcfac552adb9fd2761c095846821b7ce1569b6c3d76c9f4a857c1534dc1406de075c64e56c8e8a16f7d3fd9cd34e0b124e272c6cc2c6f3f1fe6871d46493b1a9abcb7cd208cc779ad84a0123edf67fac470a3c85e0b2410012700c8c4687846c8313576f65a713c74832400157a5163131b04a1f345d5a1ef406347e63f7ef0e1a85063f62344b10852f2dd01c4bc1d917503e97994e86051cb777114680ab0938ac9a1828745815acc9fd2d9d8594f2177b985ac3253c8081a7a25bc5ec65903626596ebc7e0f6c7317a2accd79558a497bbf44c75e38f869c94c4260d9efaede849bdcc734eabf05853e74fb114c58e6bb56aa3711d86eac13034308420673576487d7d70d7dd35c4a0bed0b37e07776ffa771d7c0ba05eae4f551cbd64327f383cbba85ca36347f8b0d1d02b4efffa56f63a73f300a65f0926c8b1c3d49e049705a01b337642a42ac78451ea1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3ccdda613b47d1e99600f84b571d124b8c52554b53885d90592430e30916597458908655612834158877e312e3e99eb5cf7f653dae17bec797702972e47ae34e70159011b4014a9e27b5fd269dbcf81335fc4f95ac057c7e4979b18d77aa30886287e7a13b5e7ce232f02448cac319ac480feeadb50694685f1c4e235018272e40165db710b8a268fd269feeefb5c9942dab9ce78e61ebcd5709536f0ce4493845b9728c8563e4c2414ecff6e5f5e7ef9fcf24f964ef5829a68fc02db2add04646580bd270642db749217ef1836012ae52fea3a516de3fdb721adeaa804cfcaf60ac3913c39d38b6659122998abb0ecfab7c365330a5de5509c5be497517f76c104f5e02e35b78b2d9802b5193377902b3267820865fa03bf36b64913117eb876e118c1685d667124c0c6eaa593c287eb8f6d89b8dbee624d5d6622fc6b423828fc973e218fb6c92098d7e203929fb852c3bf3f8a0770fcac8c896e34cb3add3dff29752c71e32184ec729de0dfddbbe752441ff313c7edc2410d30f3e43aa764d7b6102cba29a758105e3b4c57fb985107198efd083d6388d97e992501b96194827592ad697d990a91bef97f2405aaab5a6b311be861cb8ed2f7757c49ceeaecfbf09a8a938c8ec3658f6dc94a0335840a89c4ec48c1aed5bcaac34ba76e689cd3a1e740afb51c3827d11a78f2db7d0035795be3a1216a8e1757dbde79b5929941889fd5fd7620cdde9de559ec72881b185401a59efa9ed6f6f47db93ea9d405dc017522b95c2219f2f9a1fa6b4a9ae777f0221c2f582675c4e8e0ab31a554176b893a234a68e271687573a2ffa9d37b50f96ca9c086ab3eb37ed605a4123c18c3bacdda74972a7deef0627549485ec1c59fca954004d6a28bb6291b4348c5622785482084106e49a103d6d01dcef261dbd211d2fdf2be7c460531ec6ae1d7dffe54aa9a0cd285bc5f9cef7b41bbc997f79d56e9f557157f77c179f55f4d44c691d47d4a4cd3c30b856738ed830d5de08412a1a7a44ad8f3057c7b3329981e1ed8d2aa5e9e93488f77b6967212fcd71ca33a1a32a62af7af372e5e3fdcce56aac5408a3cc7b6620cef1db715aa1bd7415cdcd6f50760dd809ad5c91372f01820c23ec3fe7eef5cb372daf6dc13805d9278af393b531b2c5c518f5e283d072decaa73e03fdc5063334d295bc23312f4790d8b8c111f9b63cec7dc09a67509f615aaaa87720e9b9507e18274e40e455a966ce1a3b19b00d7a67d48543058eaf202c30c4844c002deb200b539f9a42cca3e37cb70c3157619c0b2f645a1f3c995c8e58a23455dd3658631c612501012e7f4d40b2d41c0b86f155001ce6a8fac84b339cfb354b74de6b38c588015e625e302e4c5cdd8c8e67c7d38932c134f3fb461265eff15f89469618fe7c30595327caf0d3d741395347a575237e043898a376;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h2e59934ac133d6dd89b3ef030fa196ea05830b7c0b262bbbbe9f4ec71c44cf1f5d1ce4da60432baf0d99661979badb5100a1f87c7c90baca82c4eb6c221ad58369ae5a7a8ba5542bee94b3c0fc8cdaa9e55c659637a2cfd842af672593baf4766a90964a29b18411866d9e00b6814f4250bef6ddbc555fe852e7da24a12c38c7834d340dd4c2657ba57c58e9bb16a9202212a856a930dcdbf2d19a51e1d1047b3cb3da706022ebcc6f55253a2ed9cb098a97db5b585b19322d90efac15042d735993899dc59da073616ae98c01a6e00fd098f89f2fbcdb6455b585589b689faa440e18528e0f9320e66825c594526db504f541348d8ee13dd83cd931eee96bff8b7782168c23d8f8c941a35e8006b8e7236f2228309c9815217c1edda45f7209b72b613287f7eb24e6eeb6f904710663d7240351ba286c6dc125e6cb0855e191ba7df61024bb513d48c3cfdd687c2e8180341e227f88a2378ecb79bba611dba0ee5a0c4c71d37e7a7ea6df5358d00b3495fb5de8804e92a62b6577729565ae44dbbd49e03e335d6f387c0a97b43550d31f371873c2b73c5f0da292858564485957191c32e4e5013ca747a85880192b07ea5116b142d5d39a1f8bddfe3c7d4f792759d11ee3d4826bcd6b02b12c4fa439c4ad4640d439144e4f186504618746b909c2d0d8ca98e5afeca2c9084f7f94fc02019e98a0abb3caa60fa3f9521c506ee7a1f1d022281469295f5cc58caabc8f8793d18ba2ea9a7c5de1e570e129fd78c8fbd982616f084f9a84bfcb020144cc43bf7c9e4266c4d1a444d4ec7e6c592bfb5ab2fe8486a3956bd44a8847b6c6396a9a6a44a50e91c4fa43dc92d59a036cda17a21d6a4026862f60c4f9e4e912dd23538a788492cb7c79b7b4056935b9c63e3d2c55be6a4fd49f52c93ed6bf1bd0f5b145ee25b92b557a5aecef2fee3badde789fcebec8d115bbb7cf2f37f42beef09d80fa2f30d515504afa0db9c76840f3517be97834644d25e1b4a37e96bd187f0813184236315956e38afad6ad938b228c04a8bda185a5ae8242378e23761ce3364535fa8405f6f68c57074ad22eb20b9a5a08c03d98421a719117d2986efc565c29685c6c641f4a11feb093acaef44a2fd83455832db9574d0dadb4f9649de89eae2ad4f52bb455353a5a753ee17469d90e2fa1068573d369020b782281cb7b591823bb512bf619452eddc791e7783a5053b408f59b2017f0a4c785f6986ce91afbbf9ea5aace59508c5d95d6f2c91ae8274360a3cea01adfbc08deb60cfe90e320d3d6b05070be0bbd21b02aebb36e31334263236789b79e0aad1721beb54dc10dc9e4e40a40d4b73c5436760c4c9565fcc4ea93d7397f7f1d03ef206d01ae9f92b4b923e3b6d7d082b9ead46a911744f851df9fa4a087f7b553f8b7d1891f143f6ecd4cde6f0ab447ae43208104;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hcbbe83b3661a815d087c9b4f5b1aaf588bcdce8745bb054c6fff1cbfb3ad136a5ba80c24ada5bff125d6569c7d6ee6cd032446fdcb8f340526881ba28cbf83ebfd171a9a846ab87d936a36933325192c289772d27586aea7aff8c0c2e0a35cd1d6a6dc7d15d09861634c193863d4ee61921d30393be9c75802e42ded29eccbdc28952aa768af72ac4b62b08e08c6b80cc42d506c17f3607f7df6628d3dd974045e34cd236cb87c87599500d9b9d4cdfb06f8cfd0e7d0193f1dec1f4e7dded9aa6259710f18b98f7263adb50ea081c11e0abaca5adc07676470cf467ca02329cc7699e37ca27fafb72316c9dc18244d15e016bbe57bcab1faae8db272c6e77de3bdbed51852a2966d29c4a67b815fe98011e748ddcc0c65018878276238406951948dd28abea6b60c78a850b7697b39502885805941924b037ff02e18bbe2caf2d68bee0524673d6953cf444f90e388e82cc2a953ac0b77545b41bf6f41d641d8a0f869c31de2dc24d0f8c2533278549b69759f7b12b97971d186cba18e4099189b44ed12181c00fa1940d87f823d1a682dd4d1d68233c29fdbd3a909c6d4a8d744e582938e5c986ade1e9a4c3b65d3595ca694d7a763e638292b940d7164258e1dc34fdf675e9bdbc00969cc89929875c63eb97a6e3cd46c5002af4a282b7b2d13bf22b194fb8f3632bceaf9273a932ab9daab8a0689cece9762e008b08a4f03c8bdaa9e29c61afc0de750bd06a2d77a42c81fcdf6bd4efeb415bd6ce10daf28d63e7a3d5712605d4d4b0d83e8d554ae0c5a2cb0c356b93d26052c060085e70c6c74d24e634f575fc350905e3ab8b6f85c2de6b7d07fe2757c3c884efb91ecd10d38767cebf5a464b3982ba459518a7f4702dcfeaef45e307019bb6a218d83353c8096f258fa2125d750a7612131016dfbb82013eb61d0b700f2a9a79693a5f47518ace6c31e9699952ca374cfde1b63475ff2a7c36088b46680520ed6423064433496c236f64dad2d06ac4758101151d11ae0f4a5af928d200e65d74b28c31c40eacf6394eccacf234e2f41063f8930420e58369041e20a05db71569f65738517c0325b5bfb379d722724c326466dac25d649332fe613c656de1368071614dd944206b67ba49488a74cf2c91ecc0a0f71376e583429453566889e8957d7c771e0e055e5fe744a547c49bf7a92281fa7e96ac4341dff3712953d3f97dc5c19854f0ff04fcd9fc2168f45555d10bd17999e7e8312a25d85c75965869429d170b42629655af4ea3497d626b68b42f609647b85f07d75b77ef0f8162b782d8e6b8ffae507beafa33b90204dbde9ce9d4d0ebb0403f3fa5a00758fa2552aebdca83d8c22243bddfd1efb75ec0fcade02c2000bf0416b235ebb3911f08e6d0b5f49d5498ee9bb101524a16d2ff54fae19ad50a2f51ba8f8f0dac3e5e312348fd4e229;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he1da0cfc3656315a9c949065311a6facfd69b809d2dd7d050ed961c36b9ea46021672a45aba87fe5a13ad2225edda667402c929b34d4cdb521365fc35b09b07fc49623eac70bd8fe0b543ee92e78aaf1674feef986fca99a25895931a1cd7aa504d89a36f4b12d2f6f8a3198334a885bab52b3cd6286fd7d416d015311d11c5a0cafd8659e7372f105cf87f05c1d52f95fec6ce7a6e1cc59f3840588e0defc5ba41ac32fc6c949b9efe8dc1649c646ea99049e51dd52f7934020d987cf60ecc69ce94e6f40fb16bf8eeb210ffabe9d18d9602c8a3f3e99df202313fac0cab316a62ec6f1e3e4aef6a80597a2cca537e310cff897a06c0fbb065ef59fbcfeae71e592ab092bc582fce776f1d151650873450ef40968f2395809e8873ecc452a03cc01cdf5090eb8e96a241226bfd733912e4bdae44f5a795f2678513b1be533cf0c03e64ba181e11cd7aaafcbcc97b5c2950499d4db4fa928d9691d26ff1bfbf1cb484483996020b99fd631f6a5619a909cc0cbdf0eb57d4f2d6e53f52ba58ed81fe12cd6e18490ecfbac24beed7126bb4250e56127646dc0b5151e17e01e0ba45df8940831f1734d11bc6134564af0b93e0a88c5fd8faa64d92029e7d1080aa0e863e13a0d0f79a8cb6a3c5dc8430e6d103247e53ab1243f30a40a7304519137092b4d8bc3bf2e197031625d77d382600a040aca04508d5fdea0faa5e4a22e17e711bf8a1b0af78b9cbed78fc5cb6452f2f3c427b2c127bdf593d42a08d8c14b3339f67716e695fb3c3807c607347a3855e8be3bbe5f3082b65203a0abf428ce0566875d6b47634435710a414176eab095011c907f15252082c12fb99cc62e17c15dc3e669ad6d15b80daab037d29d8a23d875423298836fe70057bce2b5c26923bb953db7bcc565c0d7247fd9ac00c71ea75eca183e1476d38cbc8f38425454bb7cf24f39aa22fbc23e522cdc20b2b30afccf38fdc129e460478b2652594bd9cc0ce3c9aba886adbfac68f291d1bb86ab8db4d69a3e55d0e5e657664b53f28b5082d08af188870080b2e02e663b7c00f861db2aeb3b5957084c16256ab3bf488fe894d91d67f07b07f78c611725fbb29a2b9dc093c1507d439c0399719919412c71ae054f9514dbaf33cbe8c1f9ad7b9ce215887fa03094ae9406ca4521e247506fca866f4922e2547e2a23fedf087854b3e835d8ed4b3f856dad1ed039751a6ab83b2fe73b380fce251f269f644bf8e327cddf55a8b19415ec86a26373d979be0b32f08fae2e2574ad9f3b3511b56c3fa474fcd60f62ec1bb2432181286d7e808a368e5f708af105dadde14ea3e8e46eb62aa1325494a974a77b556fe130a2686b760e9f6d10499dcf11de66a6bef0c86ad6b1a122db8d48ba6f2122dbba511b4cf3d7806ac58e3ce9b8b883b4ec6b9b5716581541c3f0a85798c60ff1b8d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6e7866f9890e6d347fe33d71917a3d5a2cd433fc2c04ba38c544f5607ff9bb4c2a49c52e834a5da2e8a5e4c8869da4fde700dc6bb8f207969351d2d7f02fd345116517230d950b4e2a3ed83328e43169796258cd6cde876368e72f10497122867c2e679d1562744ce31af14274652d906132efc20c3f13dfe01da890d03c5dd7021963c5aaa516355c4e418b388478764a88c45cb1d00394d6554dafd7373b125d6e34e364494d153807401bdd46802629222f622abd311347e090eb54d44e5957d9e6515761bd05f468b23f857927e27ec95df06dae1d3eed1980a155952d28ca7d736b35b95d84cd802acc4e5e93c9c1f7e98d956efb84e7717719f2215da03f646944345d944e07880a6ed83d951b26ee76ff76799ca90ca2d35bc22ce4ae82aa083ef755cf3f1b4eb49919bdce81db692a8a6b2ec9d1e6d5d5c0a496e888d96f734ecb6212ae569a9c26014c5cc5023761ca7c67f57e76dc461a05169e3bdd797c0f0320b0e5a091530fdbdba0966bea23f1087049bc51d52e3f7768825a85b38a69a29724b20f40471a0254e43d4f601b74e013a9b15cc5c577e55eee1b53bd1ba39a41e7f8cf029dc288b73baca0563137688db75626badb6f96c33352e330163fea3d0084b35223879638476a1749837607e1fc17dc97759fc519a7d75611503c819bbf08556d094238f5b70eb530fce7ddb3f9021eca3a9261c29ebef0b40a2f4c6e69e26b03bc493752c5db2a509276626a38d972d1a61ea2df42acd785426f468317fa5b0be506f3bf89cba0c1e7732d4888b23354b669f5d3c510192d6c9da8cb09ac976d84538fe465361879cf3f41d460331bd9cc09313f0d45c1196d3ef15ae14ca5fbe459595fe4f1cc84c9d8a1596f0ab49ef44a951697574f85c4ba9b224730f5a59b014fc2b78aa89f38d70777508cf5e417f0cf5a2a6597f29aabde28f1c83d6b93a254f8148bc32f9ceccba6093bcd66725c02b73e46155ec61e95271d61b61e89ea2fc765ccf16c050c3dec1604a694b7cb77339f603da4e033371c9506794df211f5475a08c67109f8db4d22714a0eb8817982e592e442e95f2a7e345d4fac477e7f9b594764accb515b0e7b02438391408547b4b19905bf8b07bb9f7efbb06f77c545522f9c3ea80ebfe7d1423cf47990d118e90d0736baf7bbb32fd00edfb3ae36a6fd86fd962eea066fe6904e5f58abfb0f7006cb95a1228569c9bba604a3eb589cdb55c278872ea3eb3a89116ae446ad5f0bbba5f6218528b8959352d907b8548d6c7e4312d5b426cdfa6bd48b5309daf22282a2e72a00d62a3202a3211ee7ac7643ea432d3f4d44bd740ee042ab939c493784f441cd76f4dce803d5a6dac30eed05134f6ecf99ce430a4afe652d6495b6491b874cb423f749876334e9368cdcaa1a7682298fb8cf4133b5dc9d9f2a3c8a949e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf276edac1648596780dca0b01a35d88a066f90d8fceb7b053ee85df46d2e0bb54646a9ae3ab869127f6c52cb8052d64eb1f61100f8cef34942820e16e942d6717c3beb7479f553343a53560530135abbd5af656c862a7710902175c6757d57add01521431b2d97fe3ec6151ad637d3dd6fdb4f93ca376ec217e478cc22d5ad31061975fa700c72551c3ec1549ce3a4af0b6b16899cc3f21163e5fb2464988d5a9d88da246b8b01ebb9131ee87a744e8d5a6890c46393428fa27e7ffe7cd0f9022fcc0f27e87449effa2c0376344674e105213f431fe47ad40d8ce72eab6855d4ec79dcd50ad56d3805dbd1fbe1c1f9adc02e8b3ec6eba951da0ab35bbab0d261bd5f532e02bb671e627e77d8b2537f0c26e7e36e5ddd3cd0dd60f7d5390e05b6c2963c2b3b69c45fc54d1c706856cda616e51f5ca11d405eebc0ed4d47df50e220e5201fe92869b667747948f48d1bf2db0453e0c210baeb667b9b3fc43dfc44472a698f50dee67f74c2f816cf03dfec09068457852c56d95efbd61a57f7e031f1551218ddd57266d41c34bb90987c28fc1bb710ec637109446742bbd6c70c4766b96a2e7b13527a6f7a29de9efe8471a614301c5f455ca084e6b4e063a5fb5f8ebfaaafefb5aeae62d36c7deab49952084d57cd046314d07c8fa12e9ee8cd63c2975aa3b1700ad3a0d57a39d041f47ff206961a96ceee2c6004a5c1f7c907d2604125c3a1af9f1a0e51aeb4115ab617c67ff4b6e4b34e5f186de08710ea905eba28ea746bdad81b8b73e0fb88c29fbbd0ea6b2ece9889c9a5c98ca349ccc0504239b460d14e2c026422151c43e6c9b60c5973df7c3df84fa2aa5f1ff84947e8603628bc0484a08e35a849c575c162b15a678534614fd3ccbdf49bd624e0ef46014379d012db664974e2af39290e444e4067f5573e960dc627af9c55326c632aaaad402f9f57dc70681596aeaf641a9115ef61cb513f1f83a06e30ecd9fadb37735bf2e247a26b2a779a8a2f7baefa2c895e4426ea809cdc3f569bdcc202066eaca2e7ac3f2b0efb7366ba3f36c47e75f07d28da4b840c1df5e0bcb0a60d0dcb5cf58f974ba13297b7a336efac0b1801adff188b16f74837a0d3fc8e22e5001daf62b5878f1d9d7f9cc889796788944512aa9f0efba96cf5ccdcadc072bc014d755c0190cd994998d1783805686f49c280d3995582dbf0f4d1a89120e57acfeb66d3806dc3fe9fb04c467dca2b3f19d2db5f9d4d0afe3d06d75c3114a5f421dbb9cb5b8040440cc3fb9ba7eaa00f52c80d8526b4034533a7805420e2fe23130ee40bdb1dcb42bda5e693c308b5e532712e803488cbecb0e334e1e0f7a14f5650bbf19c83da194d20d68af996368ed227cd12289d83630aae83016dfe662668b22e2b8e14f1f4fd3d5798feacf7f0085b1088b58bdcf86911a90bc31cc75ef21f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h32f48491caee67cd85b3c3c45232fa08c0a9a2e95d7ac6f1263d0ed9c7663d47dd3f929de848844222af5ce54f2e145a05cc2bdedb2fa470f533f0da1c0cc2ed9a275687b7656da406e36f07118478b7cb72c70c84af936fbc062519730f6df4bcd7c6e3406eb1837c4de0123db1464fb0c46e802e61b1a055cadd55563a9e77b86d308d0ee0f06e9fa29c894bf6140389534c186170187378179e01cf5d4520dff69e454ba4d3b5a2159af4cfaa7af9e1d0d9e75e14f46803ec2eac3bd226347bd431303ac4388687a58656605c13dbc36cefd3366dc0154aac95ae24a7c8b17e2f48a6b474f86f48784e13046c96a91fa928097f311ef7fe918a4907d659f38ddd855b4fa9d695b1c8104d6f8ebc9c9429bf39d3b81afca3061c901b45dc9a5972f5a28f3abd386a9c88d60f7a289334ab6a5b529dd26fd6a6506e5ccfe990a33ebdb87babb12ec9fc650b689e2c44ecd5f5b2de81f7272bb0d90522e7e9f220edb5f38c9f928fd011b5f81e0f647bdb64b01376389724ecdb0c2276e367815c10cb4792c77f090e03a26e70de805eb6558a626af6dae5bd69e83f172cbcd2ee3834ee87d8b16b77c9fe4b21ffda85f58dec934d8545cb4be2c5118ed35bb90805280610afdf1e15afe1953ede712cf8b2c04acb9b3d4a06beb8fca8b70bd52b7bb2cf4beb5dfe66f0f320caf0cf58906e866a98183ceb8e9ee41ae8775763bf472393a1aeb043f6ea554c6d4bae45ac8a6568cb5734699c8516678f8dd1969ab7f7ff7391b8f2bbe6bdcc58d797624a2b76a0a3da490a8015839e6ce34d9380f5925a2d97b2f48d13f06df53a290b526f38ac20a0b88a4a593cdd884e491eb595734d16e824405580f1a3a3661d9f3db0ed3b13f25c64629e070dca8513fd128993975d4e0c0ec1b72e8591c8206f9404c3e9157a3def952570a04bae99aedbe0079c240aefa398018bc0ab5c3c55d5398954917f5ebf943f84235bcb43ee01e5c36324d2b95aaf1296867105bbedeb715941302ccebf5cb528d0f71c47ca2736ced4308cc95bbe130cb4abaca69239f7c70a128d691ef00133448f8d67670bb3eaf8016fbe88d5ebf47db9ef58aec885c2c51bd3a86b1b3d97d0ded6624e63b6f0aeaab9f8c56abf2f65f8ee9891fe7dfa9236d9a543e5a0b28a06fffb9b1378d6a6aaceb4db67ddc9a4688044c8044e765d1d8d5c28995d8e15be10ba3f4482d9643f85d17e9257b1e0472c992c6902aac20de7e6c4ff2d3b8dca3ccf078111a16beb6824d4e42d14cc622d7c9769e9090a2906da17b3b59672274369ea96859fc0e1c7ac6c1ef7f88fa852bf7d75f1872ac48a88df595edfc5c44b4d9566c8bce5e5e2f238ff7b0b1a66ea3371baca3f3af2ee69c57c1b943adcdcc22c9352b21029bb9ce980dba6466a7fcac9eb163de9b9734b07ad3fdc754c221613;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he86669d935624aa0d456ebdfedd40bc33233efe734082bb37f5589bd269e8af9321dc0d38f1dc90053f3e7abe0109876632bebdff60e7ebd6b911dad0e4d102da455a4ce88eb7733f967167131055aeb7b15a1829c08e4c1328731719055fb3bbf49804bebe2a32d0108fe6dc8c6532342fd55302d3170230a3e354c5986431a55a1b7c8ec64c0eb150e955eeccf327889ed0783fd6b45a8ff4ff36346a7bce727c0e510bc2065639fdb3a5f80d18b9802b4fe1be24e777a88a2b146437f7122514a970d14f169a1214b6d4727d36937ac1c28ba8d4e9c45798526781ebc9d7e26b3532c0010240da5168b9b74c467f402c2ed89bc16b619b05a81880420b3a9c7a5b2c275166bc29a7cf62f5476bf8454a7ec2b0b3f1a9a138d9c92c6dc617bd295922f9772b4882bbdc2281c013bfcf1879d73b7cde5c9597ba292f32a8bf27e0e7f722aafb28da6710c79f33710f979aa3a5336275b3ce794513fbff000f294e2ce9ee4686f668dfafcbf2ad4de7197eba23d64834b82fc210b5ace31a70f21f87ca55ee8d0fed5e84c8d3307c1e76b3d87e0b00d3eceee12d0bf5ed88b8f5833dd44970245ceac363ad6c0ddd26f3795550483d2ef52f81a233d23729e7cd293035f530d7b72d8a2d75fc5cb60b79f9a52447dd43c97a57dd150b1ae7df5bf01059374eabe6144eb3e5fea2735531193975c54e2478c48574558e63814e17f502761c783d551fa7b35b396213f0cf62dc330bf726bf1e801803cb8136fa88f29459eaf4f2860fa3fb62b6e22bce42ab76cde2113c9f521702456e5cd826eb9bede1f9ceb96d98229afc7f0975b261118c5ba6f635ee061d91c32b6a648608341a9b85af7124ee6e00cf15dd459acb3a39bb91ff4550f1eee5498a5b7a8c7015c5b9f73e20262cdb0028154dd9964ba15c99acc0f2cd6ef28f8c0f543776383442cbfefbcc5c7f959007877b5d93c66406eeef1d7874799861494589cfbf2dcf94bceee3b077e68598e0c796196b4e413e1ed0f98aee00b3603017f5fefcf615c248803cda63506ce1930bf167f7e10974e929a3f9a716c6cb2afaf685077e1a3172d475a6bae0679993894d1303b08c19b514c16c0682deb76cb01cbf87e2e62bb61fe1876e0dbcfa592dc557de65a6872895aed31e1a9ba7d0bd0934239ef7eb33185703a6d5df0619e0ca2430cca09a05ea70a8d1014a920de764b0c6f876143280d1da9000fb30b44ae545c58d1fbfcd0cd53c13fe323dd6f8ee8c59542374a91e99fac8f8b24389fb4532848579cb4e2a32bbe0f25858d144ec3700106853da6fbc4931471ab2cce276b2b58eebcf9010d83c9821084895221451dc621eece42417dc5add1c64ab7cce57f9da93151db2883c937b26cec9052f73aa7ca0d2df2bad7ac2e665d24559a5f275046e9414ced74d441fc69e221f158ae52;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h204ad6a04fd9660defba25a98f275ffecc30e19ee102f3ec8dea63bc10102a8e53668e24f23fbbd5daa8cbe2699113fad945a0d054d6bdbf05eca01c4e88ef2e6e8d15938bc9d48d02371017fdfea4edce6af6c7d4f3ed994f4f8ba15d20010f6680d56b4c28140559287a1eabc638701d749b1e1c32cd994d327bdaaabdf457a5865e921feed423325c426c9003c101cb70e9c39816321a44996939812c4388c12642406679068ea9bc1841249086e7b3d4fad87636c2a8999abc36b930c3be846e1ef84f5b8852276607ca05336c9a8b7ee7798bad235476760482dd729ea2a9a61e680b35141a0fe7dd3504e4de75bfe9e3a77246d63d7d04845d58763ec82ffd69d14b487a2f4e25fed69119a3a102c37bfd8defdf2f19bbb905e35e0652941da0027f920efc916768471d72265afbf83a81b86dba0bc49f9c52196b783db2c9b938cf4b09ac95fa15b73ab9db271183decffff4cbbb5d9e32fc0721114120d8ba6a6461d816c98808623c8d29a42b96517794a27e8f7e0e30a1e7e2110894b2362f92a098d79c28b1c6916930929a58044add5fde0b96fbd04de8d695eb7c8a64c476bc890fab505ce9f9153a7898c14c9637fcf3de5635bab18625366f2b61bdceda7d0954155303cc269d5e623a1f07aca3b5af92a61d216d6fba2a1e4cb8db80513f92908764efe3ecc337b8ca68354bb6ce81b0992e5626fb8083e96c6e368f77744874d64cfd48136d69c92dff08daab8d831c0a05eac519f384ed0a7e26618bc0f818fa86da8cfd5f46112d35294bb06803281be49b383753f6fdc78d2e2539288403a480b1e36c97e7b8eb248fd0079bf20accc7157f1478f0077cffe9fb4ddce8f3efc07ee38a3186bee9831e0d053a670976d69ea711b0a75535b61a56af72f4c56f73662c67aa93f93fcb0c49efa4e73bd0a7e8e2e3ea30a22f0a8d8e6ddc74394dada15d1bcec750f74b45fa696e958a91259eb0f57140ee71e86b667d81a97fc4816846846fa8d6c10f4b85819b49c4a92a86d273f926f222d29bdbbe3548838e0955d153b035ece6148733fe588b9269fd718661f946ad3993dec919c6a294d12324f56ac3f44c76e198103374703578d38c45ce3e6c08fdd52edf61578e8a1eb08759ff97d5526a8f3fc953451a744651b76b095919ffe878b47c1932b7b46e5240cbcea0b32def66354a1979bc709f78fd97a86877ea09acfb3121139e3f3e1fbe11a6609dca3110a98ff522341ea346a7a548e3d9ef903fa6184d000062426bead838a32ad4ab1eb5444b8d4c0dd91e254d3318b318f9fe4b9db74c86a3e2a06d0f6f7ebce0e641155896d3363484f4c164524c171738120b03e3ec150ab87eb700286aeadda1c35365b21129ecc92e2c85d05f3d6d4b4b41082f0cdd6be36e6a8769f3d0db43a27fb63096724d7c502ddd61ac5b7e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3a1204e5cff68ff904e879f32f940b4a6e2b8b4b292ced06d9e0e06cf0f991aa4293d0c6513a36cff588e5c74a803ba06064b95c970d460566bb9574d1b82dafcbe176fa026994c306bb27f120ce6919bc7e5d9065de208218ee168f12434c9ecd70ea62b6dbc6283c95ab15061f0d2afded8d0ef49b495534f1aa01f5ac55a72e19e8693826f8069f2ad2b56c45a323136f55e1f6e5a91d5296cf4e71232dd4f04757929b875ea399a742a66b60629921b5419ac665ac859e0e28fadd0108195e69a19b559f19aaf4097f696505732d7a7cf2173f7b570f607d4aa9dcf5266ac99b96ede89342a53acbd1adc503f185dd7fbf57f641e57e644228afed4b95425277ccc518ee3c43f5550fab07fecb34c8e05a0a82c3b8e2c37d3bb114ab104764f7ea3bb20f80f220780a8ebca0aa68c32842bf8a1784c97684d72bd8948b92df19c316961cc87b45802fcf27c4bea3421df91748e62ad01d1b99d29f53d8d4da6c7bb4119986822456fd6f3174b140f3b854e8740881f9559e92225c85259f683b5614881afaadc8c5a9f71e11c02db3129b392707f08394431e1fa1a59572917f849441a526f44cfa5d2279333e6662c204a79ccfc3fbac8aaf47f7c6dc679ade1050a276a12309061bc539619ae92c9aa0d9d3b1112c368cc52eb5cf92ac7e7ed533bffbe4939866cf8fdfbf3069ab0927920d5ea66109fced4c40421a3ac19eaa32492a29fa14e922c2d8d2ce9c4f5517b6923392fd4fe89a749d9ef34736bfd289efba3b6982bfef79db9233349a6a4a807f4620dfc636f5e3b69fbcd8f70b5bf22981a20c89c4eaaebdc67c8563ddef23d872f2f42714908a0d77825ab2d4ad3c133cd34da835e9c16f6b313806f690e79dacc33787b0038b4bf5e33489a0571942af3a59248ac6fec50caa3cdb0523c498fcf6f64a9fb51fb423f6879d1ba1036da3f12439156284d60911af941c9b4433ba621cebc4be979aacaf8ed8450f9c4b318ed79d06dfd1a14481543add0300510930c11cea13f857ada91e83b2db07b6fa8ffc4e5a0ef8878450cb98b32d77450bb8c2ba304f06574b1da534850a5080a2b6d176d42204ede74226b487d13b7c9774ca8e7f8257bfc6d0626a8644e231044b8730e990cccdeb7cd6f7e5b031eb8705dbe77290dd3d2b907eb8f5d7cc89e4529c58568d4a1431a93f56e96d795509dc4d0bc6f0ef026519a7daf880a9d90226e33d05e62597a9fe175eb028fb170aa83286948af1fe122b213db40f639b244a01e2de6d3896e1bf49b1dce948c4a160918974976c182ad04f2e4bb0e3893e85d2b3a7e92eaad7a9ebbf900cb140a11b0f73ba4d7ff632e2da312f26ecbcdb48de28f3a7b502802f5e874a546add0359af3cdca6c34cf2faab912d247176445e2540385c0c45d6ba38334f7fba9eba72a6467fe36d31682053;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha97d6e6f52de70c02d9aff7bc14ec70316fd6154a65e385021654833d8b7df7e587fba36b410c5766f690ad148e582e6ac69739685665873df9beb820977c967759c3834f9c10d5e2659a0a9ff50593d71d0ec31822afb8f599d09724a3d2be8e686bc82f6eeb06a22b42176f1c41af654263600708ea89981f6dd860b6fb5cb4f1ac80655bf65bec4bedb6ae84dcf1a7a672c445ddc3eff16d092d5efaf9778a75048e9863034a251adbb4c4b872af1a05baf5315aaa5aa87cf73384bcf7b0c5833ef67a00a7ed3cf17b792389172faccd5315bcb08508914d2fa4b1bbeb83e0cb34c1ca04211f0b181e74cc09e1eafc18eba570e7bfdbd13a8c82e2cd61c5a0f59cbcf3782ec432feae35c515d433c12d181279bd1b037525e0fce9f6d7f38fabcea5359cd1ad777b9a4a364c90dc214927179fdd83303cf08153c86c9d861d82ea743acbd94c33e5aff36c4597f171ed7ab454c07dfb08b815b67a76ad10123bd0e9f91d00cd21ed2669f30ec2bdd27a04be09e94fb5450a587281f937c5e5d376e22dafb9eae214c626793d83f6ea75022e90e330dcd824899bb65f4d317095603ceee38e438bce7dce9c3519bf460c3209e4b7c45d132c4778146c1f97dfe979f5ce84c817281613dbac197b7a91a3b80759b4116e4f05b49882c956eb93168dc5f9c2d84c904065e4dfda547d90ffe7b5cbcf25b0d4986eb0ce40d2315d3a9d5ff540c26ae4ca7d63cd304f6fbed467a63dcd5600593931530e796fc384274dd6a34cb0e3df48fc7ecaf5ffd9f3e6a8fc7c0eeb2f8924ad24212a12b36a16544cec5f141b6e501e129b5ed6ed1168230a19d774e092f4bdaef402b06fb46519b245a37094a2dc8bd4bf8d26e93a017969408b037c79e146113f15d405e25f116e3c719648c14b5528ff29368c500adc2e361dbd7a08d4f530ff8b729e5967deaaaceeac7ee980210d18a918bc6c40ea8e343029d8afbef36c8cd1d94a02ba44e08d78881543d01d5d5663591343d9c6d7861c11e8ef8efc1142a9f003090bdd53d6b1314b748f6233a37bf51c53e8ac4c0c6c0fcc1b8e4ec006433d07a979d68bedadf8cdc79b8cd5e8bdfd716269112cca020c3c66f1b59b5809093a768127cc058f31a58fc0a8c703fc2524b8203aa15ac7b2d1fc65fb3510b8e7c356edc6aa3a0dd8011d843734c2207052c3c74c9827c1f19ca12f533c012481ccdcc0f782fc1145621cdf9dfbab7b29e81f952561136fed75d5ff081b49d34d2b7d8c89c3a1ffbde52be856554b7790fd1ee371b6bb47029b570f8b5ed0fa2394512a53e0a77dff6cd5543fd3ff5edde480271754f8d3169d416c57dc87f397e2aa20b34f27a98d110fc76b7f888adc8039694ca91fecf1fb417659d5e68510e67c7ee9249a49c96b6c47fdf2deca1b5e5608fc27b93682b470f097ae0094ec997;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h592a5610e97697c40ebb0ce879a4e2cf6c1bc423ffb9037a3e4f96eb6519665dba32fe390201adc63799adc4e27652b09b1ed26488b9b60d937b1f243375e4aa379e5072442dda99bf5e0824650c080c8fd8f00d32e74b82c805fc868832dedc306e88cf973a48bd426ead1aba6a89b56daa26d2f353196c95395208e5ee2b3b81da11f8f930a066a534c6cde7c8e8ce06f0492342118e0f6dbd84aa8738fbdb395279a681c8a0443f1c1df991883c94860fc74b179e8f1f32c402766d54db2bb49fd23fd98bfc3b1848c774fbfadf06de8a1c994b92a4bce0aab0e4a0fa511bd0bfcfdffc2538065b2940ac2e2a656fe617118809119c94d8088dadd7de9a02d21343d8d7063cbfe869ebefeee588bdce18864ac355149d417e89723331f930ffd61a6222860e7f39f0e84ef8f87b8231156d96423ecfd99c0e7115a32e590d895f19bafde94bc5e25da69ecaf5122c38dd31edaa8dbe376530d84992796ea8952aa311063ea93786fd540e65b44e3d22643b008a060ae9cb9e49e1ce1981ba56738b970d432319692b5895df494dfbfe00f467e25d8f7e5f4d2402e6e4bfed1fee48edcd646a3dd40af73455e8cccc928bf2d9fc8b68730f827295ac80d2356ef848b8b0b09cc021512df24f13b056359d5bfad5bbdff6243ee975d7841c6958d9400aae805dde5645d5d4c37d2a232092d85bd60a1cb8edf1303899be2b59862908fefca40db54de0a9c3f3690eba3514de18f4af2d76b72fa04fc4e1af601e10650afa409ec130525e363c1da2a3a2f83ad4cfc80de8d4d3604594aad6ba4f92eac75da603eb4c5f89cfaa25bffbf57c14b07fa648927f5cb3f68fba50153dd553b72efd4ff5be64a66fdb08c8943a629de477874fb62ae0168e6cf8b7554b287ed7288c1aa328993ee8aae340f781d6830889a02cf9a8d95d9ceac16bcf93646b4ecce0ad2a1f0d7a5f6f7dae0303dcbf8dc06a5df51a6deb05081a65cca4be210363f1ca7997fa5e30689bf2cfc0a714007862971629425b801ba5a62f101153c17c8fc0f71bc0583fe73eb5d218143107caccdb273ba27dafe1c24fdff4f184b91afff349655f01f6e8ed9db98fbd7dd382876e14dc2fdef36f097088ea74246e9f602cfecfe3cf1e7d9aac2e7239a4eca5bdf42eb0457c971858e16ca91466ec7aec17ed6ab9f188bfcffe3fc976fd85555d8fa50beb9a6677ce746f3dec7b3a02412f50c4005b8b2e7ce644b924bf460afc8e81f442f39374b579f13ef3bc55bca9dd78ca858d7d0fae5315d5101b5453d24d419e96990708527c0e30bb7a57c3927df37a010e58ce96d1209e2e99589309b48f6e12a46a844b588832a6f67c1d3d6a708c039c61e26d5db0ce36b6cd10c27f065515fc85b723976a0acdfe6ce8851edcf1470b9071221bd4d5376db57689d0d2e9d9e2478845141a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h47e13f32a5b811fe7110cfb889bab5b0e3aeaaaf12d7b2e36fffd5d26676a9952e4e53b517debf996576e3580145c3c662094b06725ef0c6eb9abc8299e8aa366de3396b9ddfd117d8659b26323d1caa08eea93d1b134c3445889e4caabc2298162668182f33aa7a2c89dabf34cd3a942501946269e4b12432178d02c7b65da2aa217c311407110c462ee23bf6c3fddaef65f9130c3fd2d155f662b8218d1c75802803dea08645699f57c3ef6f708ca27356d201a8a08692343dcc86da35abd2f6434c7dd764c7c96c34c01b03bf6b1d324deb36c88a68ee28a8756c158dd9bd5790fb4da43de6a20da8eba87fcb5e46df7ff294a6c1dc684daf031ce8d9d06bc859699a4d1bbf85df5ad5d9499f1ef988706b1f9ba65bb8f3b4ddd23521bf2389255b35bd9d3cbcc56e2725f79dfd9c52c0d01b7536918f3dc30070f64f42d1d2eda58ff2d7c5fc66546f3195e11534dad61f6d82fc76c8f7bc08d235cc9f8067a750d9af63ff33d8be9c04f7d586fb90dec8cb1a2433d87173c4792b0d1b7e0c57725e6ea62af8384aacbba09d87ea371427d413b5614b71e0fa554712915f769659eaf5047bb27ae127c191893a9dd3c6d908dd04fe56989fa263412b11dd1176143897e55186b42eb96e0b5f74093f4d650fe40934732b894e8cfe1f555404bebdb72c0b99cbdc4d6e477af9a222956df703aa660cd8560ef2fe00b474daab48a0071bfdc908e6581292a45073f96ae75d5f4302383aa5975e4716d328885c75993f7d90776bbf2302b9268b5065463453c9ed675397210e1d21a60fe075f0eeda32277344452375904c9b3d657408d2d438e06c9ee4d34b0d8563bd57404203ee881c82b4f3342e82d8701e90f50f61c6329a4e2d83c7652046edef49613e5e082dd5986f5c8a84a8d45a7bdf64c373ead684ebcbb5c1a3f230f3d294f821824c117a9c29289d94d3dff5cc613d6709defd5cd2049c3e4d0e1ddbdfa9d37afd67a419bd36a0abd1d9f56b39e2620c7e13d0346650525b899e367b021649a9dd630a174753fd965e55714ebeab3ced298da0db51c37efee31a5499317f632643c63880d65eee05bff874f03da7155cc935dfa76a83e9a9314080b2a5dc95759b4fbb3135697a036865c07430fcae763a681f0391c522100e1ef1508e61023c37ec29a9cbb230a99f8523ffac84dace142f17f49b8142b19d6142b05c895f2c08a5516385e9ce3e80f183fd4905537eb5dbf85458549c7b49784fb28c244d450a76c28214348d376add764b4894149f6aa7061a18cd06d7f06f177997a3772128b602d2ec00e5a057cc7fa754636e513b7265f8b84406b2226895ea9e66c36de291b1d954c416c79685695357c50ada0b67393835d76d92479c674e194f4ef22783a27d21fea56f469ccbf03b7bd331fea739b36388710f4dbbb2ace006f1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbeb31276c62f789eda4017a09c18b26f0470ad714bc1c7ce1f93791be0a0e85370fd7688b2ffbff468db325590ecd24849fa695107a48bf6a7bacebf7111851ae23aeb759671f7bab4f81ca732576fd9074f081cae1d22f89661fc31b2e5bdffccd73468d4b88b9bf14417375edd429c0084f0e92ade842525f49865911bd82a0cbacb5f8d576273b9e874bf08f4a03ae8430bb5715080791030ca13c80bc55b5af66e8cd84e5e9d402826b30c49a4eb4c2bf282541a75786987879081dc17e084f4c5a0b4023ebe547f05a5a688701cbe695dbd551663dc7d0b237d5b659b9105e806a69fc9c3007b2c5696d221fddec109fa4c631faf467b8ae7b5648f0e13d6e8a93dfc2db967721f4861e17c31de8c8069ae60049539ca60283134d20f619385c5dc877dea49914ade2cce9165bca4f5725e49aeb193806332bb742eb41a8fca3c671638f35601c2408b59f9d130101afc3ba18070aec8be6fc7c8638ae2f6cbaa23f652f4dce03ecd289d9dc106315450312474f1fa173c57e70dfabe4575a66186c2dcb5ead9bf8518b281aaacb6859db5c391ebd56a4bfa08183fd3715909248c8a60dee46e1f5babeec0bd12a34e157a22a29726b0859f38f2a339efb44d1028ba1a794b183e7df0469a132cbf9cf773a599117b52029d06b0723eb606e0ca09604cd4ccd821e179ad6a4c3e277592b335a675f1e68d38ea09e0adc9c260be1ee34fb16971483b4734eed5fe04393c7c24a92e412be894e03fb75bbe59575f379f01bddf91853c494f353175b8f02546e0bf275164c5bad336d0e9b74ecbe826c40252cfa137f9548df1c27a3f8c04c0cfe573b9bc939fb8ff15cafab1d9b2ac6f375b9ef6dcda4c238c2a67bc47c380b605c3b56d81864724757ae52d90da2936172197f0b35ee91ad8b09e843c0be63b976b7687bdc409e76f24c0ff58686d5b32742099c005454f5d857f81bb854dab21b859e253b2c9514071306fd8843bae7ae675be771f95ab207179825c08e1f9fedff173dfc18757a003e6d09ba95e6ee0c12d155e2e451899ef90f12496a8aa036017aeec147f2be3c3500df9f17be0786a4b36184ebb9117a54aa2927bd7890835a31cd82de2dbde284e60670495a18472541b8724dd9a62d514918d7adda61644f5163d8d2eb5d37bb29fe86cab789dbb3d9d74f4ffb7da5833f27aae2ef47279d1b9335e63500fec99d28154756490a33259ee78e8a66f47a561825a1c47d79f23fa897dac0f772535a5d8de310afbf65552e1cbf240ed27408dfcfad9752f25b175a2354b33ae14b93118222bbc5131ebfc534161d2ae8f503214f373be2b732d470294e4cdef6eeb21af531631ac8e0d802a39e25d6e49f45d8211e4a47f86d4e8db45895bbff62786a3794ac342bd00ead56254068a6ed8fdbc26180f1af38ce223a82dab90be44;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hef7c9546b808659eecaed848cdf74c4738b9cb70733c9eb7065d113eb1333039f393f02663011f714ab0f55fc9cb27e3a2eceb9b74aa657605047c28f1c5f3161af33f480ec9e805fa4b2c1c3ea75d3b1ac6ca7d29a5a749b537bf9073115fd355183e5caf5406cd772a68877f61356f726d03dd0c33d3efa824528919567251752320a0242620e5724f23b92b54897b5515593ef2d19ac5b06dfe9eb780d51a7148f6d2832fb8af5bb3634ac84e88d9ffbbdde85272981b0a80713e5b21f1c5c945b1a322e4ebbc39f99d86d12f6045235ea0006b400ea1e3c578502a3e4a9bbe47ad336c3a03057935059c2d30eef3f85176f0f74b53237d7b1badb2a6402739dd41b34460a30144ddb667a822e295dc91baae3f841a4c6c11718ef01bfb8bdf03e676fe4e6e351a04821197ec76f290dcce0e17a3929e9e1640ae5481ef5b91296195aade82e89b82a48abedfa10f3a33a354406c61e60b891a4e5288fd8db8910b1009e52a41f58747080bb5d0f4ff0f9662efc1550e5dfab84a974ee7540ab5988c4c6eafbc01009c3de1dc34e67af38a90068e72f8f7951f36cd5527721c28b5e1af812ee14741474f1aae387a60a80001508183e170102e967a1b06f94e6d5f78dcda8b81b71e6708c6dd9130b98426d5be41a6276ced5b98201664b7c9a99f7357148d8180d270407fde716c03d56f566d6339c73da605d2d7b87993aa32fdeddeee6811af35c34affb7cb950d2712a68ad049dadc2185f1b0623ce8f9a6ebf163ca72c6e3dd74c315deaea03c51cd190aab67887f081d6d85110fa44bdf17688923ea3c5de737a42f3c46ef694c1c485358500ee5cef3350c4042de45dc78c4d01c98bda1ef551b695b4dd3620e51395ceada187d98c04d855d67493c2d44ba59a3270cfcb3dfd87c2681b000551f0f21f55578c098dd58e9ee09a097ec30b9023c498c13b3ab07adb3f4e3ec0d22efd185b0e3993a47ae5deb2b94a5959e22d39cfb33e31b628a7f791265730d02f9bf4b9df4d741ee41800e97eae8fdfc10afc6356b00ce000cdd0b766f951f7fb88cb68b84c0e874d5d0f89118ef8e5d61f1a607bbec2954a4db6ffd2940f20e1af3a11345a5e66f8b1a467b07dfdfbde9e260d8ee0327d599bf484d22c3dce61bddb24ee6381c50b86a92c775d07b2f03ee16ce6878002c0ad26c646256519b78f706c5ca92add0b318fd1b7ec08d18989f7b410187d344feb51e02b078645d6b5ffe7bb795811a8629792d9228cdfe744c49b47a866f58b8192f761e42bddb0bd3d8586765b04ff64840118f13a96161177ec3453bad68e5bab09c73ef5051bd7211282bd854607b9f8877b4782b704404ddb1df5f52246a617576cb3155fdf7dceecd3d35e70404ad9021fd87fcf5121b3cd1fb041713b9e28711ae94ba1eb65b5e11f3b3501e3f1918d4ce;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h2d543ecaf53d72189def6f68f5edbce6af839f83a49220d25b6b104236e9db090637fe9dc7e399dcc1fd437fd771bf57a55c0fde378d2e7d6181d67ba6ad4ee08943baf62fce15552ac3c7b4edee4182528d285c5c9d5c656d0978a8857f05aef8ffc56dcf17a59a7695a8e1080d7632706082c3f3b2af246c128b8b9d86b79c97f75346009e185d7310d897474bec22bcc84c5f0dd7e1c856f009f80f2ca5d46802eb83089811a9bfc0c138221e16166a0186c33c782f92e7ae2fee2488f544ce9a6c5290517db5c0a1450d7ac54f539f1b515521e7ae9c5ce00184a3cfe4b50149691b3c34a844eaeb2b05f700fef12e25be674459224f4310f67523870c1f1605eeb25eb031ac847696afb360c045868fd8c621ec26054f73d35d525d7067e3bde71d086b9f0b42fa3ead62a34a633cc7b26c408bb2f13a0fb35876b4e879baf81e650c30923771d4904b2922f45b958b9d3765aba936a29ef9619f7c28160610449b7c68c2a5aa77a70709a459c0d858a70fcb21240ac459fc7e423e85f75ea09cb9b35f5e80cfda26434d902cf32710c8670ac15f6b1c6643220711e633d3ebdc988754bdda0a7843de2ca4db69ed1c9ea7d5bd9644112bbfcd1be02404f0a7bfdefc93f271064a8e07bb1df3012ab2696020d8d5c3d0e03f19aac340426188e45e47ef4c2498229d26e54b30bbbaebfc7e1d068458eb4ff7cb86244fd5f789ae846f9ab0080848a5404225983ff42ae9a2c06969f4802a2cddc707e2efc0e608d21d031f78fad715d662a5ed0003360cf89c6c88d9bd70d1cbdecac25d55012da941e985bd0ce983ad58c03f5c74516a36550cfdfa3041ec02e58b8a78e29fb37c1528f353d0d09ee952d8da1574aa8330419c6aa5a93f3c7bda8fb40190834216476a96f55391fe75829439fb8c088fe7b1aa51328f2d406949a6c0a170bd100beba8e2c30e2f300a839795974efb348ee6e680223b810e7f92292aff298b9f15729576c90943f04197c0bb1f4b6cd65da1fbc338dcdf292182be9fc5c327fa83df9ca6e9c02f75144751ba47027df1b411f71a8fa6c5f78980723a4551a2f0d3265c3b1baaa2e7a7fb0c4201ce907351e1cefae9a7e1da1561217ae0b07f4b2e1f7c79363e7e77f010133df2e2192209069bd0fa44157a96673b40336fc97170caa331ec47d22362b19f5a61aab35dfb2a2fccc50cc7e1124c894edbb6f5348d2bdede776e9113f96242a94c2f59ff6b1664114a97882edf3c467d2f49535d7ea951b98b732d26c894d2d2a9888b7ef4eac9bce966a8448df410cd0462b113741da1890bd10bbbd035ad9c73ccc3de793266a90827d05628407d3ac9f964169543295fed847c6bd88cdefe33f9d07f8f1ae143c1d924849f0981c8ea6db4bb52a7d4b8da3f6b9097ae8b8ecf6f16b2bffdf7b95a63e44d4f5308fec4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hdab4223406f59bdbd5f55a23d11a8245f7eb34cebe5a7e57adc17d45042fe37473c8755e61b18dfbcce62b689663e29ddc9a9537187a7d61b4df2053d7dd198021db43e4766d9ab55e5d27efa6879f16d70ca3206e80da8cacc7046d08373cba7d8ea7a9d9b36c5f12c95173fd08ddaeb88590ef49e0fd6cecb624314cc459e6bf62de6f15a73411a0fe0735777be2bff3fda7062482d5002cc736bfa2b078fdf18cde4d3ec7db27162a26359980ebf25a22b1b10d0abed88f4a71016e142fbadf6d1ee1a7fde98014c879fced73f461cb365660e90775b05f4eb196b68cd98a3f2cb53225a8e7fdd589061907a1ebb05afa622b59fb1c1ceb4dce585f4c7428a0e26af26e89f22ad719372911cc9a6684345001122687923ef6736edb10e972d658553334dbc3317fd988f3d13cfd4089d7019d903c7f54620fe0f9139c9046f915560810a32fd22eeff7f783c0c248a9d26ff30f9ecd66195351445bf11b7bfecfaef47be63742c0a25e1ad8153342d29a1b73068c3c20de49592371a9abc5504e5cacb7529748f5ca077288e5371ef1b87cd76d5bc72331a9d90e229fd8b701299fdebf92251c35693263e2f49e32bd8bf19743a0c472a858da82bd98ec5746da80b39dd9584f324453f30afda8e78876c4608670a83f07a1fa7131c487333ec358ca8833404e7172c76483af9e0f208f4e86952be917fe91545e95709fbed43741b5b80a3650cce278e8317a145042f4812bc5711cd49edfeb682c2159fea1f23c56e2e4987b3c55a944dbe065eecd498a80ccadad30c0c32e2d0535fbc1a07a7392d094f71a079522f2c37a8089ea6e89704b897ab499de6ed2f81d784695cb62be097cb61a875cd4db9925dfe3c6f3e8c5faf64d86d5d88603295cedc9fe61a851ff028aa94d249a5e4145a7a2c86c8e2852b27c4cbde33033564d6bae19ce4356c0ba9df275cae7b332a194b8e50ed1b1003b272317ee1dc4bdb4feebaa265e1bffd8b2e0d63f39b4064cb7138f8236a929573f5b5d12eff6204ddb0a0ca5b06adf2d71071e2f3c158599fe6f9faae09961fbb6b111d64393544580077364c4238bbc7f3af37f7be7512255dc9911dd04f13dc94935094ed90f4826bd99f4a4da11302338cc794c98bf6d3b40ccd58ed06e8190b6079faf6dad398e99cb836eb0e05cccc309035884d0ea1438238e911e3d736172f801a06ed2ec0262ad2a8be086418915dc6e0b077320410a8e49d52ef800d896b9f1f554a514d435a83aef1f79a03c4bec9df0e5fe6d54978b9135c997ac2199feb6d87adc50e3f0e17e065fdd97ded26215bc7c85a4b741e9014b8d3eef09f24ae946b652af38f13ad7562bf5cdac03e930f666972fbd4fa06db5018d4cdb911f592a834fb08be91e1e08a1cdbf5b5725c1faadefc2c33c1103a5d96fdbd5671036c2e5b0116591;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7c7a89e1f2508261eb307ec1612a7b24efe69324ea969ed939c921675d9101853942eb23154e35c4963215a16f0910b5bae6e7f8e5ea3bcbe8f22ac22f83023f95382fce3d32349a8d626861aa4fdf9a2948f6640240b3dfe076a38c4bcc4699c64ef96633ca65ef19df235217be9aa0d24df896b59c9c34b9fb908329d176b0a257d13da9661455b863313afdde8c28651d06a6cc4d3767e32bf7fd865bba32cff25d8ad52cf3bf4b9e528aea766fe94778cb62b87b16dfe2f23d472890b9f75dbfec637993d0bf7e02761103e5500703c0c3bb53260de5b54d67c70b51495ae910bde4b63533a9f5b4220fc9b7cd46c7cce828af9e66b9ea4bba4ae9c639dd75a5251820f5d4384560f76a6e02cea928e90e5f62107e5a7adcf82ee371235e07a8a145da8fc7759dce4e2dcdc76c5a3374c967f29db4c5c394eeaa2f772f4f1082e2614b27ce74b55346f68f150431a87ae7a4f28f6b707d824f7e9c204f87ecbb9b4dbfda912d4c9e18d0ad7c70a5a0599348b1a603f9b9b2bb3b17fd4c392c7728dbc32d5037ef97c76a2c25636bca8ff471594f591053ec0d1a1c33d3f5fd0396feff07bb0167027a1ba9681fe14e7afbc18fcc3fbd0687ce570a18c3f1d3ab0f2b84bc7f4294a22be5e08465f19f2e171da014e533b97502bf35635f0c145c75c6c65d2f6d2eb2a8a9dc417417082b5d7468daa09cfe9ce2b83b8de697ae70c604346878e25bc1adb954fe6c376077f0e58a66ab721eff62891df4f40b6bdb275fa72cebc4374be1da6ddb3a5bca185cf5054fab852ac963e139fc03adb28bea467adac98da39eda46efcc2f5b01682a779446b6b844eedf7e2fd0be98cfe300f2207fe33725a424874692644694b86313305e471d4d8b254d875c932b18d0c3c265cdd2cdfdbb1c935c3712c9e718299a4124e70b5ed7fa5d55cbc017c2b1b7129dad328cbe9ac3cc4225a82c00ac144b800bb11d080d2224e063ef4319eba75257839ae6a991377d2a3b08029db90740cc9a9be2081ae834dacdef3e0a1560c81265110a84fd95ca474982ce40d429bd0cfce632b5fa1648dd10ed5578379ead93ea651605b22bcb1914a3b0af3067060af5b66d990d9655add548eb399749a61497e115a0b7124f297ea38cb12cfe774ef21a862fadf9dcd72a110c744e78226113a56119a0a8c0999314c62ddcd4bb06d0664b495f29bd063c5dd0b1f8a594031efdd93050a4218d084d97c4cdfd100ea4dc72a08eb169ba892db165937bbf8cb91b868395c7dbf1f4d3910de1897cd510786375deeac7db9bd65f514c976428d6d1abc6a5a3fe74fc8ac8dd92e6f99452403783c16667d5ee7c144b0cc5070169dcd7f10140be1a05c141551c4a6f64117e009e2cc67986ded783a4409d611b7739f472f983f70d1b533ff3d9e195deea315bae42c252fe2a4072;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h2b9310c974257d48e3574c6a95ee104b52ced6c8a7e4a9a366c05a009c27dfc0d7b63eac79fdf71e8f1aba5b52bff031e7f8f464154245580680ca80bce76fe9e3bdf0b8f7d15cfb2cf1391e5240c6087b3f37ab4f31c0c2f95a0d3a1ddbdd2f482a378c669e4a6dca71bdcbd49387ee6c71984d7d1acc67540a4de102cd6610c1fb4cdb0d10dc8376b78f54a3c7b0fd8b2275a154f8d3678e81b7b01e53d38d0be69ba81b7554ebc639249d95e65c2992dc62d877b029786413b81bac422e3a5970175ce6f5ecdce71c8d144e2ec470efba85305aa549928c0a00306ac6c74cb3a7d43263cd17b6929bef8dba650fabff74f9fd84ead1bb3957d2edc7ac125947812892e112fb6949b79d1d2c6993459163bf5280781d49e7b1cf59447cc3819940a8504404bf11df889d1452183fb30312e856f11730914d378acbfaebbd5cdd8e763916f99194061d25b4da4a42d2763207da7eb60114b7da5e82d2f0cb28bad7d0a8445e6013014d68c55c142902b473fdae915f87eddd6b37c9a90f3534996cc5f08500f564fb3893dd3b1b5f9284956e334a0f61bc92d927ab66948921842d84e841153862c19277d1c6806842135dad3b191cd7422bf2fac3a8d80fcd673674319d5c592eb536a7884c8eeb15c55fb47cf141e2fd2d4d84161a5332db126cb28bb66e2a83b7667b5686b62bf1ab0b1cf67b5a8067c347a474dd84f58822d426bdecd08839be30d2cc062b1b2e3ef73d8662e6f84f87d38128714ac4a7bf7a3e1a2edce355d3d3be24b464c889bc34f57842e85ca7b7ccdc04c463a5ae992a325580f4e52fe42ba022b4da292ffd92a0422beee66b7f3da7dd063bd1612b1287c7926f1e25af1ac0f392279943c4cdcdcf3d9ab7280695df6ad0cd0034079dccfe441406e1922f6a71a17358a6f70dc5f8ef66c842569cb89101005d4f969131c1d67843eb99133a414eaed6552a1013122e8d7d4996dc7e078c394e67764bed0e1f9c0f21b693a544af781bd929cca19f2d12352015646382c8fb35382686bb5435553d1a037aebfa5729b22b1cf80dc5ec72cf847c606873a2a6d81835762564239decf2f590f89fe7b2b53f3b4c5e5abe787b34d2e2be8033596aa294abcfbea0fadcdb5c91be18ef25f60f895d24e9d634a4c21f4f100cf2d32d6316cb2084328f8096b91d0aba162d8a1b7872144748ffa4745498cfbe5f7f60e516054011ce7ba66a24c14c6b8d614d0d89879d8e942390a8f3b93276dd60330ee09c290f5d5c73f927b2eac3b13e29c55fa9edd066a9a527730631184b9bc6eb8f8960d7faac27f3feda3fdd4954e7461daa95b327a1f916f13221b33737a6e3503db18cc8e1395bbab2490aa79d412c3ff065bcd99f383685e93467902f4b932e7ca03c7eb7504506f9c6d226d33007b8ab57b2dd61497d0bdc66a9d7192319;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5717ce5229575230d7f50fcfa086a24c4f2ed6da29b608f6b4921956b0865f7ac97534ce856032de8f5408bbc0c53eacf2276bfcae43060680e8d84eaa0bfe96c2a2923f42ebc84489416a1ce93fbc2f238f442788b68e0c4cfc067ca75303fdc9c520a56a06e3f6a51e1395eb26dfd6d80e022ffb488ec89f564c3694837e433498ba9701fe6253885dc7f89d85722383bc9f0b3e426819f179763ec638da926b48d2419a6c33cbe8fb25324f11abb308297485a4fb468b0cdae5dd1876b58e340bda4d69eb18d4f156683185baacd0a8424d470c7f4bd2d4a0af286b74bbd432ef2841033a209636ceb35726d5d5a09a16108f73f0dd6f73fab50de32aee169f94eb99593877272df8da63b61f183879680e07ac8e9c96fa9cb3b2178ed90f9cfa72de953b01957c687dfcdb4b4fca59cd070091b8b26d78129940dc8c90bc37ba42320652269ca4b3613a50256d469b27d84182c706c11fc59e7f26fd62018b679df76538551db0a674d382ee1b7d4e9bcbcb64703173a4645226d98b3f98bf075b9f82b9f29319a92f0af51beee62e9995cc18c849463c07277535aaa46156750d249e2802d56fbfe22b925e1634772f33ebe018f5ff1a8916d05fa3362ff393a3cf707bc25776bc484202adaa63d44f7a5b1bbee3194efd8ef331e65128e362539fa008243e52ac307615648035d45ce924dbb2d0e4252b4e011a29e221c5cbf08c6b7648f169aa32f1ccee4f7c0e75b1e368f61dba50e5835648390fa306f0e279419e6a62f024e85fcafc5849e04e9b1d306c6deb113d8099f017c1c09682dccbb39bae9870ce080d97dda5c5202204bbe4744f684c6a7305b32243e747120665b35869b4746f0cac8dba2eefbf02b51c625912bd5ecbdda5b4036676757621b408e5c0cc01730798355fe9c79a75a3015e2ca715a7d2a4a5d75b47f0ca08cbc9c235fd7a6c89c8dfd7c99e134a7c9a528f9633d4685cf5dae6d0c2c1f5b1b64f73ffe1c661e84562d2ba8215ad0bd2cd8d0bedab06e94ba8de7d214edd21de84119bf3dfc6b7470a67b3d03920bbfc5a4fc1acc400440137e02d8d1c1b03dd2d78ece2e1d10f470c8b62dc6afb67fa20cd80488b3cb9be8a8de7c0f3759b10067c294a2b1a0e4a16e1d95f92eedb9e9fe9bf045d5e44657542a58f3a2e23bb453bff989e157d5adf3b48586069a8dcc96435040032d514904d6bf4884b1f42915fd363b3c315987bc02ffc9b62fd364392bb8c3d5e465e87de2bc183dc66fcbfec09be29c5ed3f156637fbee349c1136ebc26ad3cf7fd153a8d2e56280fd5617799e2c88a24103a1eac04b3117752fba2bf85084b0f48479e3c830f35b5eba053440f14876c1fdc9c3fd869e235a322d825b0f9bd4825a7e74acf12736d54a4e719b701b0a5be9c991a667f5b5ef9abc81ec0304f4e9493f1a13e17e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbb3a27ec09d065e8111c0e0134fa3b257f90a23a5449c187a74ad5a08dd61c3f5a97d258552847b1772fb59097979308d1fe5df2cc6e97957ce03e2e8b559e3c111765193d7f2a431f2942168af23ecb5529fd2525b0bd0405ea37b64cc65e87f996df80553cf74d182f3c2ca9b9ed40635d3d64aabf81a8b629e0d5e96a3245c811de3174a26737abca08381c69ff07a90bed709eae052d8684017ee4d5f9e9fcba93418faa20b73ae3a87a5e301c5bfab7a34f4229dc44786b12e88b15ec0c29f0dade9fb18a6256b8e2a9fa5e107aad5099ac61a2a9bc4a98848f88e60b9310eed6ad94980e6baec550da8286f680706771805f91e3c587955c622189030527e4baaadc5af6c535a27c78dae28c7fa0cc57b0c2e327d424adf87bd10ed8ac856eed2c6d4051c3600279c560353382c0217f04f078b31f2b97561a6df9006d9aeb2c921acac879b68d3eec31c5a9a9e6dca1b4b8e0b10c2467aa03303bd11b7e92a3951f0a92cbff3872b7702a0dd30f811c68dfdaadfd044d5a0c1febc84c960c18b029c234a9127b1ca167b1a40ba1644e165d2d4499e7facfd6894be22d48ef9b38f7090d9620313b2b0301854277b22d5265a86898889a3ad94dc5670728a525a67dc7c5721145383b908142c42d0289193052aab41f9f0fc56c0d7384a56e7beef65491b68068e678ab261b35c8abc4f0bf3e1ec072c176a757e89aebb7ab143cc9fa67a8647ece2b8b9eff929dba2722bc8509307c5e764244c2114f0fee4957e3bfe582529ee94b1b6cd6338a70ed1a4b715ce4cb1c7df5c6803725ef982d103d81574e64a6c8cedc36fc60faf79e2b86ec4b8e4dab3d6e311a2980dfd45d84c8c8444c4d146a6ce4c2a195f3b264ccbdd714dd461642f4c3dbba5dbc109f69e6c8ef32c98b2121701b3bf989b1d299badc7144722cb9458777ca2ea6e61cf9b47b83a81697720684141d3e5102561a7e77c3b8bee843ac267dc8d4441fbd159931026c9797c71f0889f9e04a5c84397fa708873d6bb008b7fa728709c73e88a4347b84055befaa78da3b10b84d1c10cf6e68202f5ccf463061ff8de51634700c500940445819e3fbba08e3b4fda547319b53b541c16575fc743cb2449a08a6657337181cefc626436846d3008eb54017fff6727e67f48931f5f38a518f03578841eef187bbe7b48e4891135b07a5479fad74cecf0cb71d96d7001e0a6c95a0c0dc9f244ee32aae266add123f5d293a66833cab156c81f50dca822cb330e52e80f0e628efc56114bc0afaabd3c406b21c8b961062ce65564aa77942acce7ecd636540799f81b2ff322c2e608322119869df19cb3b1a326ac4daca7e3fb354ac0aabe6db96550f66e93c180be7ca0ab57ffb2316c2923bd79878f6b7f30d73429544b7cf0969fa311920aa56d548323e391545581eb5b9615ae6aab2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6301e6fc1363e929e0ae559f1f226d0807cf2b7ae23a7e3cee05d150adfea2a6d728a16cb472c3942ae055eb7ba2a3e5ec277f3074dbe7035edfe0c09d9612f5d1afe2fe7ccb8717d85bafafc463a2730da4939f8b2c17fd650e67371399ca22b9340dddd5ae441a6529e41db18020a1aba2fca1a3f3406853044ce058365096a4615754c2235b9d0b30dbced4efa9c0b34a39341b56c4d2f82ac4c0bccfa149b9d83ff84af5936a50678e46a346f14d7d912db144963027e076af5500639fef8decbfcae1b680d1095e6824b36b53757e705be8da66c96458aad65f34f454ef6aa347c38f62876505fb266006e4c3a119c1fd725b3a470db75a59b56cfb3a2ada90e38ab9c1cd1b8c3493a54b95f8b9ba1a69bb5bd0836b231e2b871b10c731e1bedd82321460b2fe6737422d5525d2cedde82690dc66723efbbca49f9997d2962991aae68438bc78a8685672d2c83a23922f63171859305d286ae4be21d73bf512534d753861eee33f06bce5cce912e1c5dfd67045b6e635b6d5f2c67c181c0a227dc6d6890bfdc6eff4caff7d5315971120069142b8eebfd82f00b0d7eb61a272ea848df6c8f30226b4bbd4f56e3a69ae482ac1e7a3c64cc23ce9d6bad8666ca2e4de30c0b7ccdea8fe41dced1fcec8dcd572a0f99c342b7de35c66ee82e024fd71faf59da50d4920402a382ca450382626b102a501a87a5220e181f4d660591ddb5a4145f94d243526894bd1cc7be5c8e9ed1688ad19c294be8410e737ced1888f3a42bd5b7ca7044b80f007ec04308da88cee559bd5e4e9a97355035e6c4573479cc2c698f9019a77ec064ecc22d13de98465e5e6033fa5d3d892ec9952d8bbc80c6914e39e32ee51aa1f527cd7fa82fc9a2a7525bdbb304b79c8ad48e0410c84b68c82e150bca7d21734bfee2685b51f95a5671c0629a3afe65c37fed9f724385af6c01866bdfec69fe13c710211930606fb82baf263976119171d3a67ddd6fc0e335d0d7eb794eca00a0bea5dd6e712428d49e1ff690bffa369b55054b82ab3fad0269aa6402eb2cc541f26685ccc92abda52ea251dadc9dd9ac7ef729a32649e94906dc7f8c538734d030a38a63a68d42a9f32513eb00cc0bf877c51892f3e592829fd31388a7f53aa3290e110cbdb1b7e9e7f098bc1f5c4835e2120625c427c115ef1faa8d6bb1a26d14c3fd66124a2ed8b1da7fa43ccca247011ca1377af9bd890d55a5cb58a3777efb1f4771ac45b57d42d70e2f139fb2e5a3ee63f606b5217997bc140a3328dcb2e5dc7b55e04503f8610a788844baf055933573fd2cff31af3b356ca541b698591ce9205e0b6286c022499c2377cd333e8e35b0608554f0366471904982e12dc764d86f47be0b97806713928417010d7b4fa70e639ff6b5c667a9752cdcb5196f5642c3599e8b45a9dd60f994bf38ce1d679ca;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc5aea0b233c0feb88bb4f64f5d86acda4293b7dafe0c68b4b8f73c5dcaa9170d0d9c741b7b5e3ef6bd7c2b8c20ecc6f834348103235a7d6579a8dd8f329b10072366695de12a4cb4f0baa1ec220ff65b8077fc3b59ad13b5f78ca23c391d3e85e7c17a4b22bdf119dbc11b57849d95aaa2f0d4a8bca36d6afa7a0ce17a902f9c49ee3b67fe260a4d034010ad524c5f6bbfa7072226ea005c2c1ae2d6273f2c7d0e532b9078bad69bc4811e60c1e142429c6c0c60a6838131666e06f6c7ff2ea85d9198c05b4f463937d4b7e2e99e56004a8fa18282a91764162d43676e154e62b333a04e132792327e4cfcc35e873d37eb261216d7c2375eb22503c2ba2efd0234714c43c76ae0cb997674330e51071d315b8466d6d942fb7f50402505ec09a7ec503a54bef858c42660efb80cdc38ffd7ba404bb03f25a5c2c8aff199d520e80029eb8595a433790f9745cc08079426ae8aa56093cafcd079ab2a967721d5ff552fee141a53747128cc287d17605ef4b3b2abf5975f2eeb3498be4c0f14b4d73ea4a33809835c16aefc263ace7c55d8d8046b8ddab82e0ff1070eda4e4322369218d4aeaed3bc37d7752dd248603de19a5c4c46d6e216892aaa781004f0d0e0796c27cdc0eaf29ab95291147b133665048192b4bcb4fc8a321a2c16b3cecd8e319484ef6beca2dbbdcc49027f6a7bdb109e899606fc8e7421f13dfc5d65ab84980b52a4b2f4842cf96d4a086f9e53917376eec56fd1e94a3b7a9ca04fb9b9e8a832646b78564b2b12efa6afb8d42fa0520b615df8d34f64842b527c89a54e536d1198e06bf8e8fe770c8af4f65dd979adb55bb6192bcbdf5cafae04f43c9aa8c6b748a0fa82aeb8aa75609c738c52c71f84c6aae21cfb27277c242f1e072cab737946dca73f8487df62670552207a07b88245af4c4a222289ae9b94e68494c019fba9c863ff8aceb3c1a23982461ec3ffbb861564e5239443b7f2fea7632b87e5c745abb9ea578836464335fb18353a068206cbb47a8838cea6ec6e1790f0385497e72d756b83d3afa5ec7c821adac841961a27d87aed7298ad513f22624f8a79265506dfe8031408e15370536003ea2d13ee1babb4747e9a86ec388a4c0973ec4ab78e5fe7a617c9708623ea9417ab38253b3eff4a64949169ff1d5d2180f8f4190ecf877cce19c1c13dc170de22e9cb85fa6901dbab2f1a67e7e17e9cfdabac3af6c8b678190e39ae275b899944296f6a5bdebf11c78ece821010a77e607256512019389ae5d74699360a95aa219c674797a928302e1904af301796df74602501c1b9c16588ae46838ecdd524de2d3f3eaaa3d3fcca8527ce09e4d2ef9dbad92c48a0a351d5d389972e592b2e731c9d1ba745703f0ff5700ac3d2e49c882308469decc882960f71c063b0189ce35dcae342f713dbbcac39be4fffdcd63e1a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7750c1cdbdfc95831f33f4ba49ab81c998db10597ce329f6d08d5283b86cf685befb6cec46ae560904013d24d3d705bb150609840c1940845bf392fd6c3a9af3ca0ce7e6b8d4c1dab293148ef26b9501640ff48892d8064c49f49775415e3962d5fb50b6bb3a7f3382336d7bff29f796d839f584cda9247690d9e62373ac583684e16146660423a0ed74054c8c481345f1af5a1db2dcc3f3c53aa22fdaa32041dcd84fbc7d46aacadcad9da7d81e3207982cd7ef63ba99eadbc88f3a5742781ea5a199a9c058c4c7687068fb1003aa2a4f7f2a495f430b22624d1b8b3ca805453694c928d53b806bfa2b3b7730d73e2c34d065be6225e67206c4cbd38346367a1f4f0d6402b5cc7a0452e3bf8489d52defa1f33cf31aac906f43c4c03b1eac60420b54621975ba5cc2b1d48ac3064ae587ad07633d58b0bff4ebc686813c61e51d4a972e576db9b5240359a723760a2e1524218826ae7e8cdcc467a98cf1a3994157936b401fa0093cece296225f56114959cfdb4bead970dafbe20409f0aa68186da52304308df40d1885daf46f15a63a7cc157887c3a46aca4c69031341083f77ceb5d1018e79a0a56e6200ff7436afad8ba64ddfbcc89647996bfeeb4695a0e5b357a3c06b5d70b8cc0610b361f0d80e755bf590cdb0ad1439c4980db892ac94ce81e05d68985efcf7ece48797d530726e55b1cc0324ab6794a956c2d67e7490e71bcfab7599e9aabfe0d3405d676348b7124e3c000898ffbfb9ebc7c19bbcc168a361aec90dac4929bda47d25a938b9d4578837c50a1d06c410da39ec644ecb7eeb396fe7ed90a0318b10e22cb3de49c46e0789f66703da3fd96f4723617a543820d0531912397b200924ae709b05e7987eef9ec38e1dc653a791d4d383420ea313399d800e24396f7e5147710e98e9f0408b47c2d94e4dc0f71c89b11aacf1e0e63853caf571b6a011d2b844f67e6849177a139287fab7803e8f70e49648eee865436a7a075c05c25bdec572624b27361d12bed79f3cea7011064a2b539706a490dd9761886345a0b6da0e2bec09f8d8445305075e0106376979c16786223f32bd634a335b518c0270ea4fb8fd41aef889bfb5227f27a74ca4afe659c9a8fa7239695839f6dd92bdaaa3a2c09e5da0a35b384f274e20b1bf864966dd6c108ee54e08c49a60604bf61679b2087b0fc7f3e96a87b6303cd67082a740b20c62575545769eff88139491d5200d65afd3286c731dfbfe23a260ac20cdb3041140187eb25ff43ecbba6ca96a964b5b8ec1fda7d9ea046c68965fd26de2826753617e83c940c392cf7f4ae9c3645f0723dbd8089c3ff430e0a9a4f7318feda676391fb6884aac6bcf0ec646535e638fbce061c14a8d926c54d8a18cd87b77b905d2d22a75b5e7b7e648ac6a3c1bd5e9e40c5f5e1761013483974f3cb93bc505ec8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha4871bec3053bd4df763a4314c01dd7e5de0f84d6c3ce257cff2f9f9a98df6fb4ce40e6e089b78a35e63e10eb85830b13c0f843d5558acf73ed0deedb68d1519526edb54f75eff59cdbcfb9bb8fdf05ebb2346c1df138a45b710765678b4d104f81ff8fb56c703b98033609dd5124963c3eb285857a155993dd28a65c70b5e64210b4bc6382e2c43bfb9b141348c0aca3161c09f1416b8fa681f787a143036d33d6a0320239f30dcad6786fd50e26e0212dd16e04a2c9944a71f1ae71bfd295ff53207cd96ea245875935cede9425f7e6d29f2fbd5e4de85e44c4d953d067d95b091effb5e0fe08ab93f10b005372ba24ad53f2af70a58506d2f4ee54349d913a95315ab79bd959a5d9dde95b781c7569f3625aae4ccfbfec2695bca748840ec1b51e50ce4c809fd20f6d4a4eba4ed5ae4960c7c40f5ceb479e7caafd653c015e09e70b09781271000f15f2dae7d277563dd9f822c769114e03d280fad3c9005476aefc30c02792546dc73f24b8f705e69a0233f46be9ebbc5e4254f4572e36731f249df5b8d63dfc6ab0a3b1165f3b6c47d3654a4cd724481b0f771e9424fa4cc37ac4b0f074bcc2a5a0d62f11eb25b9a1c83ec58ff2b81ee2f4808f7004f2ba9127bd0abcf5ceeb98820fa58c12c8cd7c7b1cbf00f19549b24117ed0bab0c6b693563db1c7f1ceadfe384bc59504b77c33de3d7d23c04fe6c930ee5648fa41701052eefaefb971626c7722a2907906e3531a2f24c61517ac10d7c2898dba570cfbae4909d8da7fd1a63861bab5d7ae13dbf4293a929bf3a588bcc6bbd84a581f8c66f64f9a68342f11d5fdc551700c4d18a7f3e4942c54734951076e445735ef63f0da38a5f2767c42bffb85fdcf1680a2219d4c1a57ba644bb90d30931cb67b4d54ba23cb70d5a0466ca597b04ecc23e98158f793d9f68991a536cc6d6e1644525c79e9ee533af58b959b301d01d1e86f7759de8f485b6a341000c8b1b24c924445aac8a34b3c4c7c4827aed3077f60dbbb460247b531fffea1dc69ae06b1271c7d554efea08ca9fabae6ab18074c06cf99d19c18a432193f2daf08e34478c0616b2ce22f283e78a49a3913c32b59f90fa6d7fbdc8d8e36149da3613099a7ab0a499c613662e5db2cd1227b42edd26333d73b6451ba0eea6b6f94c31b2dd1dcbff663004735f78a3b88a612625e147bd2f92225b3a9b5ce97834c21e971ecff59f1b56a8746bf9f13f7da010e9d90e4d4ce531ca9ea39806cad68e968ba6a59ac44c74d1e59f8b8664a110b0a48a32eacbe3271bbb065a07b767ceeeeb62c15bc9e6e30336ff389fd5379aa05b684566b6757b16aaa7b345e8e22a7e2c87a404582dc23006126c55331e8869d77b372a4a09b55824f56d4202f80c990d27d7260405e043f8a9e92e972a75467319fb4369697d00e1d93c3f1a3367b558602;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h2162ddedae95ae9c3d9210032b5368a1ec0a50458a3aa61637b3dd19e70ef9847a8631833f354795a8e747f282a550f20929ef28453e8de13c1a2e0affd7a946c7a61c7579fa709b917630279ede3aa597d8a6a10dda76839cc1f22f1f6d5baf00f496edf4326dbba860777ca2b9ee069b109fba51f7d91875a9b13743dafc932a2851ff45e59ec5fbb980a0d277708271269721c457ec8ec4a9976e911913059eb0c7c22ae0063fbc0b8d8ce5d339cacc897563d5c2d0bf5f91940f98e84ab8f4839673e342585ff9b18a4eeb97a3387c9e31ca24a3954c579f0f024bd17d1fbd932eb7456bae3bc2f12ff50cac06b8d5ebdacc93d3a096304e22fce8ef4d0bb832fb0d544ef3e6d61f85fb07307d048d90def78614996fdf43830e66d02d22f8098d980bc65904cf00e6ca6bff44a5f8ecc937980421aca7d73e824de5097f1b43820905e15aa8dc43ba47a36975b9000a189f02ad300ab616c44067a251832270c2ceeed84e846957fab62ab6facf7867fa470bdfa5064b780f2c424e989b06ce4b053f0fe1d169d62e0aab92b3e3d922f335485c5bdc38c0c97684b83a958a08ef00524402bbebfafec8f557586d68b6db3b704e4eb3d4719abf3341c59f64cfd92d190cc8a76cd14d88300a7258593c83a6152151c70f3036216a1d55aa81e2c3670df4ff38f02c6d34d84493da85590ca60b1c7c483f74ca3cb0ba84c155c1928f4c04d8d11711a7d9d887ce26da6e7e98213ffa4a34acd633bacc002624de7225c727a18422331962e74d2f29abaa749278ff15f1de44d0d8eb5e113e92bec8ec23ec0efcfb2c21ea459a890d2db0e5d69f0815afa98bd4cd19949306c7ad549bbf05f855392516b50c43d672d58ae29f0eb428eef71af25e320d0ee3e6b14d28b55dc942334ab22923ec307a6c6c4b28a59b0df20078760da1fc378e1fb40b87323064a7772880f8ad4da9f1eb6c6294bf02406d87e2e8e8db7b738a5f013e86a5fb8391a974ed296e6d2fee8631747c9bd113ec6ec0c19124e73249d553862d9fb27fa06221659c1c58fb8c6d11945e2b816ef00ea79538741d2c51e011cad2733993fc3dacf626e4a5c3948dc89591f9464ff11050bcb6ea67f64dc43be5a5b495e71bba529b6cdac424f444620e83b9f249f4fae6f497f396b02de31e5197aac4e64788e10b0f3b71391e6d9e0886f3b5eb8817336fa9a87dc58333705001ceebf3599e84234275f43ff2352e9b9e42be57c999d3c985e9885c50d788aea5684ac6b4440c5cda236cf9caa921c3acc127b7fbe6d2a75cadeb186236e42680e7bd646be105c5fc98c772342f80a5edd4cc46798479e62c593548f98b16cbefd2f0d86133110fd6790742ca723095c199447974482c19e7c60f8b0c3917dcc08a1ab87192f446fe152942eb8dd74838567e467bcb4ab641c69bb136;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h83a1d8515ea0261e4174b2a02092aea47a00c3d49f94fff96efa7cbacbcdb6d4cf772c6228ec0f3584a074514a0c35abab4e9f5ae66023d4f75ca77962989b1220b333ab2681314b0a454c84624ffedd31fed05e033ea3ab2caa83975e20ddd654edc7dacfea03b685b38407f7426e5c6d99b1e1f15d206956fde4e50b5963b1e5caf3b563836382a8411602c35e7b2653322b05b84108794861d6cafc66a91b4d1191bcf9119ee8a901435fc830418fb2baf346233124c5f0b25fdd301a22b5fbbb736402f46b4d78d6650bda79115f437a9a6cc265eac1b318a1c6d8660ab47fb9797ea6ebf614939739108e070466478164b846f715290b86ba25ab0aa0ecbe2c8fe3e1406ecc3e69550f7cfd56fd613e2afceb23d1f49fadc480f310869a87eb050abf501a5c4719a5591965f6b2166d0bf585bf8ed1b51863a2f844a31d0cd54d4cbde03e49553f1dde5a215900c5ff4bd1b12a257cad63e730104196dc7ed826b0624e04b4d6b15b5e8efdf83bab4252be7ca84db7b80f141cbf1b4d47d91a4e61c0453bf1d426977b5ee17df5a57c1df8164a52d3f25f39001c1d4b66e850066cd9b4a3dea59f8768465f32014c829304b0488100ac614949d04f4371f09c453dcf4e1bb14edbabd6d4f24e452f1c3c96c0b96d33ea4f973754e00f03b2438e379d052c23a6130afcb1c36df4080eaa4474f86a82de1d72cd8acd38390a95e19f9774d0cff015d354fdd1c79721f9d58c7c8dcc761b04f92cba85ae1e6fc072b3c11021c9d82f920a02771a697edcd577978f523069ba1d0dd38094b6a36f23657f072c9d62af9e44c26dca6e723a40577796215ee29d5097a4b6c0876f35a134a6b01bb22d5541ecbbb1de0e30bf0241a0bc49f0cc53e8fc8805bc245e5a33ed93792475fdc9f8ede7809f9a6bd475dfa234bff0fb5f8335c3c10772784faabe396d0435730a3ded531419b955fb926928573bc08a3a4adbf74925588ab4cfcb906f6872739257696cb5f1f3671ed20063964e64b29270f925b1396f59cae776777657fcd4443942b8a269ca50b6db031b1a890a0d34e89d0b1a48018b3803b3918430d3a401870fa94b93c3fdaa8cb3f90950617088510c74d78291200907fecb65bf737864397cecc73d1d683c0d48a811da9e4b8dd40cb550a8e900d63b52d0eea0e5dedb486c7bca58c1d9d4cffbd02c2fb1a92b52ae2fe810bfa340798cf89a95e2ee523e1eb49c1f7fb8ef629e7f9353f4ea6ad51e1a4f6e9b5e227c1e6c3098be140a7973682ee3e2dbd298538e20c15bec97ad633a858d87fad160f6debeae4f195390c7829e949fde55712d04ad9a8465182a2151083be0d0acbe71c5a17caa399db26212d1d4fdb8bcf93dfc4ce9f89f758ae539f2c3b5bd1cad245a0243fecb4a2904a34cf739581dda8e14f2b25d0bfb287b3a2c8823;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd42e32163c27af1b817e940ad4f0deb53dc36ce2cff17b55fe44478041fb41cff18fdce2aebad201854a914ba4c914a5dfa8ae921d8ed7312514ae1fcf97f219f6e49062cc77120687731a7323a1f984250f837ce7fccc93e5cfa8da9d0a89c8cb800a59760f8f546f5282f1110e488eb9915e9823d56d79c75c72bf5048e4206f23d07d96105d92fd8da5afcd6d09c914d2aae8d608aaee4bbbb13895d57af3bf7ed02019389ce28f6d7e90bcc659d3f7a5442bed76dc38bde56f6d136dc602005e4c2f524296a51e9109c0cdc002135c53b4a46845dea3458beec319f8780dba6fd302e11ed88dc2811bd32826ee7882c6924d518fd1368fb6a285df46315b62e8f84d2d78a82e96772623d477edf99ab5df7f6d735336fbec7d91dc2617fc395064f1104e4ac6640e81283174d1a8c1ee889cd27eef0156842c67d881ef3fd268116983d7f9bddcb028059fb7657c1d71c32b6abc44203549ff51bac359833f3cb929b41cf1132d7061340663b1dbdd54d33813a4a95883c7535526bf8261e63a127bad202450e0c5df659c143890324c0d8a2f018ff165ef4d27119b4ea57d0811a33da3efa9b1331e1ee96b6d5cae274392c5e02853335d2dbc19024c542ba29350af6dd9a5ab9c076bf9ddfed1d59475942db5319cccbf546f0e01ea496b8f8820b82030b4940dd7466e706afca3113d40df71e836a2a02f118ee33b27eaa64d721de7eebd8ef1792b6ea38824b1ad90bef450128545a5b372476659bf81d92d02673e6a8e617dafb08a320aa610ee87d0ece4a6f544e6779268d6be91f7af1e8d93ef63ceeb853010b948263952ad007d0f48cf2ad24366840c88c7ad3b8be3e170377e10d64a874ab3bc7811b5d5b5ce198e1724fcc6f56ee7cb0a199be36b93e35590458530ec67211aa47acbdfd2a02fe7d9f9f1a819035a0cb361fdf873ebf9a781ebfc132ef925ebce59edba762a4b39746042c0f3e434cba9f8338dfdc00dca36c9ce229979da5a9a93ed60a2464ebd95f7b0ed567202c34c3bf976429b24773edf8f2b4793bd2ac102fccce92d60f8e4f6f2b7d25e6e5b122ac8c6ed167c4491df1f070deb1c7ac124df75f093540e2e6a7b104ed6a881417ba1a363bae5148b70fd7bbde36bb32949937bc18d2eebfca8c14276ebb42fdb13b635675b71c5c239f4d64b23b751ecd031329125c60424df9b3469b8546f818f7397ea6bad5c273fb93931122fbe0e690119cb48a372df00ace112e6c4cde8ce0e42614bf0f09ddc54272a6c3564184d6c133e7e741e9f2a69775c900aa66d8afb3eb256882cceafcff6d8eda7dc02b84d99805207fb457389be122241ff817f2f03162e495c74cfc96b9645f1b5c768dd21e476b9f86d5dda977ad4bd564e2a6dd86df28a755785ca2fdb31b0745d076001792866554d2f3933d3a96a3823f4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1a2a21a15c42ec1a99a7912933096c375e9901d8a7dca998c5ecf88e2f338cb4165aca977aa8dc61beea9518f60f51ff7e086b7901505a7e527b55eb797b65d9583a2f127cef68555087ba3da46a1f4e3c36b6f19ab5ac06e1d2692cc6e448da972ff443d8c5b8d0cd8d9431ad11a0bd0c1c83c1dadfffa4ac070968a292b5c2fe7af0bc1ed1adf756ed31215781aa28583e0f6d4766f08d16c8578d410e32055e83156d29737ff50b4fea0e5fa8a1849a6c06591cdd89104719dac0cb1a7f494ec071e74182717380256aa6c5444f25cc777712eb6ee33e5f48ea53166582ba032d9fea872154d10766ee85fe306246e9fe1588e22892e423240c280e6475dd41204b6936165e7233fe3c94193181022ffabd59ce637517cc42f3bad764f3319baad7edadf623a9be89b6fc686f1fb29b478dc31e3895e539b8bd2f02e3358c63629a5c19bd812b6aae1ce786e0526cf78ae33bc47446b191fbe0cd3b14998235b7952bf8f44365164310a6ca2da56eed018d27e5751f7eadcdb0073623d3287d7fdd3c5477216d70827e88beed779222062e39092a8e89fa8553801b7fb21a867e2e4815a66d18150f910111948d84ed3784ee6f50c80f9c578e65efc4bbbe65af38ee328e37d00887ee73127e79db4cb0afe8ec8a45d94157f785d0f7d696b2d2a0c740e54d61d2371626f14ba59662d9f01447933d9bcc503be941d0c6f447626a12ef40ad5544675ab314a3049d54999c0d08d6f6469a320cb27ed60950dce3a8573f6439ead69d40e676aa0edbdb1d1ab7790bdd5c5f19f078a1c1239c4c1919e81f86a61f4013d46a526a70f318636f0be61ba0a308e4faee17246cac2d608cfec337ce1bc3d5f9284d0946a06bf0fafc3e8eab662db7657565bfd575321748d4d295390eb4abb774a0f028d9d38ed7be8957456a4671fda0e9076bdf03ed4225a46f65aec404c71ebb5b8d7a01fae08818f1f71fa1f3ef9e5ce37881a2f2988f2e9721c13a93505b28e0f06e02e303c8a4788a19b264b78cc5af0bd15feff12e9bb4bed53b08c73fb0e604369cb61faf59233df0fd07a7055474d84ee780bed704610cad39fcbcc44be26aa4747a7569e90bb648f5eeee667ffd57d12a5351b4937b45d34ef833f61a44036de574c68cec0ea61c44511f39074d83ebf57ae5b8c35b959cdf6b73bbe8d21baacd876680f9b96f40272ba5c005080d94fe69e819f67f56659b21bb5d86ff937cffe732538b0d5b1e962e1d78221102fc6f9d2a38722a3820141c472538c2d2a7356cf99b8e1a31dc393a72da94396a86d141116a34e6ff24716a1db83ef159786f8312d171513d7156840acbb73eba88cd5fd0c90735912ae0b532e66a01d18f92b26f4d80bec5abe7ccc2fe53d22ddf2f46da9b5dfe1d88805b8c076ce7cecbb5eb1e6dee333f935409caa98d2a21e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h386219a2ab6e3c6f1a09766e79c4113498af42e13006375ae60420acaacaac7e555756340f08abc8e62adabe953c1f8e8ba9a780cf306c6244e0f08aac17583b2709641484828af724786f1e594211cff0f7ec1c72686fe7cb3bfb995a3a0cf2e9da1e855ddfe750d4aef243c2a1835de2e66bcfef2671dddaa092c0d13ef6e85d25b64bb1c83e19a5c0ccc26dad925f22fce2233146febc3dc57078dd177829d7f7662df40dfd7f97d4d40a3c3266ccc15303160daa6eb7392b4de5e8d5a994107ffdf2c0f3930b0be9281a814538e60360595fbef022a30bc4fcbd585ddd4d5d32eb80596840689390516c4880b91454a9bdb5f6dcbf9d2ff90b283f76131e3efeca0882ab23ae388cd4cb048dfb3b75050e2290dfa9a27f534a43788bef81677745f765ccb1c313897d96a562fb354f9b72ad8f58e1c626afc942f1d09ff7d5085c2a41d714bf7f1793d7df808c1aad382d110b55ac705c8b18760debcd8251ed5204b62b4001bfeb8d8545ef66936c923b92a40eccb385a7576ce9771a4d33bfbbb32a6cec72d39c77e5b776ec1deea58d6065ac46622367ef66a790b4d68fb3d3d2772b3b3f9e95a3532fde2771f07780087d717ee3f60533f69ea29e0f886b762c3d5a3b8645121390029fd1343fbee75d218b9d9e1a8fda71ed31656d6eb4f12e11e2926e28231659c052025b9dc6e24821b1b73d7115db6fe2f147d572ca6ac39e8ce371ada008ee6949a29882a31ae0c5ff3ef4d14fe98feecc28ff8a4bb25e100889fd3d46749bcdca8d020025ae1ab24d08bfdfba6e5ef56f09e3820657a6586fd9237bc4ddfc57cc5d5d3e46e0361c41fb71156be5437426a11936a3a30468d42594861ec13f76a53dc27d8916b2d8a50bc890c3e1911f85b0366e1965aaeb154a5a44772e22ad6839cf4c96fbee95122947aa93b8d73cc9fe5c6d3ba82969b7aa5a340908736f44498a8f2ab796b3ad37e2db8a44b00a35407dc419d8c7e20ec6e5f06a31310b9fc8c3113cbf171e18f3734d7044b14c4bac2a02bb952e4f5f6f921bed632607cc34f890b4350f97ef744dc35a62e9e5f5caa1f419c8a3f0c7aa13325def03428954f5ae2502cf18275f6cede70842474e23cd99a2aeb44e05922aaa220cda22ec8787cd4f7c7c5e8c1c1750bf68b3320034fae7694ee99b0dae118ff4334a11d7c741c334dbaddbc59290d1b17d7b127b6ec9cd9d628086e05cb65d88e775bffb1f68ba9c2fe918f5b8d14b9d0e0cafa7d7b591b1e9d649a8a2d050c5083ef89fe10a88bac20d435b3e7810442126d84aa652e91915d7139b34aecef2b09904a99e1cb0b1d06459be645fae06cbbafbe80fd0a9283af4180a4e0c4b435a2062cb36e3554cc1841d4af8db3b9ddc274423a84c48565fb0e2e8d314bb6f82aae1873c8ed6f470dfd474a2ea7aa5bc7f9a14432d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h93ae5eaddafeb573d3ccec3aab252b2ec5c7ed9cd0c89e370eaf4c14a44ac6adaf4da716a1d29885f5e905c3a9c579a16d4afa2b478bc4952148fd6edb747f2f75366c45dc18e32f995fb75b70f4007a087833cb4258f20400c3963513dd13a0ea2694a63f19ebf8b40657b69bcf70bbf5fbab2fbe572871e3a1d5744a8e0b1a38a0acc6a6da31c17815723cd780f7c98c49fb517dab4017f3029aa511aa9fb773723f9ba17688e26d2b56f087de85032803ee4cc31bae271a99162fac8b46491036e2a97929e41dea01622a185b348e375bd40733b15f5b9b73081a3a2ddcd23c1459d5748e84e65f27304dc37d8e9bc906e17b46f51752e884fe317de571a6c3875979e62ed6aeea89be38a70a4f44a8db5947c382efb7f6a5498f7ee5991b1371290e1883fecc83cba86a7366ad607328f151fc9cf45e32096ce1d487dd9f725aedcc150626c8d8ab3237219c7d52df088c6ee44715a67b3400fea423d47f56ad18aa46b5f3b25a39cecc1158f46f79d1fafe4e7431d19307c5ada3942770068c9858357b93bc0a94f3c2bc527616a2c1d31b78cd2746599847520abf3c47d6e310d625f634d4d36bdad6e662c7cc047188b6fc1d1c3f0a594b693016cd1e8682f2329da34d7280faf2b862e6ceeb45d316ae4e3b30f8082e8f357534e470d8c2e6b9cb1aeea70adc5800809ffc279f2e73b7cffff8973f5ebac555227cccfa899b419ed582f377dac05e06708643996629f1db6fa875e8ccbb6f9632e52a4a12c8247f54cb50ba7b874a8ba0691cab2c242b0b522dc2d7e5df9b235f30524fa14756919c2faecb4fe3bf32348ad2b3abbec103ed2c0e466fbdc523d04936392a73f39797043fee7075c6efbdfb8ba665bf0be997445ac7e8176da4d91867d622109c939240e071e1e70b5263bd206e0597262c59ae07c798630c9f7e2473ca145e9f91be7bc6a4283320e3efd77edc53dd88c0ec34c4872f144cbc644968bcf3a7543d1a531c6ac21b600b270444fb7caa5d89ea2f71f689f992025c232152d1c0614d34fdb801a87a654e11ab01f09101e7c463606eba2c61009a971946ed95a70dc8661021f9e2b8c33503ef651aa437f1d35b9fd6fe20257b26fe4b7dce79ff67279f755d400c697a81627c14b518d0aa7bbf1f8eb896b28ecd7eea28a72082e4ca758a133fc57a06897a961e4b66acca7e003b9a60b67949eb001b45de650bfd904dd5d729665af3585a25e1c059646eb63741f05360b7ca13e211ed9a09b0abb9a97c50220a6d7baaf478ad69a3235f9bc93e6195525661d9d6c4f016634ebe6c34f8bbb55b9a30bc8ac1506653738c527bab77ec5ac80e0bc978491a0c699c56b0c877b1336b62c4d0ebd452e26b8436b28e1d8915397af4e58f4c126643018aaa8d03ea99759ceb3b53e452aebe3241fee7271373abf27d2f476c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h11b56096e0bd501722ded9437a42fd4ae3e2a6c8f2671ca06f1bbc6d7e8ed69498b119e8252c00560070a31590bcb68e3ad9c7a3ff13e9a04fab32579bd7490e3c48440fb7b00f7e984d9b7658842dc1fef8c84ef7c211aa112e99f624549667750d6e154cacfcb8be85ead29c089e5991060c979acb92e63cce11827cfdc14a401cb4e01fd9fafd5d819aed272c569424dfcdff7c43929840ab40a2d112f2305f0a2d08a5352e291e86d0d0141c83777c58886a8d0be852b6db6d8c78f0faba98870aef138c846a57f252c47dbd6ed685441311a04409b8d338622155e44112c7c9b68c0be090b5c760abe4d8f1b74be656523199128735b774fd6d2781ead4f6cb6355b70119cecc944486772a1cbf2b3bbaa79def474bbc1f0e678179e7804e594278350ec6f6dbc98215d563f7678f092d793ab60283b7065d793b2f63af66f8c7d08185d6e562bb11af97ee8e003275fe8785664ed8fe9aa20f7eaac2b31cba191f544a92aa0bbf2eecd4005b814337e69d9ebe96712a05e69c8458767b317ee4c5c475faf69ae8c50769ff2699e5b68f89800e339a7f164eeb2578ae45908670b37b54eafb11a8b4987099a7c329cb330b2712fd0c41399cb3b396f5681877ce6baaec3f9d0079ca325d2a53bbc64bef1ca1e1bcb8fbaa169f530903cd87c081e2dbb0478d4eb45835c0df0c1e66c8ec04ee751fe6abdcaa8e4a687aa0eb604f6e14bfa3cc9ac2ea17409f654055f19925954b824f34eb21fbeac90319e3d35de1002d86becf5f4ac3ad56bf2965bcb4b47bdacb74ebda505e7be2495d31e4d9eceba81bdbcc0979f07f872c3477e3f79b613ec72828708eaa717c6395befc22a43942bb3d893f13e5d10b8d4cbe7d437d2253e0dc332995b33af673921b664144858be0eac3522325f3b9565f1e2f45bc1d23128c28a936c34a8f556043a8796ed3913bee3756925e145fef761f7b364c0651e8c25d4e7859c6c1bec3ef764bc329a77975d9d3ee6b2aab4ecc459d2d38206c782cd38e5703bdf952771896cd785918635da912b65b82107544d5b7ce1200eacc555502c0226c213bec1d17e05e4a9e0df857617168c3a4c121f83cc95383fa9f09f0452832577bcbec96eb5293f45f64945e82931ac1bc85bd2f35712cea13ae2560841fc44ae28331664e1c851eb69dfca0fd09561cb3148664bc274da188cb56459d90c6aed3e904ace5750ea6f912b1415a17d752f6f5da0c45ea0f18f894cc2fd9a36d977657931370974b48044065016bc936396461115a21b5860ee5f39e8d83f859ba097345a152b28b4ac390ee8c4dd91cdd5b38029a2d24dfc60ecbb86f285c199e2a5cf0ebe6a79c4a666d486cabea322ba86fb15bc4f93b54b98ad604fb5c5bf276ddb9483489839f865bd257a82ac43806b52ccb44645c3eda9499f681813b5e22a738;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h903bff38961ceac821a6c24173c91f84077451e94fbbe4ee9a4ce32f4bb4088fc727b9af882b5304ab61999dcf5e33c7dd5cb3226b46054c78059e8b96b9d6de32891a36b01fd28f9b29d5c57753482683c5ef7df6eead94b484918d8f2803334eb6cb876fe3a033ec05f1f714dc686297ad0c922b14a2557d4a2353ed116c0c1cb884d197ca2b997eee1c89ac4559bee2601fde4f07be09b141b032c59e0ce687a909d9a26479979759bca231af7ddac80b229ba6b975f812afb684e1def52c734933680d8afb40da802db8f25647454476bfa28155eb17ce352d4e1772f0951095779e8e335e6b7a085e825e004410ed349721963c2b264f7801bb91e0dc74c90d7538595a920afbe9f54ab8907f98fe6f80f78ec7912d0e30bb40ddd35ad1d23e50f2796c7633520bffa5c6e9d0c92ac9f5fbe467c1581a1322012639926fe5815e2abd4eeca6c67a11a6e53b1b9a9118bafcd64efb2c797e943ae2b6e64c916f2be786106403eec941f7a43072416d5d593a3289af6a38e16ff9cb8601196644438b8034b2a4dff443a61acbaf5d6ce912d4d771c070e4dbf7b172dc7982ef85998b96a98e27c2a06f91818fab7f4a21ebd2ff74526c94a76a35922ab17b2c2f8974bead44104b118f1435cd54eff31204f0cc1b80a37643fbe04b4c6430853d85c5b02416528eda78ad725c415a4fc536fed28334b7865277fefdc24597155f615e4af9c69d3824097034474cc7828f9ee9ca307f801573d1f778b2989c7a7da3f5974c7e69c484ec22d88d8527467157bc0a13e55dafa7cac320aa9949bcad1fe22e70d17aae1f70da6f3330e8e4dbba58b6c2538717c50ab2b7002c7fd3102b2e0d71f12cecce77e36e3b5ce86ab96c2397906eb9c64514d12ee3deabc71200de81fb50c828412aa7ae6aaf34406a6701ba3f99257f9ef51cda571367e48c2b37e8d1822290b7ae59d19406be36ea08d9c4ca9a0d21cb41af614d189852a85e6ccc2ceda867abb714b1c4b039b95e9b5fd02d5a30066f0ee7efc79b93dbe2bc8e8800bc3083fd2c981b66ec740a92156a7e4fab16d7e3ba586903108118fd594ca10efca34d6533ff841bf8c4b22e41b831954378bd947ca1a074b475943ee23d2ec60b43c5c1de1129c75710fc3aaf45278fc017aea97e44822608b43008bddf5a4ab2d645bc4bf63c9db4a2c37c8f0f8ab50068d8446d9cf97f75db2b4fd50c5f3f31e299eadd6d1dd3760813495c039356963085efb126987f2af85e35476a9286fe538b9772e6c43137a6a94f1c2335de165beedbe0c029e43e895f07a802dc5c584b02a9eda506f745e0d54c9a0b2ed4a92eca308fd1637bcadb3e573093d2678f5ac1b3f4227cccb413aec31e789c1b81cb7a57c1568759b830851662f7e26e47515abe8ccbda45dd25593f6d639b4270bc34572510c581a652;
        #1
        $finish();
    end
endmodule
