module testbench();
    reg [18:0] src0;
    reg [18:0] src1;
    reg [18:0] src2;
    reg [18:0] src3;
    reg [18:0] src4;
    reg [18:0] src5;
    reg [18:0] src6;
    reg [18:0] src7;
    reg [18:0] src8;
    reg [18:0] src9;
    reg [18:0] src10;
    reg [18:0] src11;
    reg [18:0] src12;
    reg [18:0] src13;
    reg [18:0] src14;
    reg [18:0] src15;
    reg [18:0] src16;
    reg [18:0] src17;
    reg [18:0] src18;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [23:0] srcsum;
    wire [23:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1154ed6d021cb3c89d37f16071e66b415fd65087d287a1452ee0401ae661ba0828176ad5f014ef327e016f3a7b1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h35ced8e1ea20b0fc59be0859534f22220dbe8aa7e551f883903a37b2bd4d2103577e8c45929a5aebfb78fab16d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1afd08a0b6c98ca31e0638bad4086863d21e7425aec210f82f1c948e01dd793cf535ea5b0a435b45c0d38f086cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha4746a0b55868cf598bf5e643caeb0140e92c0e183a54e2f76b70b710d7640cb8326d73293a8ce205cd2dfa00a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h67ecd53b01193836721fe561d13e6be174fb104dbb323299ccb832ec0f4141ec31ee81eb1d39f9c35a3d74c50f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3dd1148dd80d949c03133fc6845cd0125d3e066ecd29b2d883d55e50ccabf9f4797e8f10ff6b8ca76c1a5c0b39;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h143215650265e4165cdce986b48c7289a3af85126a1bef0086d58b984ae3c55c39d2c1f50525eb5bc4796b2ed47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f7164bbf92b7b26471be022d488051d93bc24dff84f0369ec338b116f114bd117ead32dabd26603a55e4810a06;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1088d2961456f35ee407e6dcaae38cc6142e5a570df2e2ec9acdc95c3cbf36e63d588596446efaaab3bb309005e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h176a15893f31fc2d13a4d37fd0cde37df2dacd5402c9b2aef318135ad42a50e19847e5f713b4581ffbf0e75e47e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11702892fff41d1b8de01b6e8a8557a75a16d65f8f4de76ca505b0e396da291ef6569d196f2d05bda7f084311e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ffc7d37ce7d466acd9498820cba0f321d735dfb5730fe734ae2c36658187ebb979e0fdda34a7a93950cbb66dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e226bd0ff15145a9dc25ce978007aae0c46805ed09488e9485f65dad2f08d1e00ad058b62d9771e7a502506347;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d4832875a46b2c6d1c8ffbbf36bb7bc764c86da7bda0ce5e244e6d7d93d35f50855133a643532f376984c59e72;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf19013a76d072aff7f56a8b500bd29b0e4cd59d9629ff5eea6daf081b7de0d049bf858e2553af0255f050eacd0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h359ec4b3c22f85fad0943a3c3bc93d2020a621d85c716b4ca7391897eee72d5f2e40f7b819496eae6234f8e5fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h81a2b83036f3da7f4569dad190a9f1a9ab70665c20e6675cb12b142a182eda156787e3a8cba6d0774a223a9c8d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12732e33eddbf50b789530c84448060407f02d90b7b92d862b8c7a100bab7e454ab24863c009235ecbdf59ed9c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14ec26eaf32ad918266490807172b377acc79e2bc83474bfa77d75d57ecbc02f209273a407d5a5a2e4f0f2c48b4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfaa81516bb3d676e54e705f17e9e4ee0d0513fdbc841148fa70c0bc63ea039df8f1b508388ee758bbd56770917;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h184ac66c651a8d4c01b319a8528a6f4234dde0a40094e38bc190fc93b4bc2790645aec9bd59be5988d27c97335a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbc1af1c99d753705f8b154571cdd9d3c32ed9929d014082dbdc5e8c52f456ef964cbf03d32c565bf1938431f19;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf584b0d4deb25fc6492f38a459b0c2e967f560aea7d9892b557e7df61d13e391c7b0db5bf67f077d3ad79ff955;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3ef490452b3b678f17122d0defd12c658d0badd1ebcc29c826435624bc175a467c0569a1d78a85412105863778;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h37188adc5bb77cdb506b2d0a2aadc65e7099c69387b49a385ed51559b70230c6e71a2b8898bfce5f3a9a0bbe48;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h36b6fada94113c85ec44bc2938e6ba0d1bf805897b594bd7fcbcfa22ce9c6ca49f8386ac773f99b77ccf9dc64e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b63578be1f9dd45fa6ded0307b9a0f6dba0c96d0eaa3d6e61fb1bef3104dc4f2dc943558edf608897dfeeda9f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1772e16395b0722c6934c065df70b8bbcf7ab59797559187611f29953fd3ec89d9eece1d62113487ff0e7c43f67;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bee70ab32892f9e49f2011641ff92e3dec0b6e32a5a980144a0bb75392faf5393fe01504c5e590b113f41881cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f15f1d1b31883f444989dda8f1e8646e7808a540de392f691e17ad1f23acc2d8341c3c97b620b006ba1e744362;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5545d70eff92ca94c77d3138abdd18aa58018d8f139d439e771c8f6f6d1b9ff4627b5ac79bf94a076db23a9c58;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf3312ee34bc216dd7feed36728198cd750ac2d873db293c1bd6feca7a0a8b84c64692a52cdb320d7528f30bec9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h677c5e0f7dee6a968c194b900fbac051cda0aada25bb599f90cc86234650b8fe8991492f6c0f2e054616350fe4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h130db7e31efea819998c1bc9a98e0963e14c63fdc9e5539b211d0703c4fdadf5324ba94ae89e63bf26538098107;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd133383355862088efb796ea6e209a678943fca4c9170b8108cf36514bb88ec42afcfaed6b45ad30e42c64a162;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h460302957b1dfba777a6f0376351bb4db0a4484e8e882e16b4b90bdf0903c18f7305b7784c14da43f6682a81b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfda106c430e07d123512cd31d7fc9ae31cf06648b2c7d3d18c8f1e57c7c21a7111e3b1d049378ba5ccf1171930;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc9df2656575e3af141445fd24240cb9027daf8e3369e2b3d1e9fb7749d652ad08b15a08ac2e69a2627df51df03;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc42e68b397805d40ca5e9de8444bc3db973da4fea4b3a449e91263a8311c748fab082a30a210a401617782dc01;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4884c4aa560259689246d4f8089ec6fbc13ef1f4ed795a43f7b1283dc65fc338d8c3ad84c96f31158677808faa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hff6f65cb62e997958a582fd2ebcfcd5a6cecd145b3adbaedfc08d0218dfe85820639449d18e5840ef9ced20143;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h143f84a8af428cc61373f2979ce06d375e45344696caf055dd436d7ef11934a71ece7bf73fa055ef56c69f40d76;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7993b1207c253090b59067887281591d104dd4a7f825affdfe6d0c962d057299d31e17cbfd13f2916974be41a0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5a781317c4ebdbb82b04438ca502b095b2047c8cb309c59552ab03eaea4bbb955cfa555a1296286ea5fa663c73;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13cc8d2b7cf5be8d77136a05eb218cd7bd78b168a28be504508ff365740b12de8aaf1ca949540db9a42c9530f9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h46d96c3f491dcb07d66fbcf99f75b21d3810124f3cc19545808f0f380e359298eaf67c56c83460306489b8e1a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h841a0a7311991fd40e99feb1745813b784876c8040c7cdae0a77935c5b2e9b1a09ba2fd6d0b2394a927f5322fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h47be1fb60fe52bdb46b4bd230bef2940d6f5490c5e78c76e3e4b36aaa6d149c19da4ded6ed01351b51cc6bec4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1934224d8c66ff433aad41a82881c3d8ca102b397a31cd47814b30029dacb747989cf250ee15ab2a68630fca1b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f63293a5ad02ac3a1f0abc236a85c3716515d1a2e63e123dbfe3b3c22b7ebd385ee84f9bb95c98dcd6def1f71d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haa1f30702d030502a00703b61c5f093498bb441026f2cd3033ff95dd0165615243325754355080200e395db37d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfacd5f396140bfe62b6ceeea044adeda0676c50af2d5fcdabf967807c5afc5b10d44d76c934a5f131d4150c9e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18b7b32c8d6ea55d28354badb88c55631c387450c50c16680ac69729a2753be4f0505cce5ea8904a6ead73e8c71;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d23ed178461ff994ba00500963e88263dfe13e5aa499436ff3bf696a6b2124fdbced3f7a5824d6731cf77bfbf6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18bb45e575366218ec8d42d5b56fa56a04d07190f2e2637f5c55d92c3752f322da69fa822555870d749cb38dd32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2c170449876536e8819bdda6096aca4ddba85f9848372188aee5cd661ca8377e6ac51bafc3d3ea543b86cbb1df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h959566e6978c034ea3609dbdb6c17533aaaf75e08b4ba059df85ceed61afdd3c55a89e441a0ef599ae3ccf2ce8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h50600aa6a4c69fcfa488609a11fb6b06204e7cdb5ba6d7d806d2819b5e04a7e810a23dd403bc08ce47d597610f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e8d684a45803e83c13be4be76b65527b73400a8c34f1b088f963d5863a5d29addcbdfcb573b34c91a6fbad6a2a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1576ed34f89e39bebc3da144f8cb906000a5619248c2e69e2bcf363997ce73d72d1927fb7e073d67a7d5ddad7cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb74d49809ac782a4c887c029ecda52df4fd83cc4455daa274f512a8a0621825520a66d4125bba68683a15e0534;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17bd36c21c538422c964541777265bc02877ee6933f6d85537c7cbff6eb6633ad6b3fb6111c9101f8830100b2d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12cbc7ef42fdbc39c2c8b3095f2783539128fff27e1fb75f235e484797ffa935b18f78d6d4bda4b0bdc5c1fbd15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he01a674c6ee29a3cb76c90d21420b15edaf045c75dc10d38139b83423f8f49721794afc2013673a58692d78a8b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10baae2a5303b7e87a69a8512fff06753dd20b5af3c16323976437aef4adfed4c75fe1ae69fed7a23f0a5c76baf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1160f52418e17888077db24749c48d5aed223fa88aa1747c69da422f25d81642ab849affa30ab747cd9603c2f61;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ba7fe10a2135dbc081782c69e874b1f996fc7c70c002e997dfa19cdb220cec7e1573073b3432e239556e9c600;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h596876a8288dc0f27223329a135c20fe714d0f6c87b9a354189f92770203df1537b4c397c8bc478d16167ef514;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb123cc1322115e47ea0f2c4495650951d6f262ae93425da66963799288438ac94bebacacce98b30e1bf32ee5fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5d7d5e9930a832cac5558b45bf22963b05abb50c150a487e9784e0ee17f050682625f019bbce4f7458684568b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd9c057c16f983c104ac00f83ceeab4edd0783b2125d9b6fc1c80659e79b4c01c10c604874ef51a5aa260942da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e1aad33b55776a5d671e5de42353d2fc6738bc847336084b630177cd6667343aab697a801bcbe208c6a991ed1e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a72421121ba8163341ac603e384c752efbc4984f7ae1319ed5a971a46fad55c9cbc74a5cf2ea23532fadc7cd47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6137532c1d16b56275d881d571f46ebef8e05530c9da7dcf675813c6557634488b639b7c56256d1eaadf7aed21;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hedff13828ab276123e01a709b91287f75d8fd490e87c52c2ebfac1c23044bb77b3ced90ac329bd5232d1e48d75;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1177c52fb7181e3ca9742636097da098e86bd19b95493596e8dbc89e2b41fa6575e5bd099890dc9cd5fb987ca4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd8701358434ac8ce1adc1c39510cc4e85d8520cdaa4605aa3ffd0665aef0668d9e300df210566993bdbdcdc759;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h823de8825b4cceb82b3d99af5390c6f19770a6291db9a93970054e83193a7f3f125131909463a519faf475935c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h805836ff8c0dbc931a469ca858bf803e8c992216331f143c8e98d4493bf1656d136f9a339884503502c7cbf75;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h132c428214201056773c8c7ad4dfac8740b9006b926bb1624b2a0200fb9dc68505edcc18c8ab567685a9958c8c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1de4ed99bb07cd73fdecd0e78df6d1d47ffdff99c83b191f6c4c9377f7edbf720aebc8794acf2f96d95d013a8af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hee1e0bf5a06b7bd7371517482e5ed51e604abf711ed4acaa5e102e0fbceb90f4f735b02c0c50a7d3475a89c5f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3c261422e925836083eb29cad8447e12b4ec07e4ef560655695b4a7117d003ccb2f6ea9a30ec178856983c78ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h69a1feaa2c52a1bca84cc6195c62415d48704cee67eeee0850ecf03ed7c71c1cfc662aaf32da57c013ed99a86c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f428396036ce92567b5b21ff4732e114f1e414f16f6c8da507de22870b55117a041a1dbd973774a6d34f8f5ae3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f33c9d4b26332b29c2e24ba05672144e558abbc698c2a678eaeb5935ffde07b813e6d098ac3afaa1be98117c8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8a117496d36a032f07a417ac1470e97058e6004971f8fd76b141d6e82005054836e63892b4cd4367e94c557372;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h264932d61b905a9ee92ddd5f3f9e018be4ddbc0a0771bf586d98be5bcf48c73e26c33e5119a1aa410e8b288273;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19df9a8bdc01a9f68d9cfedd6098bc1b4bda79af804fa278798e3bdf3ec4566be5a0803921d20342a8d9f5a8733;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd447c97e7a84067a8294477c525db42412dd22a34f44e2e23e59fb5d5d76dc7899a61a3ea888c5300c4995ec7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8e15a4e2c75c84cbc7e1a918d2711ffb63cc4839edcffd609b4e7fb168c261e6ed84595c284fe0567c4114dd64;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10957574351b86f391d27b643b26f7620acd08b5f822e1acb10a001206dcc347f244cb16f87c2ce8bd585cda1d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6e97be50040052f12c526f70bb46623a6edf061da2e674fe8d8a5682671f17944610171708d0ec60fe3b6da89d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha78464080545e2033b9e3f72a6b5d5d1259cfb9412b7edbbfc55b7225f01266cddc1c661aa45f1382d2b8fd503;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4c9c86eb3ba53dfbd0c8ff656a397abee8d86d572aa35d21af5e4a379747e8aaca34c5688c60d6146d75150166;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd62a1fbc7889fb04980c9fba6bb429dcd20464d6e3eaedec8e53ae01ad5e55c95ae1901d60f897bb33a92e7670;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h186ef9ca4cfbc37f0821bcd5309660218640233251a55d48069592561730935c19cedcf4167141146385cc9eec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf9442f8686cbb3ff1c0afb6c62579fecc9b882b7239f0d91898106ad25abccf81e09a474e753bd4635eb754302;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha087bc09637e7c3281104536057572decd66df87e91770c7d39a2bb584e3ef7b8bc420c9d049090d0485d7604b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h45ce35c637936880ac9764e862f16be96a2a1729da6189c43dc80db84ad8fe9418d2de74b49f5c9716131383d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h172269e380bbce837581efa318c1ec3e71a329125dfad8a5779f951883dad72316e3d432aa78f4d010b9a6b498e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h425c153512775e7dc73f193c327488a8de08561b6046b31f0ea2d8ba5cc67d53a9f80d8a443b67d0a1ace64ab9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h68f3d39c45057aa59faa2680a5cf83a7f01644bebe264229ca341c193567fc11167d1b96ab8b6c859ad0f80a4f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4814c8f7d3be67a7a8e8b7f97e72d03764ca000826980acbea080b9f2fae1a7e5856e9bf764a086f9c1ea272b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb87ddfffdcb4a221c26dbe1bf8d9db8cc17e2f754def5c6cb9aee4d81038fc0d5b63dce2d0a055600d4d17314d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3828867e00b244b1767bfa2ebb3e87e17773ebdf85efe4e1499bb73376aa2cb21b9085512ad6e108a9e9af0746;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hab85bd72b0d7db32e3e87326e18876e0b65b66479493e2a00f9caf125005c768ac7d050d41080b5eea6bb69bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf010ae61caafe019b2c32339b3328bf164b8d05112ca4cd473c23b523b830b678919033329430c10bc6854d09;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1863e150c18c6e7bfcbdb93d6503c094331ffc8175748d86fcf5dec1f66ac860f3f101e9b4b1d0c376bb8f54bf8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h68a0807012115425bf9b1775e4b3903a9427d2ebaa3731aa353d6519a616fa3171f5508608f77255fc8267ad12;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he2895182a505edc8ad461daf66fe70707d793a334cacd32e3e300955a87da633828229c75c747dbeaa0a32c8fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1869f70d7118fdeaafb22544f356732109a0f944d6d0ce54730eddf7ff802366f663f6eb9f869fcd60504695275;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8769fdefd66132e7128f1b0b51ba1fa0c9039edd846352d5ca13edf91c48b16abb28ebb7d0bfe50b977b8103af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h700aa10b2ebf74bd3551bccc31358068c86909292c5528e73b335c7484beb76931ee32ba31b3266c90b30190c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h105e4822ea30666fea3a67ba0ac2278aecfe32e95694c95efecf6aca166d25c2e87d4a3e6bbd7362093aa4f51b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb8e88ef8734af9fadc623b2c6bd285a6f773499b33a9f000c597eaec39d88b70e850e7ea348a0c77d54b5626e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a510a648fc644f0d0db796730ada931c3684f61056d64fa423caa16a01f3b92d91d8196e2513cfe42470f93af7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7e0ed9edff4dcc47e730f250ca99baeef176b899bca468fe247149754ae2c50a31355b8a0162c54638ffd3185c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h93b1f9c91ee1cffca35a829905fa9acbdec8c8fc14594d0f5a52f74729d81d905a1a590c32d0f10d3a316b30af;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h63a9db65e2a11bc2a5e59f04614dcaccd3c1defec23fd376980609371ebf3bd08f622736432ce58e77fbe3389f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd8971a8cc8e463e3881db66638ff76039181242c421499748558361375539844e912d956fb8bb509932cabdbf1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf0bdf5ecaac8e59af2232fa49d963e3eacef3eda99b826113e1aec0d3233eb5313bdec236ed3502cdd1d86f9e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18cefbf2b743c072b0c21008735c0325280e9fa3c0f8542e87688676fb6c0b1abe03434763068e52928ce899ba0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5cfe91be49dab123bb48599a78e386eed2d1ecea8f023dc6e1e7480b51c87cf2d001ceee370523446b299828cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17d6c40ab2240ea305c788edf31607bade625651ed9447228eeb00b03d724621bb32c4605feaa01a40c9d198394;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc65ed9038cc1e94a4a0d898b0a1b4b414bbb50348d2ba2fedfd3c2272677d3e4dc57967772d9b24fe2f1a41f70;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h78c0757c3c636f773d2990544cf1c7e4f3d039a128777bffb916a3d704024099ff6975197faa75efb7c9d443d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16f7d615c31cfffafb72212811b720e34958dc4effcada4fdcd5e4026f4f4c2b04fb36c542534cf17127ced3f2f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14718e591cf12f655266045d32d32529807c4aed99cccd389ba6dc7b957307f7ab0d56f87b16f2015b1ca703b56;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b6bdf39fa4644d00d9c2a583cd452f17612757a551653cfe207f30070e53255fff7a659961cca500eb5a630669;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb11d40a66952f4531b33f3c7190a307da97058b2277015894728f92941d80270eb74bc0d124a4bd7d01a5cadc0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb5847dd0543e7611ae4f278ca346a28c24afccba9ba54a6899d4f3fc0fa3db6061b5f66450cc5854376b24022;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11f361097f16b340c41c35cb1760ebf64abd6ed56fb804ed7637e605789e50c3563922aeea6adae7a1452d57f53;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c77ea444ee8697c1447759868a9e8f4d21d323f3d49119c7ab4a2907d790deed1929c0d4b72f0f0e70caed6d20;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5f2ed29599bccc9b6003f838aa6d0dc69ee16bd70e43a5403070326db8dc048b830b754ea643614dd6f0cc429c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h82108420b2a0ea2571c1c70e63861abb971b413ef916989cb7f29cdfdca9acfde8a07d0acb0c5032a1f61e0dda;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h137583bc4aa264bf9dc932b4eaa4f9a061e9306782192d9b6d4f1095c610822a66a1e3e249ca93a5abd51fdabe8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha71b7b33cbe2851702a71f295ed036dcb7df19758cba0d0bb7de833604bb661649b813fefefc3a2562d95d371;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha217320cfbf0b3e83df2f297ab504f5cc42e1fa8099b6bc61228c3866e1cd6106b4130100b69f3014eb010966d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e25c8a8f612e9ed73d06a24da04799b3ac70bdfee3281e6a79eea2025785eb5ee8e17800080fa4b4b9cc0fc988;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15c31df75da55e26b0eb78279ae80fd861e89c562dd40e08cfa366de8c81c85dc9de5f1300fa4affcd6fb7116a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h134652279086b697d2092d826317c3d8506c9394ece8ce0fd94811382073c98bc25c89aaca5ced2724f9f3caae2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14f612b5b0fb40a23f8742fa6e0bdadc16f62122e9a5d890522841f4dabe3293087007d13487d1ff28fe8a0fd04;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16263a63688cf83da5423b6a5221e9704621e28e4a4ee608a60c0442eafedcf07c010bdd25b8b730dbf39e61b46;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e98f7281f9902dec3118bd7f739470756a737047587d2aef1da69806468d6b02b2fc4ca0eec800085b4fc1b23e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e7fbb67c27affab4ef66ccba7ea1350dbe29d510d5c24068492538d4ea0e30ab931b4f2160045089055de58c56;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17b369df4b189ead444b9a9435a4d9d4a4a15479a2415be9ae951445d93e61a91beadeca5cd6728ecc1aa2709b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6a08ef94632b6c4911359d1a79650897fc9e26fd02970be7492640ae861da05527fbb6cab9bb6b9f16c78392ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d84175456984adbcce3c54cbcd7104ce95ec903d11b28b9677fce8bba8e453c20532fc1a9265ca19426b2b1bab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h43f72ec44c24c0a8047a2bc990b0424c0a705b136ef2326440ec37c07d215eb0a311f3466a336bdd76b1a79400;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cbfcdfbdf9d4102dcdef835e3eb98acf69a4f42a204960ce385df22e50b3199ae845f6114d8ddd439b3b2dc44c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11329d50e2e0e75f9d9708fc6d6c13e4bfd630be4f0c2df44c0d7326ca6de8fe983dadfcf3f74cc2cf6dbd0bb09;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h190657e0b5943f947fad9ff48816ba6d7372cef9ff127ae0c5b6975252f42b5dadbf0da1c16cf161eb7e921643e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h458e438de7361efa1231de3be77eef663215c0c2750dd1875c472c372865fa933bd5cee7f6a2f32a7ebd19703c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha8b3109015a7541d1ef5c7a84eaff3f5b3927d80dd604ff05e6633f73ca455949d2b45804c4996cb26b81a137d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ccf7efa2736a1fbaacadb7a9888fa6060e46502fedd4338126cbd3b08d2791cd679f2222512da53a2beb2bfb45;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h80eec5059e9d7ec046340b93007f5eb528bf3a2951f1436a5da40022859b229f2d13792317cb59572717576174;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdad776e3a2d5835ae001990015ac7dc63bb8393b0e5c1ff7f9a2373598bebc90951c681495fcb47e1a0fb26316;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16de39609ef582c5f0645a99e70218c68be9ffa8569fc8554360e443af15a9e9f5d95241f7e43ed5c1cc7c59791;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a11b122ab399f5df64fc60d9f1ceb0383d8d938bdbca0c9a0ef40d03950e16869fc9b0c4d15ee9ab54c23cb71d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17f0b1bbb8f2115be50cecdfc8cad66f66d5b4245ccc65bf8399d5e57201c01963587d9e03626da3c0820c892ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h191af46a80ee8eeba07fe11a90df15f3b801f75f89ba062ccdcece8bb8ac46e365d494de075b4b146f1bcef78a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f0261d719a949892628767b5742674da4266300cd9b20172182b39c2957b19c73f6edfbb5628bcbc13f72fe309;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4001ef0d304a59139a71a4afd4e1cd1c18c4edeae5d40e88dff141cea3dd9f7f81f48506e7257911edb6d98ab9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he9c184cc0f2864a9868a741dc6c51b2b93c4c0cd53b3d155c11a11251cc65944b37ce2586660c9bfb861e5c7b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3a913a094f6d34ef341b18f3cb6969b7dacafd2410d444e7e959fb8021061ac0c07e3663f4d896df8e287df6ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13d675346719b0731485d2c9d011344877ec0bf81d817af3873d1c8af6144fa50959bf883d6798fa86f68c0bc98;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h199ad28e740008b57560f1cffdf0c1278040b8619b5ac7b488feb76acb42a86d28bd71307474527d22a0866a6f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb7b4e9aa7f452e3875e6c7eeb42a2999b0ab864812d84e0b7dfe2cbb1d86dc5c0599ecaabe05e1c6149c751247;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha28ddb14f120d8371f10cef6b5d3530d6bf3b4d8dfeee7e3089b3321019f1edf7337c89ce743fdec0a2e607d41;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16b40b02c3c6f39fce7868028da2505d7f096a3aeacf8c61936ab72409a54bca2bc461dd8c1da97a8f24240a3e1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h858de20fe13e322a0693972d2f6d8c1a11a39dd45077ae6568389907c76566c957e5ad015550dd5dfaec6b284a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15ec36dd803fe9d426f0533e68329895e637a3f8979f345ab03e33d063a974a624561a3b75bc8d73531ff152228;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ac1d64bae4923583734cee0f262cfa1b1bbf565e641a507d4ac3d915c3ad0963492a150053d35944d695c8017;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha4c09635801a2a96a61ffb07b7d729254054d6ca36ca4ba9424dd54403f04e9ea3056df92bd6dccd7bd4a25dae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1549ec1866b5f8c25aea7e4ba965e2e5ad45b3fde19466d265c986a8780eca1538820b3c9542c33cca5ecd7698a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ee5d35ef2f0289be7cf6db623c244ac993af4c707fc671075d08111e142abef6481890eeb87392af1038f96bd0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1abd621a4a22ebbdedf5a9c6322dee1c196a5ea239ec95fbc972c2c7128bd4d2691a62ee55325a0cfbc3115c32c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14cad9991d68e152f2d48f57b4185cbb6ab04b4b6c0d23d55b457a01bec10c136c96cdeb973696edf117eb14ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc9e2a143fb965e939ae65ddddfa75de3dcae9ce0913db840a0765af58c941600b4df3395f7e2057cc913a51cd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hede1362e73ecbfaa1bc1acf73116a174dc58b5318e370f9d9008fb1278b3cb821c9810a076cc73bae2378f840;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c0e12503c713d3f9408dbe917f5b5c62f0ef7a1c79e3787e000bde6f5f920fdae2ed825861aa285c26b0f627a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b92d20614d3572ae0594ce55b608327504f3c63fa03083bdd0ad08dd1721abb97c15ac9a53af091221026d5b77;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c07c8a6b0c1e2fad9337bebaf7139add0e3b53c4d9de7145585919734a4c50ccd32f10ff8e1dff0146ed52735c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h160985e9b15ae6fe711048dbb1fd711293253caaabf84f1ad61f279b389e793afc0ae8ce9c8ab9d3ade7df97c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1be69c5409baeda1e2ea79cb2e7105af0e3cd10df061f7213cb24ebab001afd9ddba3df39e2a5853863e8a5ced9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ad076b0e1c0636a1eadd9ccc7fcef63a73f0b9d981d2e3eed6027ce615ff31676c3c2fcb91d855ee528a1f2ec0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e91161701873cf75ae922a6a0ce696cde55903ad50186a37d53d1f9df62f8098ed46c4b12a49796ce8adb7cbc1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h695146bd16bab0f483ff497463a38ad2dc461f7985b5960f69a79886dc814984d2681e33ba65a0c1919b0ca7b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d91f392d03c87a7fcf017ff7073df4259403f37b96aa82f67d6d95e1485b945ab5e3774fd03933e2172fafc30b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ad0f41fd458fa8537e9d8f1077ce04cc3e150354f76d59f40a03a78b6ad4dee31d9f0479d4e6e1fbeb4d7810ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fb8e656e40b9c552477aa00935707b4b2a56d11c02aaede21a0b01694fa2403b261f8d1987f72044de0a34bffa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h165a68a68126a8287b000cf7bce5a7a07b2dc48795438b4fa17886153a1ec275917638d34a2a675e7c7b3b734b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4cfa245f6165d43022c3359cc994c24062aafb40d20533898f3063c3d1b0f0450c1adcc59096939da36a96c4f3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he237ab204d6bcfcbea0afcd09071a0dfe0e1173042917c09df8ae6cbab693f38eb0ec1b1e538599e1db08fdfed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haf8a1b223044fda32fe9cee14546549e67c53bbe82f934b73f373087722080ce0998299cd6a72cd538c4cf72c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1da1d35acad4513905a804bcb36d259978848b0eded7b52c2c655ac868b47d1d9511b4b93aefdcf88df0570d2f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d440bd3b5553f0147016d7074f8c3280d70db8dbbf9017bf33b70e17b5764429bd7c3116f651f6fd2d6db42010;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he8b2f1098486dda0629f887cdd2e651e56503b81fcd40ca2489aeb22d94e1b99d65d0ea202c563bba983e6ff9d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4e43475da3390dbfa6f7989da5fbf0a950f7935c5c8b5e9ae24b5a25a7052473b484c588e492a833c0b874857f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10d6873fcb9151e3aafd216b7b0e6376cf207a77409bdae3733be7c4c2b36b3a0f29a5bd984fa50f2c01646fe01;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eddec6bb15cfe39abcd280ccad2d0b210659db108529577f6d571385f5976f5f109745951b07459e86b02524fe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18aff4482c6596158331152c9f304495dc95aed1be45877734a775423e371a47c5bbd15ebbf37f1f27478b02134;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1419f270c5288deffd1db8e542b4a0156b00b6f837073173bd7de248ffe5fc85d0012a17536aa64e4bfff396ee2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16271a9790114ed216c93541e829d7757b55ed5eee905c336cb534936ba9259cf15657d15d5916e16a886e2a426;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9dd7c84a1824a1052c5854a113bc2493a803e7c9959fe82911afb5c258df45e963839dcd90db9c9b3ed5bef93c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19305d2896dd7b28aad242ce900906bcd2718f4885b1d5151c2ffc20672c34b0a0aa16c802607e989ec9fbf29e7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h127594a7270d1a0815af54dea0aa6373e56e343728398f05d02c8b7435846cd471eaaac76b4fee40e45ff1cc261;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1150e8262b4ac1f86d400b3365a34ae4fae66ddb948eda613c57545c1a973f3320e014f4a155da9a90b834ee5ce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf31690e48f28c3bf9d8e2f67738cd03092dc5a5ab1f933b34ae33993baa46e3fdc66555eff5164ba00a3dabb32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h161d16fb3c28cdc7a07d008a00b1ed94bbec471dd34f5e429299b14ef41b164800b7f1cf03191aa5b6accd13526;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1186be5b2d3e451df2177187c27372d0f3fbfc2cbbae03cb7d852a45eb80bfac7ab8cc3d4c1adb30d45fa7b8e36;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h172d50f1ab3b52b1e737cda0f267fbfe7f4e4c2d237e4e086f104ef949048e6294ce1c776f97bdff801b2636c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e17c67932de5d31133cf9c46af682dc0da302ae5e2dc1a52a94c1875f9b19d630a8469e1a598964710fd1887ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h940cdb3741c502c1ec6a34077ead5e004dbfb41fabbac308677b317491797f4075214dcb421906ad2bf2566a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e9ac31cb94ad1376186bf0d7ac90029b64708a475623f6d55e10bfdbd2504bf9d21042febedcf03c760e634671;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h463340d35ce2b61d7aec346196da27d417ff50fd4f53b85e5a5aaf0edb204722ada1045770c707d081e4e4c3cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h146399430b60d196da6aae9a8a4f8ed8c8c119070b8d19aea7df2fb1392b2f5d0ec6fe7d1550d169c5fc8deee37;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcd97959201ac89b45acc5d835081e06ecfa92ac880bd45b2bbaae6ecc6fbf665e821f5b3ff680adf937e15a017;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16bfa602822e3f7387e025e183452a2a56d1cd7d1b4385f8bba4ca381ad20b62480112b2777d42459ba18d0ec7f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19f256972987a03dbea39d9b9cdcd27827588e59b9cacf24050b9c92edc67e4791ba4db2634cd4af09784eb4fc4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h58fa9efcdbb81ada74589214e6eb1663fe146bbef97a574f83970f78ca3787b111f6746d7635f868ecbe8dfd69;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h468e02c14e63af376795b9c7ebf8edee9c2c85ba31f736dc4a2d270680df7f2b0a9de63476ab39fbc5ba8b9285;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbe0eeb8c2b8c273828dfa54a472f6d91a9fe12cb74b02ea4b7afa0044028b7f111726ebc80bdd86256ac7850ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha104321907ad6b5e6fde61dd335c7dcd983ce670e274f9cd043480f5604c70fbd68239e8870446ad9c2df2d83e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13cb5388377a38dbc7a738892ddf9559002e3d8ff2e8befbfe848689c9f66b7822adbf5fa25b4711734d29b6e28;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha8bfc30b9e6254af0c0de558e65a47277de20b23cf4bbc28dba7244529de5d1fc713140c0d75ec9db7c5ce82f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e44a7ff55f1dc216f99bf1ba99d8ba412dfa0f5732a1cc6dadb9d64a326cbbca7580f317c9ac66e3f51c2c9bfd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he4a112ad210bb6fa3e3974b7692c17b370ed340a191d5991f3d1f603033ff9d9e1a8f2798c1c153c4694998028;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h487281b8121e2fa095217b25c8bc2455892fc4075f275e7daaf9dbb9b2156075f75db8a3cf7f0f889c2e585d26;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf6bfe6cee0dc745d2fc9e3e72eb9bb56e0948ad312ce20d8e9241c75c1f9026c327e18feb899e9260cd2915e7b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcb7a9eeb276df963196a486b422ff1547844871971ccfdc22cbef75d7e44a57d312dca1a273b86b6ef74b2179c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8eb216994e37a16c7bd042658d20df5a8af3371c1290acf6fd3fd840214a452fa24d39d4eb1e37ac2262bd1f02;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1065342fe597193885906ea5bf59f302f43094a2d0bbe258dc100ed6711ac5ef988c332d5fc22b3cd733ddaa9c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc98cd40b1cd1ad68adaf6517f3f25abfa8109871bc712c14302be856fdc88356aecb7035f41c2afdba74b396c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc4007f1973921e6ed3d9b82377b8e55c4666f4c126b4f3e91025ecbd9cbcc60923e5f9926a37b6e2b3023339a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19783d735993d1ad66737b2618cd1aad567fa41e9a257d8f6201ea3986e1a02b855bf0ec23ca40f65a0c905998f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc4e7cd21524942a18cbe0c2529de405dcbf0cde2b978881606d74915d20d9d7a6337d61d2ee3d1d3b11239ae31;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cad63a0e8ec05d7afd43f9d1c6804e97737844f786b2b92c3c68e88e0452002af138c289973a16a3ed00810c6d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h122d0b9c8526b5f33fb81245268b5a323eae56f699eefd5eb9cd4051b6b30b737dd29b33d4b25058ff70a10ad11;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d258fb63a71d07b3948a765ee4b48cc195b3ce8b48923f25d386ad9b1203687dcb021c5d0d82a7ee204e74c879;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c402c9a8f692f32490a2684619a024903c0e79132498e4e447d2d3731d9edf505be306de80569ffcee04bff3f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11f1262901df0e460ef4e5de09b5addfaa2525a7f8e520da5a9dae1bb0f31d56b80d86b56545ab34b9209c7719;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h133ca3be106c818da6f33a2b6109fe5ca7eef5975ef422e9038bb570d20d3dc3c73b25cfbc3f04254057b1ce53b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13bc75113b8d11010a418055f27e918d5052215a909c518a5a7803ac841f092a7cf5425919b9dbd6cdc3c86040a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h186f6ed4fec202d615935ebb2e2399486ad93e785a957be47ec71b9c7faa0ae7929975f797aa6d321b7469f0b4d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h42177f827d6c05c3e2aeabc4173a4cef0c520b0b87e3593c5052b5bdb26cb4ec26e94c873768ee1b43ebc31e9f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ac3de49aa827063da5f37a58d80f66f4e624258fd19b489375fd1f06b720a49140c578d9f6e4e8eda52c71b75f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f49e013f7626e97307b9ab7559ca82c60825412cab50eb3a9bd89ea766b858eff9ae292a2ee1742f7bbe4164ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h34f0f4c03fee0a7dc1cdcb9d1fec328d1e8a98cd4224993fe629b5f25c6dac28a745a81b4df9c03ea28de628fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h125ecd82cbfd39d8c0fa1a0c47203e25dfda9822f32e52e339e4fc707199b9ef331c1bf9ca8f4fb992321def0a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h89cdaa606be6934f413ab88fbee03271b6b4e68b439fcb7fc737ec8eda69105ee021c9f846e5c55b8d9284983f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ada4cc9eb505fba8ca087f1804fe9fb9de46d6b88f22db3ffbcef409d4e467838a369e8d87f93d6956e7e8fb5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfb4981eabe27f1751b3bcbed607dcf61055ca1491d9df8e02d0e899447ab7a473b80db53b3cef43f78476ac0f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bac803a2ac3b5f8299d03d9e76519de3fe3643feb62636868690f5aa1be48b975419be32f4b9996b0058cc2e97;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f39913029e08d7e2e062e51ecac65b9c3eae0a0c73ae891bdf407a649defa62c459ec1071f185dd0279a6c452b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h108a31caaa6d3dc1720871fb31b8afc0d6a9082875e1bbc010dd6df3d6dd8803b87b3cd0871906d83a1734e07b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e89057cead4095e5ae1fab56f2e31b23b69548a5635ee01e8e7cf0d38cfff6bfd8e1b3be6a6b278e8e55eaf110;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f0a2891b90ec7988aea9f9d7aecf4f7aff9b8d2bef8a17494454dd5b10d40f7b4d92d6cd1b447d4355972e33e1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h161abe46dfb6ab41c25159c6fadd95b0d395306690c12a5ad9bb6aaab32053eaaa2ce13a9fad2a958ce2a812ec6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1914eb1f7992513a5578f048ba81eb2780a4f4368812c7f1de5dd3e76b2dffcd1aa81b814ba9af6d94858631bd5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdd715905ac88de6af66fb6b90e24573846c8df67f6ac008348dabd291d907372df6a87260239430b70e742d873;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd6a683b8f1a5c54055ba43b17dc6a7583bc9d13c5833a0cdb13f86e2a9b2e7177b542254a0b83e777b21560f6c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdef216f048ddd23b23731baeef8f6793cd084dc6c79f4f74324ea81bec29d05339834298495325043dbeedc758;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h111f82359fc2181021ee948be3c26603edd1df1b82731e7e86437b9f291d6de508430d57c5c7659cde62b08a247;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h22dea180ec15f79324b7737655b38e1ae7ca4efcc93cf48aef1c17e23dca0d8d911cf3c86f6103a5f9eb094ca4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c529bb454981871db908c94a393ec9f336145623e60ffec63af3ef92a9fd05d1766371f070523c52f524e1d448;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fae630a3470ee560ff34c818c4ddefeca36cbc5721b232acad4c91f291417b5ea69cef4af07f6391c833d9d063;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c6226e70c932bba68cfebb3dfdbb0f83e692905b1a8d0a0ce9fa4b8a47a27db1fdebb87ab97c3ff96d17ef3252;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf83db59685e5e3a4b499b3eb3dfed4ad9430d71d026694dc9238af0902ee6ea60f2aa4debc87b94201b105fc2a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h271971fa33bcb1b59872497629c7c5a2a76047383eeb0c4f60109c6cf4d3c2a555e784621b2237108ae86af106;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbdfa6916885c8a90157202b0355f8712c6b8b285f4b6da2e5e38a7630235e6a0bf0ce69fd8620c36cada83c4ce;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h156fc47b62055b76e0746343fa57ff558ef64491459e379ed1cf490fb1587952c9ea86d86e249cad6e7105510d0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd3835c2377ab606565161d46274e9e22ed68b3e4db9b2ed50b9fbd0a0a620f2a9da12dd0e2d35556eab02bfca1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h128f1884e67935eb014f54c2eb60989094dd8142dcb35069d6243be7a820ed3ec12802613e528199936e4e628c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h69c266017d51a6973217b34412985394e1755494ddc3019bc08e1d811006062a2ac53891ae0ac0d36e459657ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d36f9499a497c31588fd2ea3a9d3b91745cef8cc711eecc3395af504a4cb120171326c1e43bb09b41c44322a6c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e5df9bc909801116f6f8f1cc18574d29027cb6865f4110507538032019d497b134e0c7ec938e71fc96d909070f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h55b511791807d8422bb39eda064293d99ab7dbec8c1a0a7e0c95191c44de69f8fe1586f936c45eccd08408028;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hef21e9b5af6d2e9ee4426b41cb3a2a1450907f05cf4db7418f6384e46bead67cbc9bc7f376def8e53680af49ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hecdadd254d605c8cd2d14b910713e385620e88074ab0b283e0c063a5bf90b8e0f36147e7a752de9a126c3456ad;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb4c07c330ffbaa29bdbad34123f26e5709012a0976cf2eb310ac69c45c7a607317ba9a7b1b53f16556de2eb1a7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h41060b58a2d4c2d44ec716b6fe2a6e65ed53c8726ef4d0bbee00afbc9e235c348a151f6af037aae3d684de7b15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18c298280cc7783e90c468c0a60ba6fdcf70e55ff248c0aa433fb88330a07c5a91f85b72f4efeeffd24266738d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h120d550e532bc078ce1533f5a629ffdf951836aeff6a6c81754991ce8bd6ae1508579fc8e9df746abb0b065a60;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ab585033faea30972128cc2eef82acd46571e2f28e08d6e423ec0f39495bf9ebb2848f31a26417f33920726c6f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8accdfffeef8fe36760644d8a202112b2ff6c2d6c80a91786862ec60392fd01c2c50138e807d2560cb5f59b802;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eb3b9ad9c96b62d32cca51b50a09723f1f069657bf7fd7180393620758ab533644210f87ed618e454efb8ecad7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9b6c0d5a2457fb89d8869ffbe94a0afa348f00d40c879a1d04e3fa0632c82fc2d158857e6ac4ae416e01b95557;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha1a1d0931bfa6390e179dc898f7366c7900bc1e0d0a9d738210356f79bc51c31a548d05025abcccad66d93728;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18568ef17e2e4fb393061c413f16f87eda6ea21d2e6a68ca6bf3924bf11cd378039f63adb205ebf5fac0e7786d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd146caa79bc3ff952aa4a9e596848273f3ccf9398fb9a4984de5b0e1ddf8d8a582e33e9b0c1a9d8adfd085cb3e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h35baaadbc17b9d3decdb3f427ab7c29c6737ede1751a22832516c6bd05aec6099889bbdb595ee4015d3d6c2cf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19662b3cfdbd646853749be5d2ed97a1ab326b5e887bd4a4fe66e6efff61e921ee5461307b5181bc13dc5ab4246;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h811f9672805b3f17ac5bde6d73bfd52429d47cffe791b3f86b3650099852791defbb915e9ac859ad9286801873;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16e9cebe4649b0c983ccae591d39ee0bcbf0afd77d90b876309ad5ff00896001cfb1491853bc0149ef64469d0e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h118f9e6cae5004fc2aec556a85a7c8d57a753a9a90993cd46b66b79de63a4614e1a3a64a98d9eb082322a94553f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9da8a53a80ac6547329c43c73a3d670cef9bb4c1d90b061b2290b1ebf967677c0a0f4938fa7a21451f229a5dca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h338ebcb116fce94389cf97f51a1dd0cb39a0dc0ef497e9e028022dff29b110d51237eec56ba22c1942a734350a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h138409631fd06a713a9250dfde380e49a74143e8ec95fd63363a592dd815cd662c823fcc7d1303c92a0594662c6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h167a782e8ce534093d8777ddc7fed3b7e2c75d0eca5cd1fc3b61355a5f9328a2b8bad736609cb5a2fd280c1c135;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1065e3cd2e73287b05d2969f54cd0a27b257197525fe1c5f4343d0b538cd32f93a7a870020e504876cffdbe20a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h570da203dc19e947fdbda6c8f8438894b193fae031235d2d618cb1c30af59a5383372c9caea9ff125e022cecef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9de4365e8b1a73eca8763c6f71f62c82eed2054b1837484bce5515305b3357c0f7bb99b2356694c52dfd6941;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc67764c8d5fce38d249be5131f7ebb431e8c982edae344a73e5bfa335e59ae8cb3a95c24d43471a8ab51786d89;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h78dbdb9e921dc41e429fe830a67e6dec77dacc0810cd480bb24b9d347173ae6613a8571bdabf98f049996c8819;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11bc50cd1ded57b3a663ca813218ab9311cb5aaf1467adc23a2f59d7a8315032557f2f4677f7fd66713a4c659e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18ff7bb372dcf0f005ca4650a72b490a19756b2cf5dcf64e6c333378fb6f97dd81c92de5b24dac7ebeb1951d4f9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h126b8fe35a0942010be96811e2aaff5260c5d6349e499c693c945e43af41607b6a27aa8cb909a581a71fa3740a0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13bc1ebb2d24b52b139dc497ec87f212685e28aa35c26cdb48b2a9e035e1f7d1813cd6acf2735ce5631df6201f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c5656dc814164b12a6b87b65d8b4969624eb801a9790155eff00d4ea138a9c460a09de0e214e0df9884266d2c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bf6c020eb221c8cd5deea91189509014e72f2bf9fac2ee1792f4bd520576aaf5d4de3a1d39707dca2c5efc31f6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h36ee982b04a8b979800cee119bbff5ffbbda1cb9f8b12f2d3b89efc4afe13c2675a990ccbdb4efb95ec997857c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h168edc30b2e0d57c56cf9b3a3f56e0babbfb802a5d739451f234e21a3b5ef5c6cb235b3336152ef1eb0b62af3c0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb2e7eb632da913c62f0b64b9c1ba07694a81494749639301843d9ecdeb40f49b9b48835caa9735536329b28662;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h121bdc193c4c2d3c1cf954eec11c2f89bd90018eca6a8a4713317de2aad61932c223587fda80425d5a83921249a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bdad233c4b0f6e7a4c31ea6d06b036c4387e25ae9333e05f11de9fb0afbc6619339a993576d4814b926230caa3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dd7cc0893b96167c4d5d805adc17db91da1d40f1297f7d7dc4594f96f55bc9b239f3fb51963bacb6ea248c87b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h168174369db11e048025f49e211b4e4ed1dbab81925f6f24010bd70dabb26547087e92adfe6d0c6e7af437360c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h47e738e95a71929c99a684131e6789b2dafb21885b12e7471319c9f73806324bdce7929fa514b55b9c1297c70d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d1238786781dd588e12aae644425028b76e59928a85c2fdb49cb36cec34d48439a320591ac10ef636c0843f212;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7ba0fc9ac3d3c241ffe5ed082ffda15f494ae959341437d7d1c0c6b714186e8edf0df31a268b36091bc6ecb2a8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14c706f416774b102e74a194c74607a5db9425bd572a8d09bc7142b8a0316ca506f139c7323f96de5d0760b2388;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a75bd3906578a435adcbf1eea0fff6447173a7f6673e9af23fd34b550d60bd33897c8131c52d613fde68f86442;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hab685a5210814386f64bb5e27a56fb73db9de876600ee986c313fe60dd48cff6099e2fa3562a1c37406143f53c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12315a88640b01ec6273b466d52d94fb6e7ff5bd22868abd26d94b164adcfaf5d460f04c327ecec8df3533bbb18;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h475e9bcce71b2f195e8207ef0fb593e3aeac6b75bef90772851aaf439522ba53a1dd852d4259f8b3576b8b0f23;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10d432d396d8b4e1c0b380cde5d1bd1f5f0dde6412bf17a307cd8ce6aed72122bcf3e3ddccb89da6f4aeaedbccb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb5ff1206e009b70708096a6f6c225bd15dff93790dde25d48c0ceea460e7b8540ba090726a0c1b29c980d0b06;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19da58ad9a30f10f2e5ebbf338016f55ad10b47c59b86060dc9451a3fd3249e0582478f001440f0aed22ccb512b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h128ec5758b35506e43dba5d2b342612da33bfa5e2e9869c7a2f213d813e107dfe1650d2ace47d6fe798ec6a4534;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h121d726f00433c6778acdfcc587647a1c26a30d6cb779d0c8885fba1d4b1f0e145be1395478e6567561ca925ab0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6fe160714b644bd78cf656b4037acb3fabc42a903e3526b0d05ce5dc7c1892337dfcd9708874a115d0e32e0bfe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha48837112563b0c02b775f17e66460c5697495632759a1988a42a302eb81a307a95beec528aac97782a7c4fe21;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14c8cfca6509eadacc1323c51c4d8939a3afa2731812f4b66724f50c8675eb401d4887ec0a76327d5b62c715fea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5b20dfa0e3cb7728907521e4bbe20f5a2a29beb71b7051095823c7414b1aa03bba02d0550f9724f6841080672d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h60a5afff7fa4f1416d6aa20e6a7c016d5f85bbff05a34a836e24e83e2a273466af7187fb9893e0f309e0aa5ada;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13a50d6fdf4496f0deedae5664671d37c6ee1f59e6f203f126d367c52d1795897313a7671e8f71814fa398e40d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c1c1ae03daef119cbea921ae5c6602b11d484c918b4e99e9bd35deefe767905a9e1e22ba983dc2ef237488db3d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10bbd636f496ef5161bcb25d84bf514cd9a99bbe8883e2c9236a0a28d94ab4f8577af7d9faa46c22797e3c78b58;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf4c6c5d6c4a27bf46c5c78953592aeec1cf1514f8f3919723824a1087f128ee883a1fdc99a338187eff1e078f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3cde3c5fd2f45bcc14692d27369473a63400fc8c1032692a2238baf4bf3b8588c03177f633139e1ebb06e9f914;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7e1fe20cbbaf7811c6dcbba6d175f2288571f5641d7066b1ceed7dfe60702c9b69b26d23e5d22283dedd59169b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eff3cdd08efd315a5623d845dbd3634ff36938c7607984a853867ab6a6a5f59d2e4af8e8a79c86d915d4b1a341;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h70b94513ce527d3fbca59c5a1f7a63d025a3e5b1e4dc1bd516e0373763a7c08601d3e03b5735bb81acf668d115;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc91fefbb15aadaacf7b3686d1c6c9792b507aeb888c3312fbdc09564468fc4df2ea47a428f86b28305baf86e05;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9553dde51c6e6eca8b010793e144ec5d7b5dbe7aa3e5fe47c24ebd6763cfee85d2fe8aee9ab13fd5d802527e3d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b079bde3e328902b4f44bd450a73473ac1f1f9df8df9aae8b46333271538e43d7d5736c3e9e26eaf01f65deecb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h442a05072e639b53b5e2d764b94c65ef6587fd68b8ffa8ddab858b623d1e06468f28623efeef34d1cca18837ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18fea02dee38031dcb2f5881e6817e41dd2458aeaab193970b85fa196caa121d95a8d89ca6e690ba5227a1c326f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3eeb646c5456ae96a0a053afa1271c930f4ce196965cd975e38510541db3730759aeb567a61fc23e3880edcb5f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ae9622fa50e181a842b11441e757c778e4f35afbbc1ed9cdc7b225cda8bb2d7b5fc09443365914d618ae32e2d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18d47c82bbac433f8f2774182194b57a273bc97de7cfe075beb05cc09bdfcca47d231f993f959623b6fc37c5481;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbfe72f030e383ebb723895ca44f5d305c6dd1da13776cafb93112c6b3c2e314d3ddb826a7aa694858fbb03a9c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h178b35c43d49b80728d2a69be1c4e5492c8f235ba1d17e904d368aafaeef1e9149aeed4d7f652a0553eb081cb87;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ecf6e78b943861f6e6544c6c5a9bcb111a6fdebaedaa4b19688e4088ce24d59d795b15cbb308de5fb543598225;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13288f893ba6f527bb8e93704e5647dcb7d614ce9a68ef893564d8a52de58b1c6ea9d72585f79ae6d9e33aaa1a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7ae07d61d22d81f986710bfabab95825f39a6879280bd7074c5cc7cc6857dcd39b14e6b2d84c55da2181d8fb68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17994b8d9b0f3e2a173e4fbbf496fc99bc6f26de98794ac12152e106ca6002d5304c5a72e3fb0d9bf4632e60da1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f0b6c6cf5b980110e0a47c9b32f46520e5fa31489fd17a016091f6e1295ef5baebb81181fca0a6d84455592e52;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6862fe9332e2a6b6774e98b5136282804dd2c08a63d99ec000feb510bcfbb8f34f48f831b6b9d5df5ff5a7e800;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h142ad750b78992827f82095f52418c99c36ede2050cbb13aa79665af42ec5da7f18b1e888fe45391088eae00ded;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3290f5e7ad3faf8be3c62664aa9cbaf0e9c13a93b48d9ffb00f0ff55c46c43ab7dc87bf976f7bef7cea5bd8802;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hef01f04edb5c88952c38de9fe6f71531fca27ca66325317ea553fd29ea10dab27cfe5c249b939e4ac5c7faa1d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h110e9ef4537863bf7fbdf9e0e54a1803445c023bfa6a72d74ebbd252de9c6dca3a54aad92b4c620a7750ea87c27;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h412538cba79facec9a163551a930e95bdbdb344f5697571ddeb5736c5849822ef4135c7424a6296ef3627dd8ed;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ee77407daa7d0613147f65620227be281daa49a5709a525ceab2fdf0cbdbacb8fa9d489c0348c66a11d058b9cb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19370c4262293e6e65f8b8711b349c3e34840f7d39bb044151b2b8c49adc4a8d796906357e29dead79e000ad4c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b4e391c1732389f76863a18b8c4487adc2498b18a0cf63604bae13b215b8069f28371d97a976dd61de7d60be5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h430ec98cd7fc603236a3227d40df465c1db1830a4c5954b0915f5d92a0f7d285ed9dcc8678ac12fda9a126ce56;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcbfb7710b85addee5262dc4e578be715f6f8579f8cfce970ddab973ad2722599f78136d9c0b691f4f64aae4a01;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a400a83cd78c03face77a44888b4ded712fdb70b941218a756dafc7af175687587d391e58e1cbbefb55c068860;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11ac803a50cd21076cf64c57da31b8dab2042852fa621e1cc72e82ad94cee55e2f81c6427e72df5eb9383b5db94;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h34fc0ffc0b06043baff15432251ec5c9ecf0fd4b32fda3576eab72007aecd31b2e724f939ecaf559bf03651ed5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h133f1918ae70501212954137a04466449c6719f4edd63f4fb3f6e35fc35ea1429f6af2914595c8a437046c45dc5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h29ffe07009507eb3de839f67133949ba560173695ed8eb4725c9b09b42ca2043819727d26abfd84f7dd5091ecc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d9660b42e6131a1361547a11840ff5e249083e11f8c77360b63c8d20b050689cba6aab937e5ad26531ebf38714;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e829f56d432ffdfc7adb7649d81fc850121b5b0cc06590e545e638428a890225f5c416126e4e5e0befdc21675d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h78ce5479b3cdadf230a01de473f63a72da0d51b5e37f7abd374dc0ab75a3ae28002828cda802fd072cdea676a8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7aabb857c491cc6e21a0ccda84388f2aa100b792875c60cdfa931055479b08949436d076891c9ebdc9dc36ff15;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1be030e1040ee136d2ca6d94a87c33caa6fdaf2cc52895c4c00623946e0187f912ab0aedd2357db03614ca3cf86;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hce1c46e786d5b94c65d481cd91cbaf1c896d6cef0a662c60365d67d28d80ebc786c7bf825e5ad3edca979569a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1366ace46d3f998796c7d20c5896b402fb7bc8af04b712a24c8b877f43043e5b6438ed402072a1f39414c09d56;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15f2bd8acefea72e2e757278ac01316817925f491d8344831c957c39002d77c6f23fd0d312941e27e8f94348057;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb13dfbd155875c2193e17e5fc871d5008a71194e8ed832a5627464e631aa293b4385e6259476f6df2bce6ca85f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h116f6503267484bc16215d844f3e9de68727a4e2d976d71ee49408fdcb1dae67cfe7266654e765dc07868ff03f4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12dcaf7832372351a1170b3c862f51cf91d4cf6b6d7832978a1bc752d1e941531bb11cc7f622638be04397fdca5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1906bb9db34cc71bbd7bff26eed69c6605e13ec2374f504b5593641e6ccbc9ba36865af82f9d6d29cba696b17c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e7cfe18d7666648fe473e2db9fcb7490fcf2238a71e88811c2daa1db421b5ce40eddf6c0130c737d42a531a466;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fad710af68af4e486e588ee82a9b1e1fdae16c427d18e1706979de5024c76dde6c95f583b0011f883d55edf376;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h70b98aa2dc6660c6c88e281a7bffdaa38d04e74eeac1e435ef08eac4fd5832aca78f71ff3c6582a11c8894c4e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h250e074efa85e9cd495ddd6e768b7a745373641f17b62ae643454f8f67a799570515347341ee763e709d679ca8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5188677555d31f3c9baf96b6c61d33e7629b86bb055d66c3ad9bbd4520d249f81d44aa21cd5556a18d4ee2f4ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h28db03646c26ed5e3b76993b58e32ffad1bd2b27f9152a3d99a3011d3ffde0999f7f7f9765a76bca9789759c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b314f466235320d727e63a7e213367f9bb95449eba4832b21cd19db3ef1fba3e455dddf81bb6da6ad60f01138f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h120a2212b5514d0d146b74c839ef8dc5d7b393490ee78f27dacedc3cf04e50ebf44be2fc5fca4035e9702cce3f5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h160b57e4e89177795c1d2bcd2b9ef7a04108581deda053dd3683289937aa183036e65d327520fa83fd21c7402fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h170a7069c2f727f151f43a7fe19151c074a40f1c4ed866dbd02ca8f66998383192cf4f2a93344b569193abaef3d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h101bdc555b0b38faa65e21ad8b2ce4b9d42a63e52be5a9c0438dd03ddd8f35aa66b2652e7e9c4fbb6d385aeae95;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b8760fafb56112876f5c2612828433e31c5f29b46dea5471d04deed58278056d48b19d826dda086ff464ec263d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12a2e4f225be60aa504256a2c1ddb0a1c829cf385b71ffaffd9d3bd3e2a3aa801244127623a449767bb3c15607;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17376cfe77d88374420d191b79ca072da96feb63ad0ef0eb88659c88bebf1df0b8857bd25962f70c1ec94df30e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d482611034e91e4198333a45b61b30b59ce12e7f8669fc84499dcc6ffa9cf9ecfa9f7ef3e50e61ed67cbdb946e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16ab8b8ac474a705ca8c4a955256d8773047c5e27904649f6c761bc324933b0088b079770e0efc8e9c8c6462324;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a8493d4a56cc224b5966f8e9c686c94c2761c94a96a50e5c08cd182fed4d6a529dc3605af47ba7fa1af2c919e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha7774a45b92d3468fa3758c09fee07904726971b90b9cdfe1f066abc7f3ccf3a0db00d9fd208946978d52c877e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h160c876e58b4f88d5f958b014fa81d64bad546c9b064126d1906d957c821ccba44367cc98c413404b63852b8eec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h908100140cf647b78541969d252b622169f57a6156c83e9ac0cd3b713646efe3908af027b700849c63a97e0f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19dbec78c2a4064d819185847b575830c76ea3d3f94a2fc56ba340faeb68e3be2b64f9e63bb72dfb5ef4cf7089f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9e8f06fba720f62c938c520462a374622390e0a536a6c7c8519db7298a0737a4dced4e1c47809231ca5716ab32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h142e13fae6f426bae8a261ee79ec3def2c64aa76832dc84f9fd16580358a0b24e747db158e18c584b2d90cacc5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h196a39dfaabb6665f26844e0779e8a54c6e055ee9fa4e7c38ce341d4fbfdcbc0e42a7a8d83669c8e49c0c68c8f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1209f31c69f152d3fd30742022fed59723f3f441bed00d425ca50e430c10ae31e9a02f203277f3e67adf1a92fd4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h26d0d32c7c9e2e5e318ce06b75c28360becbd86dd32d3fec6f2c0672374f9f62095672b96eccdf7895940ccf36;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdf209e1fbc6161b7dbc86f5cb76df853bcecfb2e247d158c41c32181082046f9ff29002c779e233bbdc3cb22f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12ccdce4365404c90f6dfd04038c91433dfcafbdd9b246faa49c16869531e5eddeb8bf15ba399082a259c8bc6b5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15a6873d16ceb9a532a15e912d833aa569bc5f5ad6ddd73e44e0384f7489f17d3c484386c01b39cc619fe248c66;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e8845584b0f061610722926ad234f5af3713d26b562e8337f8a1ec3ccb560980bd78a33668455ada40b1892098;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h110353d10b0f3a84406de6785f843936e2454c8971251db446c736dca0b096fe90939583b1a92778cee1919601e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d763ee26e066cbdd2158ef8d0541d82209c5aeb7a6ce9660e02a1a63a09aec2661687260c83e1a2f6ddb1eca8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ea58bbc8bfc50c8eb14a61d07c4c3af9693266fd23c2942d8c0a35a6c058c7ba06894f8c0dcb3012e36936b1b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf7e3a57c86c9e557fa35c750f3de5a47f71b85b47b7ec0a3600b5839993d6512ec77c5fd8bb524d8d1f6824d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbaf294ab0ceef2b7c81efb8bd9af694c2824e3e1b99f65153053ca3d8d1ba8457871443aee7b226f2758e8d10e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ccad4b22b0b9255d43b4af67a3d6aa79d7aa792ba16ab6f735e4c1466910543020131cbcf6a875757760a2483f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h122197cd00bf0aefbb8bce13ed5ad461b5651a08ba75f6cb5c2b0ea587b5a87e68685b1118cd45ebf59a1a54f69;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd445b5f32e14038328e55688397e85a315ff1ccb52c808f6462057614b70fbe3aaad241cd326711b04dfd25fc0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h26a4e7305da91294fbfe161610f125663e30787b8d220308b7ecd4d0ac1786d822f8ae34ea90b65815d5859da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12e67fc1f6c60e7126ba6bde202961064fcd5555a747dac57518c51e3a622f5005b5dacbcd879ddde6b01e5cd10;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h27841e8e47c42312bff31ce039dab4262e39440a015dd08b57588ade57467ede943998176525946e94bd98217f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1856731bedd45d6cdce26068c27cfe8186be9c91b73ccbd9dce95760af56e705c74516a83c78655b4e882d9887;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2db1fc6a45fb6eae929f411c068692ba30598c061ad46a9a01a332f7bc8923c922ce1e52dab82e5f1469d26f6a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19d4c364d21ea7b8919fdf32eff83c2f873bf9d0feecb56f78af86abbce8856215319bd543fe137918e896288ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14919f42a0933794fc72f50fa49792df94fccc7e45ae24bd418b2dda08d2c447491c1e259d5ed98ca006e788737;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5a4ab6e6b7d2193e0cc44567179cba6bccaff70a81cad29a07bbe6abf705c9ed12d373434e67125b4fe8b75ad3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9f0eb8596aca4d116cefe4c1ca6a4f6852bd553782d555b0d3e448d92940e17ed42cc6f6f3c2268abb9134763b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e0722ef6ddb4e8a230cfb2b948128870a9e5242af519580d9b5028ee31cb267b5eb7c3058e2b67aad021918641;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11fe57fcce0f2023458a8d0b2e2ee07118edbc2e32d10c3dc16f7ab417c99ea0cfbde249297593f90a7450bba47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1db0fd983d12817f5e775a312cf9a3f711b6d031c5e5f7fa36f9a87b78d86121a22a726089ab043a13bcf2eda91;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3f51560291ea195e6776720340aa3d310b8c0b88c03e5992d4c76d74dec60275c240791f7e0795c88452ed351d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h179bc9fd2653394a26e4adf70abae13e0ac8eb470a2bd12451a5c28491483f031fc005773ea74ab2790bf42ceb9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b8bfe7ba6cb0b5d8494d1bcfc950becabbbacb937b67b300936a7dafed2631e77177dcdc0d7ca4eb1d2bafc148;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h191a883758a8bc2338cab3db57c17c6bd95675631fa75eda576205d084617ba5be09eadac418842b06dd7425143;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h731ffa39ea728ce907425ebd99124b9875891afbf3c6337441e17c4fbc570fda98bb943767adaa533478ab0db6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7c67f3c3bcdb93800abdc3108c613243292fa3626f49dc79e5d212a1bb42430cc90ec670c9c6957fd3e4e8af0a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18cdcfc2460818266712dc06488e4ac479966d8cc7513ea4becb6a1a3a2de921e9f738b7aafb3166061ef0df1f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b8b840c13bb3978c54bd8a349cebb51647f46d8cfbe1c931f7cfbf4412aa662438902f8c9f8c03300ab49b692f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13a4143339e99029c8134f919b245d96bcb64375123e36b93bee38acf342e24a8df352f933dd03f12f420406a90;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa1cd342ea114a6ca46eacd685cf9ac6a9a43aaf33ea009f46415a4d24c8f32bca384ff2f74a4b2c85aae87c25;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6f78491dff150b16996ea95e42b511ff0e97b36a224fe6e22a5591aa313718d6365a17e1c29eeef4abeb477f3c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h128ef3684db6ec3beff2a363ce0fe654ae9ef32541be883f2a86346c710f99ae8e2029c86cf80853e9ec0fd72ee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10552a3cd000b51f41c957188b4e5975ee5f0b59d8de889de851150047da6cb09c70eb20ba42f1e1dd002106180;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ea2803fc48940a52870f77c6915322da9484f317a659251e58a34dff2a7053d680e6ff50f8d6b0306cc3855708;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11aa629ec333d200aae6f99472904f52c97a8a0aa7b4a1d1d04ffe1c626e6a2f8fe8c9f0de8c4200b450d432d84;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbfb2ab90fcaad6e45d923a59744556fa56c46799269f38314333e11448a5ee5d6b3b2e5d115ab7cfd11499e61c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hda1909ed749152f171c6ba034a08da6f23ba4d704a20b80933ccb8ede071aea22fd86b0386470c4bccf21df771;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d4a27968f58f1748ec1822a4c5b44495e388cd6d8a62500a883216f2889e7220340e6a839c4b61e71a4de3221a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1af839c5806c946c35f77bf3687f82b5359f7cd3bf21a08443530745aadb1e617768fbae8029f2875ecd67b2322;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd69f177997556d19eee2acef1233ac6299c4c15e3b88f43c15e01bce667b136c2222ab021e60a8fbe933ba2c03;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16c1c1e55bfe67be89a0bf7cd3d9a60308f4b2bc801ae82a70f0ee341f36673ffb30d5a0aaa638183e66d10a7ec;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heba3819e4cc5e8ebb22699bb5105bbdb71e851ca558581427a804e3a42cbd588ba9846a3206295b1ac8629be76;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1091485db7ab2a1980da0681ecc44e53290f12556a6beb9c16ed29fa132be8925375e42ad91ea603afc5fee7fa4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc7ef0b4960d29e14c0eaeb918a47f58c2a4843463d4f301b33bef27a86f37dc0460a58a9cce935095297ba062a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h100a5f3c74ac739ce6cf137a7a26a05f953962ce5a42bd17fa4d2665ac16f6523166a1199cae815c31bfd821cea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1053d8e6f0974fee04d68baa867df551a5e148d79fd8a78877148551988a94d373726c449acbcbd3bfe520d3070;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha5a893f735fc4e84b467fbc63b671041c5dce70d70532735e815cb2cad2da6b5f21c609ba70ba0431a1c24c221;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a46459b184a7e4c4b7d4ccd7372f84208e6419b098475ce53c6376436fccab0214c5519135745a9f20e0fa9c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h541eb3525f0f83b88bd6ba63db7852ca8e4a4d1f07de6f2b5f48a968dde701fa1d9c89b55e8382983cb3c5cceb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h170d64947363417598160f8ada1ef3fee8dfdb9ad25beb82fc9194ba5d7ef4832f30fffaca635652081a438c7ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h124c6b7bfa54550c873c570c48651da2f4d10dcd2acc78c093f5f40f1cffdb4af5636884d20e04efbb30dab5bb9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc2a098f11a161c00cde15b04f3c058499ea948a6f4d09f08ff13f11dc1314253a6c02e25f3824f15c19539850;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e93ef5aee9ae198bd9a2820c7d5b06bb0cecd020699dd628188799b8aa66f37aa96b45d9aa7e0b977813fb4403;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbf4c0638f5df6742d426014d293dc3e6bf4b47dedf23e1ba7e24d27dbdb5c8f72968d9b744b25966b76c18a71e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a145d724712cf9446beb94b17c11be653453db1a831edb20f46e857b3d6c2444f7416e0cab95669a25a5a32a90;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haf62ce10a312c2dacdf58920bfd1b071b40a400e50101cc31034ceac600879dde466922b1dd2ebe4723c13586a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13048bcf22d785b09c1dd3c9334c91d530eded5c5fc96a17163adabfb0fdef92ffcef0b2a3ca1e4e95607c5b69b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11f099e7708a7367e13c32b7f579edec1a3e84d93924103a4c4121e151b924b2de3307f0e1fbd4a407f1057488a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h190bde5103e786a01fd313362efd0e29b03d74dd592746e08bbd71e9cccb879874240416a8c8fdc5f45b9b5cdfc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14ef9f37bea45f2b471394aed57c9c08a9817d6928250f0ae3889b90374cd86e2b5c1c79b4167a90b49613754e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6415e33f3208121c7de39d3e32fe6f8d95b5d46fb4247428604090773bc2d93f96a22676197045a62e2d6b8b37;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d84b21a147e5f35aead389e61066714eded616b7d5bb85ad792dc0fc6cd363da56796de190dff7f5edc149a675;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha7392d1139b2b70c39df2e40d68458be22024d10b4f4674a226e773109aa6090a13410a8145dbb04020045efd7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cfc7e44e1b5445a7c0dc4ffdcaa1990fffa72233c2fee032f01b7b4520c2408a75be208b3dd17c111e5f18f052;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a30e8411e0e46c80e08e0d4f13995d7e21f752a036f86ddc5ed1f7de21284c6c15647751c4998e3c34d432165;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a244d74ad337991ffda898ed5eec957407458cb8f725dbcf63234fda9c4aa39e15e02a5e5a3cf13d14491e19ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h110f290c2cef5e2ee85979b2889e3c80bc4277540d84b3e67f1484212676e043558b88da49aac9eb19743450c62;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a704ea59b7411bd8310f222600fb7cae070517275bf456ddd202ef2307366404d41da932b25994ca47dbdca0fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18afef0c9f048c08ea40050badae8901edbd39ad7686f313f22dfb6387c3d3ca863d70ff97e0c292b158e344d47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15cf968fd01b5c45b7a86dc5948968dfbe7f9ab76d2ec16c9b255881139a8d682cbd3857b5dc77278ea4baec791;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f80810c44670fec11d829de9d7c6a49a27c5db3cac212da271403433546b17dfe97d4170535d7211e5a015916a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hda0d36b7235e5565c90bb5f69c303b656cd697ccbe39bb1b1c2c325775611ccd838f73c6231fac39ddda642581;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1213e15894dc2ba3d6c63166a28069b2056a5b12e386b605c2bd07303a47d7cc09135ab95dad51f6f9b65ad2497;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d64690ab2603b01ae0a4d6d2397148e50e79eac480cd1f1c6924146ffb78e71ea613de34569a9fb8a562c0b61a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h184ca09788dc3955edd92dfa9417635daa42da7827eae4e4e3ae2aca12fd4f17080122593c9b05bd00aab8587f4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10b01364d32ea0938a834cc4eaf5adc9406fc0f34888f6633d6a6ae0a4e1a2e469db38a11ef323e9c54f6745614;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd3cfed0d69eca83c9571f52ab1771d42ebdd83129c2db1562884668c1e8fea77f075274ee164c09c26af460a2b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2b0ec9df6e29edca6319c40e9d7ac8148c234b066f73764871fc80a727f734682fb052879f4b42418c98e13ac;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he53acded167c515c81abe8d086de0720638c4475c01a6e591ff2cde245eb50d3951766829df9807a3b04e6018b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h172e39bddb55aacb81375c41b95d2a557cda89e248ea18bc23f3e8c5d5af772f1c8c50278c8fe43daaa7bc34050;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f66e6b2095b17a033977eed6e3327de0578350ea7ec57923d42825e7d85a60f31de4e55cbd1cf7c3241f5ad9da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h719d7ea9480133f605eae53c19716bd503ee8a0fff4cfbdd0e6f48e78462982b25cf4a70bd414ca8d5238c5b68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h79cffcb0374a013e3cc251a1be1b63ca13890d785c27c6478bc99033412531d735b0c3011e66f67d5596263014;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h55c856b2d12a13e91639dce2b0aa33c5addfecb3956be19062de03c86c099ce2193fe52a6641a3e6d98606274b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h374bc7f7d0cf043da9a80e0ee7607a0cfd771458b27b97bb0e03bc8af3769af90bcfd867dbff7b28d8ba1d9463;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f53668b3ead90df699a49e18719c27f2bf03958f9a4142ffb22d4976a30734a12e0e408c16623f2eca2ffcbeb2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd95c65f774c58733ccc5d039e9bc0c5ce5b21623b7944d996a5bd8408bfe8427079753c325769c6fbb89c6f202;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10d3727651bbb0ae80d542266425a0524f3c43eb2448ba37320ab97070b7a9dfb882e0dd8b74bed06a03ea02643;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1999c7e26bc4c679396550861e862d7d3a9b9accaea92c54fb8ca661ca31b94a598cda8e9f9a79551b2015402fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h138e7da09fe8d78a6c2860460e10772fd2d490872b24e113ded3ca739e85882fafd9eb59e00b52aa77f18a5adaf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f1ea083724b7770a15e3a77a70e5296692681d52c34e058bc25fddf0877246f676994eb90032bf24b52e261e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1228b61275a8a7c18aa937d733c989ed28308fad4ae5d81ec005731c10cb163196e9521de9ac06472b5e518b902;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha8fe09945b592452739e5a31d0586733fde973e9269da3ab6df7da598a8908c8dc7d4ba13a07c88e7e8f93f296;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h984fc33365ece975cfef5286af799334822c586d1c2c934dc28278bfab9c7fcc551c99a6cf6b649c59d969364d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8b42c7c321a23112d99bf23818da220ca56384345d56e0baaed51d4fa79dee5dd5b3bb103c7325a467e702bcb7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec9c93eef9a447c5ad610efb2837eb80a4fedc74e50efca5aeee069469094af5b2bdca5c1853fd71a223d1b7f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hadbd77985e38cfc2c67b84a60978897d38aa0a38fc807ad9b8b1711142d0150b90db3ab41d9d04609bb3519c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h489a9c240d2640f7f7130b11d84e0b282173b7486c76d3c73bd57660cc7c155fea9de6132c7b282b1f40b46486;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5dd54071032b85c22b89783256c9fa01a27352e881ca22d3036818d89cd770c3c394b6671bcee755e1992294dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18cc5e9c56e4454112abd8d33c34d3e7aa065e22bbe3ec9bbf2227d901f40f36e8dd452aa91ab0883a53effcc41;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he31d5692add9345add1d61da1f0b41b57ca47ce6c4be056c68b1518541b7a04534f330d93e910ca86dc51a3ae6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e3327af0be98030eb45e84f4e809865250ef02f6ebfb5b1d375b09ecc120ece867f4cb6b7a4a49565eef1eee0d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h179f2294ce428bd947cf5c4164c8205677a8d2f8ea81bdb94d2f2e3be53ef4dbd7172e350b0d7880b912482c981;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8218489d310248739fe8e98a3a44371743bd9a287df3922841bec901d10f124f7a1e15f214b4b8d339299cd49d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb539db9b479c2f994094b32eba8a395c54f6462184460dd75e91eb10e7ceab4ef8f7fb96f97f3ee4f66e3e6085;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a36b206905ce79e8ad655c856dba7428395cd3a98eaa68765f6c28565d28939ffcad845d1a4d55b9e39cc6d294;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1050520fe15e9e2daabb7b67a6b3b4fcc34c348aea193a9f7242938059aa69df1ae22f41996f2999c0e1f22a4d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h648e666cd7eae5a3283cb56a6885a10aaf575d4a04e3d199de30f520501604d7a056695c66667e8e112651aafe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1af7463a79852316a181ab3793d096f048902eb442e1d610eb01632a1abb759a29ce5b7b1e8af115cfe3c037509;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2edde60db7f5fed1e7772b9814405f2dfb0a3a8148ee32686b810d8ee34e79b8df241276a66a2453a1652aa5db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd97cb91695c0329f15f7bf9a9877dd6e6f78a430d24e377609149d671ced07f2aa83798b87fde804411dd67c1d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb5168c0d0e57fd541419744b12bcd2241fe36111c269379226e91fe4bfea1e8a179cbc848ad0181b257cbc89d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha70cea06ae1ad14916fbe8c4f47f65d5568df6c25c6008f5ccb33766f1cf552d42263fd5d2ac3015d2509c1411;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e20f7150892c05c8b2892f55eeed0fbb4b27e626777f332d0fa12d9110588ceae777c8b74f46bbbf5a93d863a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h132e751e47620e015240a5c07577be76f074216547991b9f55532ccaf84f23f3c72ba7ef4c40d229b0a048aa9dc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1453eee01a06a4fc08dbc9d2f98361306495bbce86f5a1a50fee255f599fec59943a1109229dd5b14d0e3717489;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h114a64e10cb4872142ccf6069e0a0a93ab504f741f06bb322752b82df8ab1aa82a486af67356df6b599b0f3a019;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10d133aff9e9b67e8d7b98c17af0bbabc53fad20f7efddd380471357a3d18b3d6835f3e85223fdfff541d409ac0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6ae0b1e9afd49d2853109bf5b2ae597f797abdebabb16508acdc0fc085d8942b3cb698f65ed1b1dc48d076aaa3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12822a921ea4bd67502c2b9070be4e07819bb15e3d2934eaf3394cc004854ae1f64b785a2e09b36230997106254;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18bc238441a1dfb6a1d5783f8fc13bc6a0e4beaacf414c14e83023a48fa3c94046d3355d866e85cf23b767cae27;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c573f7f00dcf1d456452bdbe9e57090f5b8f4db48a6a83ec9063bbbaae68d5eefcc2a9ed3ad2239ea8924a0285;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h194b533fa88beebb0e7c89beeb1acddba9485ce60a04f85c4e9878de502c28b0c3fafc69d98b560b71ed2a8fa62;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbd6381fee036a1783eafb00d1c89d12f3ab692670dba1d12832562085d4f2a08134c5fc7a48f0a0b3a665a9133;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb1250b0ca9fcdcd3765514ef27a5e0167957641c6b462d671eaf4cc684d68339aef050c7a9fbc635d7203661e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a7fb5d9ee6eb1fbf95ce0cfba7a3273bd48c5855a62fcef000580712a88a46ae7b718484245c61ce6a7ac87e25;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2df9f73472fab2043aa29da2d41b7dcab196770aa183296efac91b7226ddde4f5b32e17542cd20406d1d2f7a8d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11c8bb6460f5947e4d6469b580216dccb05d06b3f8fa5df7df7f7a8971503c5763c0ebe1cea3e7e9a9852e27894;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb1a615586bab4fa6f647d57ff748f804d3956296e5b0431b47cd787a43ce2a17247af59a12e1a71aa5632e9c31;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11daa869c24c16ce1486d18f897317893c2f2413a538ed23a9d0c061b1b1e8e58da637c7b68929cb8c80b28df1a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13f07dca0ffa87dff3cc3d3a67e6ae15a337ac28f6c8328c5bc351253ac8a1c660f4e62f3018ebe511886c6ca64;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8bda50767bb23e3067e73017a9c0769765bdd3a74a4ec336ed03e3f5da9712fd3c2bbbf5f8e4bf5a37d718c52d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha3a1f05d2bd9624744b50e5dfbf1350091abaf30a510edbbebe4961803fa42b036ec9f38dad55fe234b359a74c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h93959989f18e376e1b0e6621e6fb72a8f60e77d59d3da9e87b3dcc0900d13f90558a0ebd216ebf9ae243698ba1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d925ff2b84e183a3ab680054583ec7d67fb1b6fdba2fed177b191090e84899180b978850aa297fd2a4a50f640;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hebae20a3865f509afacac2108afce33d58bf67fcbb69b60e5c54faa227de2499abe09fce48edf4e584f2b887a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4aff748ac20fb15991be71a0b61cefc23a9ddd2d212ab493cfd884a456e2ea7a49dc050fbd336692cedc55e6f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8f7b422c590e113aeef2df68730661ee7aa56f3d3691c24e2f93da84c45e774e18cb506fab6a799c483e32a55e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3c7951f59fecb562127bcdc0db2ed22febde1f820c7bc31f8665b01421bd5982444689e8476ef7c18c590a73a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9c09edf682c9409995ed762e3680d188475938da811e5e2b285b7bd7d5043009f710de4d46dcd2e95a69cf4cfc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc3d7e98a337acb73562765294cce503c941c76ac345f5e8fc7587133849cd9601c8af47157d676d2905434b8e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11de9d70cfe010445027b081c8320e65fabad0d240a1db7ff8fd9cf66a0fcea5426d7779f3dad1eb7bd2ac096df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc030adaf745a7c7794a8b2182dbdb6b5a1482240d100b86b4de019e5c8a5d38601c0248b251c46747e01b27436;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12d4281c336b8200e07a78ea23e16956f1cce2157167b0076208eb66def2da3f37b5770d13257d5f266e480cf82;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a0d22b10c3d2c8f2e4cc282d23f75f4dca0f11f06f2f5cf07cd03aa0394f9764cd5c1d2f1927fb2e6a4f0183e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c28148d5675c6a22218f4749d3bd68280c3b0daa5f0652a6f0c42185aae1ba98e2d56019abebae10b5d8e8d95f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ad69cae0907e0a5767003927f8868440870d326930fa5295ceb34631e41d50a8ad3df8504b9f35a2e8e4a35881;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfedf3cfdac7a92abf77cbe11aeb54d94e0829a6e50adce3f7a4e2b2f5d6fae115e9a96d074e06ab443f6f624b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2231b071af776fe223cc84de5de368034034a8418c2c1ff4266dcb64374e1b8bbd8ff6a42b47088022dfe0ebd1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h763e8cc2dfc6b2dd1247dfc79dff678d60379bf0fd9c5e954eb59c6b8f9499a3d72df732af11409e2e2236d864;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h441ab0f76fa312fa15bad27774378ac61a3d7b6a253a9e86e0a8ad3f19180463ffc0afaa48d5a59b717848e8e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14a88ad5597474e8a79415de3ca206bc8b443e1ea0e47502dfb5ce8ec73aac0b40f60eb81b1481a77cd68c6254;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa3b4814087bd1d0e32daf017c1e1b809f660da0f62e2fc242dc645a6c7d444146be69834d82f903bea6a0ca2b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h23f3507989cdf650aa13dabe32eeabf6945e67a680f285af8175e1079606ac2b49ca249720c0aaf1f8e732164e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf158bf47e19d2d282d92d4c29f58770cd5ff67fc6e8c0fdb45c5613d0a43511a8cd2dc302a4acd214d4be0855b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b936805c8d04057a8a36cc0cd70b2bf0cb460e78a4d88f05f23d6b3e39f148cc245b55f2f24b2015237f51d12;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15bd507b57d56e7b9cd095ca94d5e6de49faf6fa506c2792b85d9b6fd330d8ffa3dc70a0bbf362834d1e2ca5429;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1380dbd87175d3c72a0248199d303f77cb78b25c3de272f45b8cda93ad54bfa806dc038b527fd0702d713c82162;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha7dba76676b7eaac4c97cd807d0daad2fbf731af2561fe89be93aea74eb91d5f00ac59b4b233d4d1d51ac1a45b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h117652e8605a34b2136d6cb389fbcf1c392d2c11d3d05e3c017de5d1b6ab9d240a7aa1b708d64814aae1d04abea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h116100b79d2057272ffc1773b65ddf45db48fe54abf5efde236aa65053904b4a8af03b921fc12ae561d831a9165;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h89932f267a498386f7f97bc4bc12bda53153aafec6aa855eb4448894825c97a8c90607a6cfb14c61b55ab7b36e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13e62f16366ee84df8c78bdece774589769a2cd9389159fe7ca8c50101207cff905e109200d2a096c4c51723c31;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7a44459c71be7acfcdaef36b96de0d82557d859c859427857e01fc7693c636017fb10a0bb9f06f90596e973f7d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19d41598c6bead387d06bca336266e0c213f7e600d91a7e942480227638a8609ba6aab9e9c0f2f3bf96356d28d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15ecadb9726ba4700bbf6dd19626d8e65fec998896201c6ca77e79e7e9b7f25f59d90f1fc6bebc45c732ec9d59f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h102937fdc43221832bb493daa629a882792e60d603c7ccae5c563413eb336426ae0ecaf2ad1d204471080bedca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5868b63d55a30d09c938783d890a3ece04b1675d5516405843b6e0d4093b887b5a3b992e0f1c9ab0d2171eb45;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd41f3d1d9524132d2293e57ba87f29ec1099ac66c18df605232d465deef3ac0bbd9e21a986c6355ded038ab6d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f13f60540ac40612fe7c4f5870afdaf3fcf9982f1766742f33f9ab12026a38a4f7f91786e0630d364f03b6576a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ca1712f8a522fd7772594904234fa53c1cbd4931a76d64316da38b5821f895670ff5c07ebb22aae61317f33ff5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd1126310191f8f12b640192e52101ea5995c43d832c4617a9484a01d543cf00922cd11db7f939498262e7dee28;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a3970aa10a9a6b110c86ac1705c1336b91d3a30862c5bba459eb9bd7086c9e7e1464b4a9a65f21b160c383b2c9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc5c7bb96ed72d9dfee9e30390690bc0e61cc48c6f8bee579cef52847d1b8463f7d44edbdc937954185c5913971;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he713debe27a730053a1a6c38085ab7dbf276919a5548701e39407e1d0c1873f3953b8a05f5f9517ff38b453497;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8df4ee9565f6e0b1288ead016b7834b494d0c56f158c1e60e328434890a42cdb3d1a5a0540813b0c465de859ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h106bd2e3b36a3d198c83d2d7912875b9dff5c8d9275357b7a1d759dd97fb94287f154f5bbcbe0c5ba243aa1e5fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1319b3ea141029533e560053ca616ca7709cc0231ef065e979106ffc34eeae464cd5b74063913c5597cffed9ab4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h890d19448d328c900db43cc74bd5f3ba928255fe3d578eb1faea535685fd02f4106dafee747770ef9e79613acc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd77f89c33c977ddfbf42b4a0c87333bed64fe6883f202016ea401a48f61c128f07cd452f9fef1bcfa282fd12a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h131475f0d054c95d2a2d20fe186daac8c2996606c4ea90881e7da5356ca401ba9634e41aec418f0372b39ffe41;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8a5285378232357d33a1b92c23ff053bcda413eec533d25e8361688d08ac77ad301764d3f93a4d884196e77910;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb50a1307addb4d5465f63615451b90edb843fc9f42f36482de65ef3552a9d4426c9e2ce1fcb7c2fa2fb31ed15d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he34b1b4ca72649d9cd66656c6589f17099b935817036cb8ac4eb5627bcf56f4f042ac52e30dbc3dc2cce803c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hbca787cdc1c378a647ba1baeac54d4bc4f5c7a3be803085f50ed3d82092a419c254fdec49e510cb094d1b4dcda;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he3087c07bc5ad0b415737beb0d9be4efb212d1833aa437846e96ef401d3b00688ebf2062185b64e7d4fcd99929;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d78d1ba0f79ce4db6f1f0930ae000c9a1853e4574f9078377966424beff8eda5dcc835defd727156081c94b1a3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12937a7461a49265a6b993d82a0048129a38f16547b8ab15bdd322ddd19943d6321c7c2341221f4801c2a56b3e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h116b5fa73d288f29625f2fbc2ed5208c752c888fb1a03588fd658a56fc4cc27a6be31cb2db9227ef8948c770ca8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19555daaffe44a26914065d437496f048c0425f03b8298ad560e0f2874c4627936726e2706b391a746b40e22d75;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10eb648e9bd8e27ae2b8d49cb90ad7ab9b7182e0f3de8ece4d4bdb4425c80519480146fc0929af7e99145d7058e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcd60b5dc662b4568aab0c51c7c2f6184d164570417be8615e382913ebb54c34cd41623af31a36b8cff3e1815b4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1362dd4543b01f9c59d00af13159a56c63e95d2cde9bc0ef67454b3d24f7939587da3be216b1d45a02172ba4749;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8ef97bf7648c90d4e910c59afb9d541ff4a553a63b3c922de635002181fd167ac7db86e37100f14eacb814bbf5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a9c6b5641b38ee65ece6beb8dfdaadd13f52209b02e8abdc81c3e75fb67170c92ca7dd04eb6827c627846af5ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10526b5606015df877dc5e0b24bde324a875721aa5325d42c0904be0a3cb89529bdbebdff501a16b6b2278b2997;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f32e79b6bc7bc09ee846f5ff0c6edbe25c18ea0a92aad5f089e61fd671ce9a949f50f0bf1c68e9f675886b5cd0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b4a434327438fd31af5a03c12d58513af152b81dda50a0c8261dc4ee0d8c34c67271dbe85c742791b202377643;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h453064829b5c3f1d53cfd7ccd6f3c4ec37d90a9a84436783f51b80f22ab6ac7d795b5624606612680d9574ee71;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb72ac37977b1d9482d6c1c34a71b5cf2697f0279620c7bab99b2df4b3e0b506b85f5bd45e0c85381aa35edcd1f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d463e5a9b663143d1bd9793f2bb755746140b82de9b62f6f8ff6273388e32ae53a837425c988c1bfd687264166;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1de11c4a7f46afdd630889fec384313bf6cf8cb143d6211cb3ff19f2bcfe80f342d14d4d8044088c27ddd1ed582;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h163b35162ada5641a1cc907999adfae9c35c76f5e0619bf03da12dfa13f60ed2e55ebae513572a087635db25ccf;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h109424d46a52016f1a4b8121a8542c8bd19be009542a105e850b194a6760e168c7ab748fda8a6029ab1ce7d9783;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fd767bd9e8c8df9f157530d45c472c68fb9c31ff571dfbed3b682e58009c627e4586459e49436b428ae790ccb9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5c48a000709966536c6fea1305e0ad3d8e932565789c067c04123dcd2fcdf188292da0e443433f525e47b8b42f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c3fb5376178f5e2f781e1a014316413806e293ffba77331a6d525a6b4713c74ee9e838490ba793482abcf27dd7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8cc4e0240d9cb9104fb11d13c1ff598e54a7d286172821b0dc8384e8142983287c48b61d0481ce6200645d6245;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1332800df4cf1246eb7c9b20ca65ab92de384598ce21b0868178785b067411e516b85c4984119264d0c45f5826;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h137770c1ba30502d19b6752d128a9b1c24d20af615db33f2cab4cb57aeee1934316587bc37e6d2ef3a355115f0d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11e3c847640f360a57fc2881f0fce9a915d4dbc3c645ae126d20dba8510fc439c95dcfe8d826fba4015a80e1e51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3071a95a3679f1e875a7d9a667fffb557994711148ab1ca8ebd8570b6743d811e3710c92a83f52a2068071f7ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e4e14541f827a6970c6d2f73dd9b53dcb045c11eac0a6a429eb96a0d3d0c262c44e57defb22597d36d3eb33a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h59bb9cd95bc1120e6cd5b0b9817335df850510452940dcd2902a58916b12f0941cd7b6242fe0b1ad76b768c672;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h53636fe8288d92b8b8929b56455e160fe02bd6ffc20a7e385445bd114e65a456478619ec85ada24d01fe44069a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h119fcab29e460df631b78eefc6e19784ef87b9399630bfe49ad924560927f1fe1ac1e976da24026c65d91291956;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d676220a98c60f79e4cf6e73498e1cf74d5615ae17086bb0977b3efbd826b4c363ee784ae3ffa80386e4526a05;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5b434cb073fc5e3e5661de384afb7f92839e30cfc186a8c3c7292bc505e172cbfcc24c62e5acac558fbb4b6a61;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h320fc845b37d682494c9f376a2190d228dc1b045f1d567dc654190e5e178caf4a5c9a10b2e6282ead6e10477a4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha5cf9fcfe7e94f942e245bf36b5af5f4edab31d6fd32620ed08711d5087988a4c8406ffc612ea3054904efbfd2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h182b72ebbe005cc8570036e70d2dfbe9505eae58a3012624fcef1e9dd8e349e8ab2803766eade6c9dd8249dd901;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf29284c6081dbb0d3c81e4845040234a8f96c8e9397aff98f494ed446ca02b2834afc47d28ae5c2c57f33e8ad2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12a4cec3e8be7dcffe13a2f51884b4d767d53b74644c94c91ee06e952940e02d304543bb5c483d284b3ae2051e6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b8eef3ff91a069d787dfc89e227b2c17b209772e581026a6c9813150a8e150441a5a9f7092fdb3c784bfb915ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haad65f4af659ffc6322daa6c26d8bd42a604c33a8b6629d6c3bd494d60cd97846c75bef6ef62568beeb7da928a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17b9aab9d6a73182aa08aad45c48e42478ff6beb93bbc90b32a001a2ec8404ba39a582a9ac8c3ddda45b31b46b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1732f4d20293e68c2031432183d1ca70a1a8bfd6d45242832a54380ffa81cf521d1399dd4e8cf239605a656fba3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e9c4c8ef7b6192c1486c54de5b6d6554e024706f130a46fe1da6fccc7efd8fd142f11737c2bdd227e9d4fbbee1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h51eb7610ea6702ed61d02b4f27fed4c1a7a972892b5224f4fec2c913598f61d3cd040db68755d9b9c3d9a013c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14cf32483be6bc3d5779023f72b958643141fad8aaa88f88b09eb895ef7c85e83b346c3c13a0b9df96e93566d76;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18bdfb2882df2d6c5f3855348e7731f634b62bac23f3208832f24e55f35af2a2b620331103b878be857296cc12c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb2c4156dc928b7933ca198e1e72b8b47c3138d4e4f1503f1e6047569309c7a1f98007f719766b934efcf6583b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18e4ec09137cac6eeab25cb09adaa58b3ba5dbecb3106958a00399f7a03b358ae6b1b0f21455be3f5ee4cfee474;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11343eb448ace75779bf14551af6ab554a9d0d4cd9769d05399597c43e9f38d016851cc81a8c6ecfe392422e7d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h62b771d6e07b90a5f6fa59593a229181fcfa3ae1c3a54b629483c3e96b23bf3496a6bcc40a4d1ee43728032247;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ae6b8e99a97186a1ca9d398ece7788d9f648fb99eb7a60c2ad79c75b38f5ebad659c7ac09bcba35af054233179;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17b1218eb7bfa7b3771010e2241f7b9d7d5d311ffcbc210b07667afde507a088ab7bed34ad658628c1381631ecd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f1eb5d9f991ee96a8612e1a547ee2d53bbcc1b4b552d83569711d6fd76d924237d63649b017011ebcddd7fc423;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hba6aa371439c5916c6146cdaea7aefbd8066dfd51f6b9f676d5362222f0657633cda4f34c553a0216e966fea7b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb7530615b6c50e5afdde87e8cff8be2989117f3c26cc764a82cadd4ce7035c77f39e1aa868fbd9a7e939777989;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h227d63b324e01399fc86bde2844784e91fa588fa0b9d140f4c082a1094200144f0f1f96a10da32c641d9d848b5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7b0d056acbeea9500bea75ca3e00afc89076240c116bf18260fbaedb90ddb385117075e3bcacf400774ddf85a8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17db4a5903581bc4dd2da9d2cb89d5e535ea246702a29884c392727879f21607f49d3244e0ff7190c89d8d3ac44;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dada22df2a5db939d301827474f6aa610bdfd1eb1b1ae808504edd878ee6791f3e91457d8a9be58337f619b08a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10ff3aba9b1bb1c5dee595736e0cc5052281581ff3dc8637151cf8bbee2dbff95a2649b1646bea23d6bc0c2de2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd1ec6fb7c67329cac456cd4823b7ffa3c6b5b90cb8190a92066b3ec8a92d0b41aaccd141bd92485f0ad4a4180e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10a7cb4c131e11aa13c75c352c03b66cdfe84a8a343401476427f6bc373bab32542956f9a190466bb0f22017cef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e679f174a34b73c9c64e0a7f4de1b7e6510bdb4a3f6c3808222e2cae7dfd776b4a00c47eaf6bd784d31be87afb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17efbd627d90fa9d05d227ace9586437bc5acc9ba38f9456aeb8413d745959d4a2978f1b094138183ea44d1a2c8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd1b03392bb040275bd8578ff747f46d726b1a6a7ec9e7b95240a0e76bf1a3c9966cf128e100823bcb55c0e4e66;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h187f2140b5b838530d52a8b12d7de94731efe2b42017fe14eea07e41ece0ea48e89082ab72129d438bca8eff9c2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12a617eb2d091be099a1fb6c61c06b289c3bc8d8736f270a1248be9965d8d2817ee09a6f8866c6cc70478024294;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h22156e7acc3c768bd4efb4bd06ecfebb3dd9a6a09baf41bde22ba1580757a6cdea4774018bd6c5c221a892f4e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd5cecff61d3f46e90731e5129fadc22c30498c1ff16abb1c34553a2997a5c742b7d2b3cc65d8a5c3f87c9a06d6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha7f26e5d5c2700a92ec3f2af1e55566387dbfaf1a5aef5ca683628ef90cf6db44ee72549c456511f184d648231;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14beda2ea3ccecd05a131ca9bbde989bdb5f2480908fe13b0a0f6fd1e9991866bb504631f2e65b2352d50d9b63;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1550c4a5af723da33df6e18b9c1a7e98de9a942be184208fe5694129dafb7109c0fed4eb6c77b863f423f27dcdb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1544d7cae745bbf1452dcd6429fb7998f6937833295df3beaeeadb4cfdaac9934a9d900a53f3a78ca0699688643;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a672d3f47ae561db59f9e4b660b074fef58dc70cab726996ba76d59c9ce98451e87301076520ac64a4d30d52aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc920a2a85d36b979689ffd388c73693168f904fedf575746e0452acf3ef35ad05d16b88c502ef88fd5ddf5879e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17cff89f7cd1ba29a80d898d800e13cf642abcd540bcae2fe53aad5697274e5375a1ead8a55225e6405c99b8d04;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1397ac143701cb8446456bf8543e11c52abcc07b603bd9eb2a617e2fe8b71705ce976b3f3f5adb4d1b6fc4aef1c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he053c9971210a25c676eda39edafef4bfe1d06b162c2c3cf3868bd0a81d41abcf5a80d053df0a5ff444f018709;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d32735ee3b6f08c728c5a049cc1b77cf69d9a9f591731cffe40225627b9e11bc1fa3a9e407cd6a33d5680edca0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aba37f41ffa50e44e3034122a509ee5bcda9f9658472dd9a1106d88ab97ac5bd170d30c73bfd84a79cf74d894e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hef06e310382243aefda8a7b06dc52a5bc50be6f43b5656fb85e298b8f46e917ffb12148a4f564de00a7213e94c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7f76a9790430f104d1767a51f9e398700253939bc76a1cd152cd79b71473e0310dd7e1f535fa611e5a7ceadc68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10762d88a3663fcbe0d29854861a8833ec71ccb1e50577d4a8d01c6ba3d51b8a8aa0ec7e1d238eb7d7ffbdb3410;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd492fc4c5799b8c0cc452eef16dfc88b241dbbab2e58b12e59c9d40b0b3d3551f214ba4892d71337716552607c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h159b76e48d5eb3f7039fe3722299c1d2895bfe6c259d72c4012dbc8242bf20564c579a03aca691297b9af469aea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h186df1fd6fcfabb93f686e067a22f31c010804dbfd8505c66819ca72bd49cebb83a6a8e42443bfc3f47080ced89;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hcf953e08333178a1f12982e8152237000275129fe64ef56fc2cd2d4e45b333cc22d8218f230309548185c71286;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ad4fbda89e52b6808b1407bdfaee5442e17bc096b942b3b2afbf9769f0282b7701e58bb6691ae1bdefb82693d2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h165aa0e7155eedd4c507a120a770596dfda6b64883e330b24f3d37948ac31f900cd1c8e7e176d93873f36002ed9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h25c24aec2572d8be78609e410e294a5a530acf4c9b4fe4b4be7ab21b9586860d76df361d676130863b2c71ad23;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h72e68d50ca3d974a6262a420378ae884460c88145a9d9f20efb3e7357c93baa2668ca3a16ca983155499834d7f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c0a97d5f182e93e1f98dda9b75be80128b890f3089e030a13d54fec5695d8118b4ad1738057811dcfac07940b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a966ab7d0bc8cd0bc22f893e46ea28a8205b88d92456ab23b8984eba341a044432512e6b36bad804d84152f8a5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e8adf6b3d3a0c949e252931dac2c40ef9158f10b07c315a040f1ee4e2d1077126c400abfc6904fdc55bb816bf1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h191083a8c75a2c8d21e010bf09187ad28b3b0b85b1ffabed545746086e1592ecd79ac9118fec7902f84a7bad36a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h50e04368c88cb94942f6d5d6062cf62e9dbbcf63c654fde8bd4e6a13885a03c518447c9f35fbd25f7eb2bab3be;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc3268913da45bd17683705aceb31c65f376e821f098e768a369945f1dcfe7d23be299bdd727f1fce4a53f086da;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h70529637805e51d4dcf7774b14f23a21941fb4369016be0bbaffa0ea7b88b6a8654449b1ddfdc60e97f27c56e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16982dde7611cb1705e2a5863cdbdce589781770f98632b546a0926e79ec535160c41523b55df308517f27271e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c12b03a34fbdaabdb1759f1baf963580daa3d3f05d4209b861c121ea06c840ac237eafa4fc77df97b739185223;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f9adf163b4d9443d1910c649b74ef826d97927907002cac3663075da1d4a266a94d19f94b61a6e3639a8a061ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h33c614780ec1deba02c2e5f9a0342f67c08a6d54e074dee8b5ff2f4b9aac684d040b029f06f1c15f02a5bb5016;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ca3c21b924186590216eca824a1c58ab28da2204a87ba7ab32d524803d8fd1e3035996da25484abb92ae0e7078;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hba5a601c901024610ae7cb1e96a3f7efb7a6979cbaec537d722ec406942efb6c0085e419a7345516efe4bf5296;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7c1172ad128c52cc0381594d0a9c6f7e41a32239cab0f76474ca8f6860f7eec9f163a3737a420d791a2f1cd407;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ca9f928598139027e3aa9980a8e08000d42901efee35eb7ca7e47fbcd3cb383a160808af41ed22543c2a61593b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bb117c0d9005b7ff7fbf7ba1c48d55092f778804fdab2decfbb14105800793ab2c7a20a112ddd0749521dcd08f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1686bd5cca4936abe0f4cc3cd9f95ce76576e4497c9e650ae7133c24868e31899cbe3ea7fc2c1979ffcc5224d11;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h173da92a257a9f4f88132a9622daffaa2902e629a6d7da6eedd67e6b6cc0a1f30a3db1602638f889a0d0b9309fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1007ad89b9fbbf015ba269420073bedcbda7741fe26d17215ad9b1c80b482a634709306bbd3e13099ff846a17b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h144e4ea603742136caddcbb5fc3fdc0786b9bbb9256d2036f5f813aa586af4c5d825a0fb87d755134b01ec899cc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bec3c98f8b23a9effb6bf11511f9fef20daed293916de86c82e58f7463c662ec3a549fc0aef2d9a38e8a970804;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1caf9e72a657552bad21b10d040305c0629f8082a6f3596e22bf21663216eb5957cffa1656301bcd87712967995;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf81d2d6f6b8f32b239a34fad03e5f63e955cd49cf0cecfaee3ad8549cfa7d8bec9ed5c349c7d65f456e54285e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13fb759acf9f3d82c94e31d3604616a6670a22067ff81c4d9c83605d6f6cd734e4d5257bc0945a932b27ed378c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h75ed078247b19c6f7b37483f341978d3fe9a60713c4bfb38c45f104d6903a743bb512cfc7584cff917c5975e43;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11dde0f4e37535dd6dd68150781a05a526eb66cc0cfb27ef29bf258c77c155e5d4d5e2ec8f86bdf19f54234662d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5e98bd731f3f9465c88f8a2028b64c85056157f653299d6bcd4bfaa21d2e026d8845ef558d8529f7be28d695f0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he916e497b12057182bf8265a434f024e85672481470ad325925dc5a7cd2e394d717e06707b6f01b426022a9af9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1139ef33a5569b6ddf3500123365145845db2658b246495c378f9074b9a7b3e093332d1c62ebed71c5179da5d7e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12025b9601f538a959675dd1299984327683aeca22e3a7313882c3e20ca3d87eb4da1c5ee6f4e54076fbd246cfe;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a30d8c937cadd9027bfbc33e3c6d60a45eb1316a393f7811f7668a2587fb9e292f47c43fcf1755d7c9db670101;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13706da24ed22a69d5017866fc2b4967c073fa9268f70fbff3a10eb69687e6257d28f9ee3bb10f77ae170883215;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13b5a30835fbf372e1ea1f6497e7f1262a0fe7e8c843c3645f72790795c111c11cc333c031aa775d4879b42143f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h141078a4a70135ae35c49d592a8ce9c388dabf13f7eb92747ccb4568f0163232d105a0a709ab5100fd6e9455b32;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h83b9faaa8b0319672a31292e5ce97e3d20cb130923f71ede6042a14ba7401c2453a32239a8a896fb3d2fe84d85;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h106502aa1b169129cf879a37b156f25c979dc855841f7430087f840488db2c960ec17339a28d0ad6c7bf3ac6239;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f5f35d053489880a796ab6bb4b608de22f2197c78794c46af979fd8cfa5a1b0abc65a4c0420ab3788e127d1229;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11d1ab812416096db7ec790bcf08077b6f31b0aeca6c54f19f79daac890e8bcade7571f4566624bfced7bfd85a6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e9c189b099741a08735e86c21210fc0e0459e1e94f8079bd0fc59f086892cfb97343da696cfd80dfda377cc16d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a10515b41d0d033e482a43d83390115aea794e10f6415c2f52eb0849c78543590b3b52d137c6f58d381c61b560;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7cb41678ed3a359a9ae66101526f4d2475d3ec15353ed3a12c7754e490466f27e8df9c9c6bb5c4d24eb2dc6a1b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13f259b9a30beb0613a5c9777a7b426b22fcd085e046ad86532ff4839adefb823614fbbf869231892783edb0910;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hde9123c627b702959a52c2f3fd901b089a729f3309efedf772fc82f60d693584a75b0b87808d8ace2fe82432ea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7cc26377b961b61e7ce03033a61217fd6be3983aa47928d875593db060a6597d05c12d5e42b4fb0da4083f095d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h67c584de95680a9c238b197a9f3b06b6f66cb58859c3a6d6dc054e0e284788e519694d414ebb46b841d2a605d6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a9c19289d585347ad085231e8e8793e5653e97bd01a31f410c92a800f68cec7e78a036f8d68fdc88424d44848c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19f9465af22e3a7dbeba7e5fb3b511312f3c43bfe89dfae98781c82fae4099b9b68784fc25f9dde5e091bbd8ec1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfb9a690da229e0120c8999a1478eff8e7389506f22333fd0edff188fb14005cea3826db2337d0a8c27da8ceea2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdf1d4514180451cdd51e4918b473745858f8e8159833f04ec930ce0866908ed44f911fab6a382805e2a63bc8e3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4d521bb95b2e0036b29e151a56a46cc9b7d230cea150ad109ec03c6b85d2ce8c6896a3aa8341fbc359a0d43964;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7103fe1b7e8dcc754a543a97330ecd52dd7afdad9c870e5d43e413ab93d04460bddb8f4e60e815237b14ad9932;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haa159f746cbe912dc0e7aef877fc2ac04547d3dbf69b7ae3afa8071e3106226495b36faa7cb91c5b2f461e03fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f74f7a22099de75757bd3553ce42b590ae5a46cbaf0d759ccca24f86533a19d5e8ccc9c0563975999737cc16c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15f0bb2c6d29245fb686f256f710f79b1c0952a17370bb240ae2bac94ca7e4f82d2f9315821e3fe433616c4f91f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b01945b1b00f4703014ff0473850b90e460d5c4c2417aa17f27cd11f41e8b4a088453a74dbfb79c32507357570;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b21968d2ace2414b29d47be3e9e3da420a230cef164c74edae0299e9c9a5b1d3499be96cbef3a02c887b9d2604;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h114435da4aa26416695a9b5a2f6836ec906878ff92d7137e53e4c7aa2bbced7f9c47351e220d187f03e350e4604;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb14d294ec1da9c7f7e0f3c163013752bd2a364dacef3a6af30a6d0d45e2241497f00e26e2fb10f66a54e2847c4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc93509443c46205975c10a5cb3f3313d4eb387fd208493bcb72dcf04f2752a0e366468dcc3d74bfe9aa5e23269;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'heb68ffb48e94469f4b3ed8955086d845b67ee809aeb43a4fa41d6a03e95d900a60586ee22826324e8cde61034c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h186a0f751bba8101727633c07ca430c2e9f89f2c3dfd9327470146173999100b09fc6f9a70376298361df3ae6a0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h997dcb1914873a3dbbe6e1a891d40cefa3f63365c2e3f6fbfaef15dd0a128c4bea007b1e81af9dcb23c422b805;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he8bddd844b2e94fca92ef8a2b577cd3ee16e7aebc152b6021b3c7305a989d633f13abace08ce1fae8711b8e79d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h490f4fbcb4dbd714fbbd344dbd05cf20a275c46fb70c1cd2373b85db757c7becc4a20e673a3ef250111f14a5bd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12e8f3258d2b9867b3e4a20655fc9ea451efbda831c2ee3a702d8ffb0be3c726e5e2058fdb1673bc70f92050411;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d0503c20c70d21d61dde177db3d83e1f76f75eef0f5cc7749af6432b88c9360333ec02f0b216f9a12dd6989e31;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd3c1247a7dbf58742e6211eda2c45c6de8edeb4b829a5d44b029bcbd763c3d3070f53fec5ab5744fdb2416777b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12fdaa546147f85aad3422e66d5704f3cc720b6eee75d57794377d39a254fbacc7fb276c3a363181a845e6c5f79;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'he725bff9d0fe72f22a4eeafdcea483d55c78cc41e40dbf4a80329854377165d508ad431fd9bfefa6203c1c5b0e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h61f0010ec6ed8759d5f268280d6ea64556fff61e94abf8baf3b641583ea5cec83885fad92cc79caa92d3c1f952;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13f5e5c277eed95a33181224f9412acd46185dbbdbb583c93c1a5234b6c0fafc08f333c4525a77b2b4e9ef149bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9dbc1403f7a84936070a7a4b7e66469c1635d57e4f872dcd74a404474fa5f598be3e655ebd1a487264b4406195;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb65e54edad438a657c2e0a78457d235e813fd18e334b9f9957c09c006ca2a860e91373fa95c9243154a71cdaf8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1db2b0ca2d646e169e2252ab863dc01da8af3da264983ff9a1db9305c1c786ef4900041e0685fe7ccb239700cd4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h199622b0f404ae0f835b8f0d24c33bf60484000e21d6eee4a68729142330d3e033ed7a9dceae693f0a2a06e2ec9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b071cfc6d4a67221bbb1094446c3479caaaee70503d69246fbe3585adf12158e3c97bef472c470a15632b12415;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1122d003114f14e7e5ee53a6f695dd4d3b1a704948a174c21def62032e382c0f5f70ea0032810772128e502491b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fe35864c0ff3f9a32b071f8523daf4d5e72434997b1116a8ba69b30553fafdcf58b9983b4b50b9895b3f25889a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d7c6f3692a1c8e2055dc2625f06c2df05b1687509124168b1f99bed7afd29a8aa7be9448f5ab40f67ff22b73b1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b9539ac03d64adf2da7250cd6d2b82c486e1470fd2923563033556440753e5ad0db8fb779116ef1a8840fa712e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1414959ac547887af95943ff625f9e94cf5a6c442882ae3c7a40dd68e620dfb79ae5bd9641a8c9254ba76989a2a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf055945367b9f729027f7bae12fa3c0f88e989a3d0d3815824707374a68a18fe05d9294244d421896abe1d7af2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc541878c6b87b44b2de6d4141dade8767585a4bf030d4a5ebd79d6ff95ac2b58cce55aafe68d757e75e04678db;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5a4d2cc75579dab5b664cf648df9881ca437e12819ba7a31e90fc9651922dafc7351615c9bd935172f6aec8fbd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h191b6c822a6b9d72ea6c603c003fe85b04f4579fa7c663e9a51a36a494e8f29e3c2a668d978e4e58c5f3d7431e9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf7992e3fbb42bcaa578cb37f21bee40ddd759174f6cb2ec5a91313e37a9035a79b27b959dc666edc561449bb3d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9a375d7f6719303e2e0f7dbd38ad9eeff7310dc5e3e736759f6ef6f792d3426060b5e9dec7e5e2aec3be11f92e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9192fb8438c63991d1e418cde886b387b360294f2c52246dcab03602fc0f643b6963a8f5e5dfb010137ac77440;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ba02664128ecdabf3b5a12aeb3468c5f0625548a194a534e7eeb3dffc27cbc3553a803864afc1d3c4deeed8029;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h256dd5b9ea6c360debef3287f401b9e100008d5270a87b709607e188ab47078f40f315be60686bff43fb54c4e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h132eebe89ffee143225f725cfe3394b5fccc88892fb0de4184013d718bce9ae8650048da62eb50d7d9ca2e528dd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdf649083cfe8ebbc2d24b389d070e46dc92f45123fa0df05e0a806b47aa23fe79e033c220ce6e552cca4de512d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6a61406fc1eb9cce8e53ee2322310d87c673f0809e0b02e0459c1dfd3d07d325dee8767042aaaac5aeae545fea;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfe554eecc5c44a96a9dcac5afedd655872e7acba4773a414b50e12adc28d8c88e694c4de0f6d53755d56e7cad6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hccccef2cb85d803ee83db8602abf214d2214dbf8ef021eb378d252ebc9312baf9d68a441a20b5e03fbd1343bbd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd980efb90a112c769a9334d4b842cd9760a05d1fbec6683645f7507aed1d07b3a43c9aa172e2704323d642c13c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha66946ec3a173e982898fc325c268ba0ea0b52a4ae07d6a00b063e0c19e49c71ebeea8aaac8e238e7f32b03a9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10cb132953d1281009105d2dbbe1a55c9bba3f78f0d1f9be03e1c962c8f84e018b5229097e654b676425447bb9d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc6b0f66ddf24ca919b17b0724f352576da9136a39946a191257bb22b03ae19c4216283f9f3c431a2da284c5d37;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h189baac59f8484cad65c541b04d34fdc0ce7c5b8a5a2737518b78ea9ec36876e762c21d0f836b835409ef5fd4f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd2d35d089df00d1b884444580a75b18fdd055c9a28dbac9acee085dd25b9d6b0c35bba88c194c27c1da5ec7542;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17e1c5fe2cc00f23547485878a5b823cd1a6e39d80974144007b9f7310beea3d3700a486b981ac1c4162bdbcb6e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14a02d23fb5bfefd6c420a1d59a636d9830ceb2fe0a7c095335cc96d750fc1736f69a147a08f8a4ab40ac4f7b33;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h133892b8e949a028c09db5f1bb7913fa1b645c00d8a10020cb5de5bb228bca30433550acfadbeb3c444a660dea2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h144a8fd3ec54f8cb9e6db55f74dd74c030ff583e496904d081171c27d29a5219ae43548f6bd931574dc7d44ea54;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h315774d8d00844f94fbc9e1920a9cde4f3e4eab80ed369c041b3599f66f040f37d905b0e9463ddf798eb586cd4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8fd7c22c2ff933dbbffb0b74c8b16de3ada2ea93755f2056a0cb7c908a0f56f5d6201f4eca4aceea59d14d30ab;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17a25ec5720b1f0e990ab93cd419a1a827ea868c4cdda463b639d8a3a6f12222727dd0cfb7720900069bafb1cf1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12499dc4f324fceae0f701a3a5bd7b9ceeffd4a8f6ac1e1ad8eb88a45a5a4500d577cd4426b3e4ecdae9fd411c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h117ae625eb40eeb243c33fd2e14e683db26fd9137db347b149d67f2c2ee2feee60f35b58ef1298bf3157362a361;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc66f046b55b2348bdc6d626fc30589d3d03c3a526b61ff66e90541bd7454e75f857a07165dcf341a36e34dac0f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ea9a7a841670a1b2ff9c7564f1cffa2b94e716d2c2eaa4c48402048ba9781e77b1f8b1efaf813b7fef07ded997;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h108597f0820f96fca1124b873cdbdc80e03e4b1e157d051a4a11a4ac48990757184073fefc028690c4eed2409f1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb1bff608baa06cb47a6e8bd000a71a2aba5de1ce2cfd5d1e079a86dde00a2aaab8b7871098c60fa674e8b5588;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12c1867e5cec7e97c0bacc436a409cd1c43e29bb2de64a4b82367e12e48aca4eb6411f948db02ad2b88ca37c051;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb5df71ab71391c4114974b99e86d48f10cb956d334615f3d3269b1456cc4a9e3ea1cf4a07050cee8968dba8945;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha95aef8bdd793dcb920e452c360bf5fe148e02e66a5bba50bed76ab0d537013c7f09043589810a5690ca7a8879;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4c8f9d115827719886e70a88ea7ccb4b7cbc75d7599493615f6b8c132e269bdb0c3a7aa91a74bb69562f299f58;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdbd201b3e7ebbc347824ed269e33267674e58235b73790a57e6a0b22ed576b7d68ae13b2a726a293074c600eae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h141ad83f99f71fa7ef3d85691d8bc6a387f71c3e92b50c7da12761c1b88e6ee4a4795dca903d43c8f6cd6625a45;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h112c4f97a7042a91ff9b18d2f262d47c7539ef3573ab8d01a7e9e16292f2929fa998c4e9dbe8967567f75fed5b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a73316f0f453ca576161d6881e45338fc7af7a682e5d0d52442134652c9778aa02d50ff5477f7713a41fa8c11b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hfc1eab05e87aa7dacef29ff14f20ad31a07d6447df295b5c194d8debe57ffcca428e1b2d2cdf2e683b2e62193d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16a13299d9a3d9b987cd56560fbda8a2c3ca8c61664d35b97c656e633177c87aae03a0dacda44396c917198befa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf29d5aa911d883d069b6b9659aa67c00df5bdc2f054cbdfa9f8a985ab8040a12e541a31602ce7d6644f8a1d36;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cf61ac32cc620b0b41bf5b290eb5be97cc2729303b8f4c030fba571797de11010957a293c5662248975577f310;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a07dc74603c21ae6d04bfad63b1aa544c2e1faa1849a3211d8fc6549c5d31f1f4b2207c99bb80b5f2972e4a9ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12cc36f4cdc166df1989c194fec1bb710d191c3ebc4b4c781e5415f0385cc3fd95b26bca1714565fc7f3d835d1c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f884625de5a512b7000fda1009ee40e72b91db161014b640ef432037253f3197b5df949c38355017f42aada2d4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d463421e52a75c3609bcdeece9b8f370e777201dfff9739a18be3cb6db69ccd84d63f7666c0fce620906a48024;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hefd1ef791f8bcc9717572c8682440a2d3c8ed26e8362c7de2ac60cb77b2b119976b03450827a3783694757cba1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1252340ab0182a99415175ab5f32939436acd3e24aa2c6ac2e7fb37fe0392e898d02ee2bb9a62e43224fc3f39fa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd430c1e3aa18eb3e1c9a9a29d3b1b0e82eb5ddf40d92407d30d73189e5784e5554bae112adadbe0cb942b5c073;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eef2a095cc855980d7af791c6bb9d7c2aaa8f6d0b5fd5351d945d1274e78118e27a53bf285041d53cd9000075a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h150d4949297b4c54447c9796d310a4a61ec1010e77320c0b3e4dc8ab4c721493d92dfc3bad7dc86f6dbaff67120;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h110c52457ce4b1cb02e54ac4dab649588391dcd739dc7fc46ef015c24ff1b2e11d011ef007f765616b48ba385aa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2f88fcf10a028b24db8e9f72122a74179a7921fa679edee3f20db8a06d4b41986914d519ddd32b34053ae0f684;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1348411809025e77ebf36dc058b08cd191bc1cc7a1dbc403b64110af650e28379297b2c85ae79f7c8ed927e77bc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'had2950e3e8be1f89a1765a756aeb24b3d3730d927ee55a908f8d0e9ea3d7b0b79cff6479f3b4c90b2b247ab41d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ee8b99208b490272fe5a5dd4354e1836bdc85397e2cb2de647406c084428b4d49ccf4359d94b58be15a4e0bc72;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c459fcfcac26f47fbe798c56b7c1c761432b2aac5efd1ee88ea72c2406d6c3af43e9ff4269d2e6c6303ee8c4f8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bd96d259942355707c0e60841077dbcc90e1501a22a7833fa6230166488b7dbdb118ab9872f2ccbe0b5140e926;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11fecccd4b1e95b24cedfa797cc09d395127efe7aee9697c237a485bebcd3f66795f22ba348f6ea11ded2d8dcf2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b30491c079cb9d5e59b6da0c8da0bc0cf07713b6dcc620993cf3c3830f60b97e1f114577c51bfc8cb12a1d63fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fa73b8f46f54d4a22558ab9441556549f290efc121cd6713887b763cfbb0cba08e1d4f18b7e3628996cefa1fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19a33d94d74cb83fe4ffe2134400068271a5e772ad5385eb34d190554ef7271ecbaa5ff975c309197fe021c4d23;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffedec3dde6ea3f855bb77c1f6bed9e4a010a096cbc8f6d322b1f9535bb42ef22612cdc9de993167fcdf9e03e0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4bbd8ad018589ad00dca6aa586a60a899b763ddc0dc5d4b1dc7b5e6f344320e3435057caff9734085c00ccd95b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h534844386e082261a96abee457c00f8cac9ba0d754879a77909d3ec220f3728096493ab514397e12b5cc97acee;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb72bc86f8e84f894c42ab0ab24dc7107f80d5952e8bd7518dae0180b2e40e8a2b37f5c1abfca5c13d0ca87281f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15119b5fa214b928812c8b763b758bc0b0c785f4ef5e9ef5886fd6873c6e38a8075125adcea2ae6d23a2eb15f29;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18a688ba15a692be27be086b60817c319dcd7a4864004b8a67e693ecd2986e3790ef09987a7d1d54c697a2fed62;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ffe77b6c21eab973bccf98c79c67321b73a48c368025d61e7dc367a3218a344870ad416c5eaada2c445410b6c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f8b8a0dd86b7bd93df6d74f4008310c7a1143de4d9c24e93c9217687c39e88df396b329afa0c0157ed3119206e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11f907abc86e4dfef73f2ba08cc6e6385e1e1c1cbbd8d96e334a45cf1b6fa344506eb30a354e3cb7047e7646867;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h112bdde66798c8636823850edfe40f10b5f3e4e10aafc9e4a5f5e5596b986bf814b4cc79410f620b1de60f1bc21;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h88a1d6707923481f6fbacfe7a0508d0b7baa16b5fca7609bb4c43983c9225f2d48005509a2cd0d8f9c3ca48408;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb8d0d0a61cc746bb503eb4b3a2d22cfbaa478d36943bbe33807ed7b3ccf1aa95267319ce1115c6f7f9edab341;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haf16d114eb65cdd91cb61fa71d9ed6da73986823c3d9521edac87299c98ffade2347e64753ebb7e7ad0166d587;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c2d0d6a33f4e5ca11d600ca28c9e60c399b1c73887b937c827e4230095865d24d825949329305870e1d161064a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hed21659363318da67b728dc5912f65539c2da0ab6c720cf14698ecdc17cef8d60b7b324f07545f8b549939263e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f05c92c7ba8525f3079fb28cafc71bde4e5a52671a3ef7e1dad94ed132d83e16dc3db837fae80b7768a114b6b0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haee9972fb1d312712f583001e2d6d05a9c4528c7975fd17df7a3d46127c1e090bade4cfcf086e25ded8999e752;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9aa8ee7000427b5e1b9f2d5f18cc89f7ec5dc5aa626993949b77889e8d64c4869c4279745313f089dc4c20751c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h166fffbd87523708179455551e9d6485df22815e2c24cc9099a1741d804a8b862688b3079953a87adb3f9456671;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h182bd7a5d789a1f82bf8a2675965fe8ea0ecc99569fa01f24777eef9e5278d803346daed71e548b1c4898f547a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2a787b714ec2e55d17236c6c901df16382090e2892fbe62ccf7ff9cb7f6df1061df69b6e47919d98e86a5154d9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdda22bbe8ea84517aac545554f5db5669dcd84bf11a19357fea3e0dde5d0d09bf8360ae45ff720e199aeeb54fd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fdccf33180846399cd2ea1684e8fca42b559e738ad51d202d98648b9444c25b2788d4fd2d17796d1780cd328d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1730d1ecdf269fd23adb2c070c563cb0e02f56543f8210c4454c03879fc7c249e3de3f982bceb5beac02c2ca54;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h106ed51f5dac35838a97379aba90f40eef8b9b54f0e2503ccbfda23f50ca578cd50ea9ef06e0c1d53e0faaa68a0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h197a6a127175582c0b06bbaaf51761067cd89a54646d369d209ac6bfa363e023e0f272ccdae6996addda99082fb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h865d3309bbc56589f15b492d3a9647767d1c68ae0048060ec237de27d2844dd2f08cb19f22d59fd433b9e91751;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6d7171eba60c141045800b10cce0cd26a47080568988940018eac2336bbd9126a95d889b73b1d8e78a8ba6f45;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9dcc5a837be3e21c97e4c89b9462082ed5e9b0d043d3daf4335600dae2382e5f5b238f983e414b6ae4ea8c4ac8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6f242fb65f7c42b35f8541f149772abede6caf7ee07f04f7dab3ee3f59834816c5aa048c29cd0f5532dcd33dd5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h79c8c26dedf58b3776e355184bbf392f2819635b8f14f1fc71fac140b4fb40a6c184f370101f527e79a9c784e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c518bbae3b011363989d9d243f5843ea1931b4e78b45f054757d939e517a8060043eb16198a497ee6d75d7579;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4b3a821881ec21bb1b24cb921842fbaff9f55fe06facb9b4662ac8c6ed1681ed935b35a733f4a47af1ecf06c5b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1eef4b294846febaf080e857a0ff5cd18fb0a5b126ca2f37f8894f634438a5e62905e713ee67446b0bd21486448;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ffdd3ce20755adbe565358d4fb6543c3d7b9224f2e4b1713794618bc77ec3ee1844d021df798a505f4898df2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h14de97bf8d2cd510f30972bc7b49f6ed1728efc8961e54ecad50c052bfd4c3fa948caf096916af2c0d64e158584;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h383c4470a7aff507ce0356f9e576eb45a4eaa8bc6e66b4f149c027f590b806287b67e25d14703cb1567ea0e969;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h142aa27a344e2f326c35b54d76c43cd60397a0465235bec07493f74782faaaf872024782c6235d4d8a75f9149b9;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1dc06de305c9b2abba1e9f48dc563d6ef531bd73e475705cc122bd45f4fe05d3fd6b3736feac7c268368e1d47d7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h533835f7520f7d32cea6b0991702ad1318b48e2a951a0a815c17018d2894f3075591c67cf6d9b9eb4650e4d840;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1acc1287dfd1c9951a33c0cd40a679539d21ff38caa30a7c44c2d7eab30ed44e9f60f5af38daac505027eee1b82;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1820b4a6e5167be4a014a9ed16d8708303a76b3c446cc94da7e6e9ad378506f38a266c231f4f0f0390affbf0872;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h266ed9a1e20df66a25ffb2b92008cee7e64049bb0887daeea621d84cf2f2c85c63396ca3b0d971fc8f87fee0d5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h19b13d503b61a12946b300609564ae45e438c2bc7c9c9b6e9b05f44df39df93df037ad49459f9a37d6c60eb753;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h315b23f46a2f5d6c0aeb24f2abdf2aafbfc56c08685ce25e1904d37941e10ccd7a48b251a5c0c448e72c8f8eb5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c4e059baf44fad46fe2d845d67eca8652437912a6e8329d8207a89b6ce953c65f698ae40b05e399b5a885d516d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18eeb06a7dacaf9914ec2e0ceb74e374603850e573b85f7cb9f4b9f3556dc257a468b251fc97509280e4aa3abd1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h34bc24a6f3f46e16ae21a63eb2c56e5f1a75cba58519fd80e06237f07404326a8b1e800497bba403c0f5b6a366;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e57616dd76bb5d8e59b2dd3715b413eebcbc38e78bd12a331040fe1067ef51574e08c1d6f3ad0aa6810afe8471;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hde937fb2c161a77d3cc22b8e5389c636272be24de266aae6718db6e5ce8fe1fbb530ae41a1ba2c2ced0eb9203b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb3c57b738c5ef6b13c9cf2a6cfdcf6963130690c5366c84f29f4b30f3a9647f281a283f7b623cfd450964e7acd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h626b6cc18bccb23ce2292cae8a50c5a569933ba7b06678bd3b7339b9e64640b9093d3a674426ede7885bafb8ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ba28727b87a50ceeb15711ff3f5fa1da9d669c09e3f10b49126ebef5b53ef7ad9139357b8426fbb58c0a346d96;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1fc15160e4d694175aaa4c5f4a93ac9e49c0d346116a9cf850727c7ff7376f304b93aabb2eaf3efd83812eda538;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h175f0e979526141a6d51796e1ff1d9f61b926d5b518365830b7c95d40a617f905dc545e563b05b0066470b881f2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6de6ee34cf14caa062fe6279589e2ddf542ca043abb73e04f1989ca4ee39389f202ae58bf8ba1667c2dbb6eb91;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15c6dc382552e0d611e98da92b96ca55fa92fb67d57bdf2ff6aa9ba9c1c6dfab61cbc7801a0554035eb11fa4535;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2d80e7c883be6ed183d54cdaa493f950cfbb138617c4f0a57db6e369d7337273c948a7b62e0c4b0612e77630ff;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd411e1cd951e819b4ee3e41d4e26202248ff2d47d0ec461002354956ce90cf527508e27d9952b6168f93c4cecd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h112ea69980653b4be279686a60dec0a508c5d10f1d62733fa2bafd1e7fc079f4732490fcbcdefd0be43950bcdbb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f03a32cc018f8885faf4b1a0111a4171c38c1278056d95d8bcb04ff488b826d360eb6a6d8ea47bf34679d6432e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hdb2a389dba6384365ed4817a3db8c7371cb2dc5823736779960af12b9b4d7cc50117434f9218d037a72d577512;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ddc3e66e5cb3e20adafbe27f1be1b3a9ab23804628b1d83d29fbf380b016ea1c19a8cf1bd14f7c59e45e5cd5c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h117beb86cf1b2a0da211437ad6f3c0cd560e6035d7a774eaabc845a19346c3953986e30a61d116d6ae4fbd3a02a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c0613a8677a6e62c3eb078f52d74b700e2a819c43df7bdd413bad277cca5831ce847f35292cff8ea25a21631e4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cc81152c516bf7386c2902d7202338552f45c6540bc62842ec0c205d0cfd265eb8dbdd788a80d4102a79ca789d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1b264eddb8f381af27d3dfdc5673637b25630ff98b0ba73e52056f65272ef9a3332c0ebfb1a7c5517a062fa70ba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c91341764d7687e08f169799b08fcd2a385ead7c13949ac309a7df23f121f9482004e5118d16151d777745335c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h47f5c1704d3b78595bd6c068098016e60e9b90d36348dc749a179e1a822211ceba736c7712745b8433fc3bff4c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h29eecaff666bb91fc20fb2d83e1763360d2577ed4bb585275b5ba655cd4032c99366704dcec935804a70ed2fba;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf7e1b850261c77d3f2ce2d4856100994c4ed31ba2ca84751ecb15ee36706d71f33778722ba282f8d1ba499a889;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2ed226f7b1342e4beff740c0d53bc67b6cc5b91bd005d2fb23e6972b7d97100f2845afc9d7d0d84b3b9cd267c1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d2408d7e726f64dee11210bbcc61d1a853d394000109627a40a053f3cd01ce5830b434e6edc6cdc4433b9b9e8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h94e189317d5e2845b7aae63f7cae95c3be4391f05987f7ca2586bca969448afb5d64d7c3032d265b2f45ee87e2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3076ac7c8882c49a1fd8e4da3351a49688a49c088a3a244c7fb4985ebc03a220b5249b6dac6e9391b8a36eb50e;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h197e2fe3ee6cdf61174c4d84e6b0fda9ad67416d421131acff38be276ec8c60e4562b2981e10ec1c1d1467c4475;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1868ff46deba6c9eeff3c64d072b7e2c0fc6614ee26bd34b60dd7d9ab92a263efc2bb28b26d9a3480641d4593c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h93a3191a89a95b2015a47ebe48ad1322c640c12a08dd420313ce7460ed1121709b831b048ff1aa651582234de;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h444ac37fdead070b6e0d7b318dd4b17c68b1d4f343ac3393da1b719d681209c50c17183d0c7cd53ec1961b83c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d9f5dacbe0934c5123d4517666c2b22d4dce0b4809424f0dd876fbd27627eab44eb9ef5fbe83823f81659d1738;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h503a1fb73b4fd367c35c2736d7d5decb98b238fa8f311630b74f91c0cc7712f27c551681733f0a32fd4b2e6965;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haa2eecf321a303d6037f1cb3d0c0a508686184e72ad79dcb37bc7e4f9526938b6a8068beff0ae767d1901b79ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12c6a4a13ac7979bbda76b7414d7715f81843d2edaa243bfccd3054c290f2fddeb37fd797c89558f38ce6263c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h25deafbc6a8f613260626ac773e3d75a311841d3f8c734d2f4dabfcc9ba4a91d0944bd3f438a4fa98fb3c06f38;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h160e755a22c0cb85034b410487bbd5060837dad7025a9c13d42a738ab25b6458bc8c64fc079e317f2ddba90c01b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h116c39d6429ecde78b53648b1d36495ec75f61a46da92ccc6f00174e37d8369254928ca42ebac1d912a540ea423;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h9645033e03497228c27a32fe551932c25b8f0593442ade7a0c3a0e5f62251ce208f14d910a0b888c1d2654415d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a8424cab2d1e754f4cdb1c8e9bf20078779a6ade84fda397d4dcc12fdcbf733e07c449fe41e5c154e7406d40ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h185a97e374243414d267d19ec96d7f80c2a6a72bbe03c16bf83bb8de3c31c0f04ab075b4090b9bb28ed6180c83c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13c8c71344707314aec04578312f659f4b6209870276ad3f9f2342db44024e7db7614cbc76c8024265cad193db6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hf645406bf3ba3f37eb0ece11c270b5b368bdad005191dbc221779ac966f49be7bd6b9aba19980f4d58510a9f59;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h545185d891ef9645b5e7311ad6bba3a553ef4d2764aada8713a8def7de4fb214d408bc979f58535dc60daca0a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12384046d07d07024d63c370b2dac9fa5f98b8fa53e1741346f365032ad4491119af67b795356a423c6fb7f51d3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec477119501fa4d9619ea517b2c28a31cd8eb582cf3c6ee734702c9fb497248b654a04d45e77ff636b5488acde;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d061a067ca1d7f6f4b87c93a17e31eefa8d951fb54f505a32f83cc6d245986f66580fc1659ebd20d43e7f64ed4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13a78d68a775cc9aca891ebbcedeffcd1f3ad007944fbb884fbbe62a443d8fd7e936b523103d458ca864538eb5a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c2d93e487788a54f865f024ddc4187c440f0603bb01d5cbc40ea43c370163af13676a7e494995dc6f3b64d27;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h71e5f9c9c6c69e7bd0d39ca2871306ee78c67b11a94da390d69d05cb1321cfadc1e256c77b86a88b0cacc70038;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc440f677a184fa992d010d1a403bdbe25044c3e815cac31ba9d39f66aa38dae2a91646ce314fad2eaf4d959db3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3db6a193cd48cedcfd5cbc0d07635816bbeb2b887ae17c1c2953aac49c8fe2f5c760616104753a22a156518a01;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3b4b8b843718bf677c37d8a128706fd0a1f073b660c65f5483b73c0ab7afe5a202f9480a5763d300f14b7591ef;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h71dbfd6b795d21e5f2afd1e27e26c964d2d4ccbb6c7736895b1be551250873c7cf2155187627ce7819e0ab1ada;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h311b98b8874120c789ab7c0d473c1fb7b4ba0a54f6470aa3354f3627c2b7ce8f97acd66023ca3ced71df96269b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h86707c58fd4c04813f0548e780ae671471bd050f0cd9383f5dbc31e9fc9369044f6f63e10a1ae0c1e92f23ace5;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17333d791cf100c0ac42a669099b1bb307a1accc9572d7922715bc86e235ea938ad15296b95711e17aae78a2fdd;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cc0496d78c2e383d458b6aad7f7e1476e0cc8263db66c816525037b272ccb927510b1504f0cb5bda5535401a2b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1de87743414d7055a6fbd4250513fa3ff949bce42b1e88ff152d64cdeb8bcd51636708f7f88eaf1c601db40ca7d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h69e113c742e8fecf7b30468a600c495a3ff85d82206c1a2ea74b2eb442dcf1186a5494a5cafeccfd2cf04bbb2f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11157fe26edc3df1501ed70a7c458842c500565e0f2638deb3666f0e57347e22a7c220d3fe7db8b7d15d8bd9080;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1daa5c3d91a34b71042b9ad380d2076f6238283cda265ec05d056174986109a76a96ee0b9f3f8977579934ed5b7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1787501170f8de9e27be435f72e77700d344ec866a96ca9c6d80714b94a8b4ec9a9088794d55cc438864216a242;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ec223c4bbf48a8e2e5c0a7a6a91bfd9a4efb6128c3cd0ff4d0cd04c057da2bee5c6889ab06240d723957013e68;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h716c096739f329bd6f87d7b65b1bee8138db036388d9984c9ce9752af24b4efab0d25bd9b728f1ee641fbfa6c7;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h102b1c7a4de63eff32fe8c553e92282b5966cd760d90e44b47757f3d1a6b153b609b38048d0a0fe4775efe676c3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6c42f24d0cc9931d70bf959b47b79c2cff3ff93a23615d1788b61d1a8712bbeb715d77324906b3d6ba1cc8fde8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h60603b774e3b4cedeb23333efcd5918fb9227dc718c38d6e4caec8e2b915ed3c0d8ebd0b14ad1d60cd729a3548;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1bb222af8586b6d86150b4a16eae68d15cf1085d251f43ab96e62cb053d75f151f816b67a89528b97cad02d8ea1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h8237e720b9398dbc8cd65f901d9b9ac49d46e28ce122127485c8143906efe2ba43f4ae1814ba8010b4994d0b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1af895608f91ace442bd52debef91858fd28e5a14d41654c75721f9c0f12fdd93f7c9af7a6ad92f821a0b6a7d35;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18e4f06c3c2a48345ca429a42d986f7a308f0dc87d9aa84fdf335428799d9ee4cace644899b470ca5c0e1a65f41;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb33cf6c019772548ea440b637994dd9fc1eb9dedf878a49b6d6dd1a9a6faf7379f3666bfbfefbde4927d433523;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hff33b7c1b5dc3d5744d1cc12e9c0972a5c995d7749db9b8483d510e6b9c7e6f683e7a326c6a054b1d8172b2d58;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cb96d75a2f67a11266ca389914df82ce4370e03e1b4dfc20330d420f01a386e8441428b4e58b184ec6f5e54438;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h6c1cf38fefc60924e64d02b1505266dec038e060298ca5122b74d44d4e295b9ecb13793c26dffbd31affc1f7b3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h520e214eeca2645e0974b83e8979ccc0f4c3eff63162104955e1bf57309c377439ee23e1da5f532228d122f4d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17900ce1a03c41be245a4522d5d3e110c1886b214b30e8d2db275102e6c0e2de9a90e59fe0d04279ed2a3d78f04;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h12652794bbaef6c2703522a0b1e9abdd40c335728dbdd3165bc16fc74c54e009909928ca119d8648f3fd53d9bc4;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h146b54e6c4cbe63343bec0c2d0c06cd0695ac2b27818124f3aa11231dc0b9ee1f2d47e708e34cc533daab2eeb14;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ba5d17849d24079db1974847bf3bc76e4e4dcd17cb1391f05b12a388332e808e52b9d1dc1e3eb10778f2f1e9ae;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'ha34f6553b8afa5e2b2c9a603c0e3c38f32233b6e4ab516894c4c1e8b15d5e8f0982026a4a1c2ba025f252bd1f2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1d5dd55103f8cdb63d6ce68190434c07aad6b02f0ecfde4d548a62c2b4cea8e83c857e13dadc0571203a9589cdc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4c52ae8d53a94d46aec312b7170d33e8af8b66094a674a09173a0d178181d86bf843461dfe3d4c2316edf3bc60;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hd03e7bf33447fe70ac56ca21c0700e53ecfafdd1d6561ae19dbaba00148e28e9068b3664c9e4b1fd41386b41b2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h112798cf57c03ad843164fff11379ee89be234c8efc6b60821410c0cd3ef8cef082a656718c207bc111a95cd397;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h76db4a081053dd4c0446cdb86fc3d20a0e4b580c6e3a585ad231de1f4a00b19b295916180cbd9ed57123033f51;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18f64d4198e424f6704e96a6df3721636f580996c6c8153f74366074571f6540ae5c30b27b5a5fbb23e0e0843b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h18b3e6b3cea0be1d56720371ee74f9c6bcc5efe68f5fd5803c8c6857ee5e39868f771a1a77282e0648daaf0c7df;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15d253d4c0c6679c13759dcd1a6d612e53b53d4e9c2e1d71e3eb240bae17b44e850959a0b8049af88ee3116c172;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2f86601ecc6d1eeeeb620b54a5f9d3b90c6559381a3c97de6e9f26777532759fb5b5dd4acbaee6346abe961af0;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h848ec04904b617ccb1f481ac9dca1182a29498edddf0d76278407d2e54bd4bbe137f2c34c47d1df1b79697ff29;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h4f99207f95a8e8e4bd0f109235197249a2803437b19075cc70332d7eb7e1d56dd1d9d8ffd3b91ceb0745bd52a2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h2c3a2136e50912753c35e90580a8e834abdff435b3265c6e06735772898a5b3197a6fae63cf6d41528a3b46e49;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7ab63b29dc7db38b80314b53044f74f1cf00abb785b4b24345bc6a43fa9f7ce7e6b9cad46f890cd85368188fb2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1103350f6e9b09782dd1f4a5eb82228dfd637f56c853b5480a1956626ee14a61f499d905fde667c2f495281ff1d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hb7114a22a9ef351bd4bfa9da15321dbe4c73afc565454fe2196573c27c92397fc04d7c0ce80a58e1a415482986;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h62bf994e0cacc7febdac7a4b92c05eabadf55e8fd6af0bc4980974760cec77bbe2cbd23dccb7a4f685e6f4900a;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e6e84e630883bdbfa5e418826d7087029aba30624e8ba06c81ad02a4505969fc63640d9f5fcd008d4ce051a363;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15c71d921f94c47cad7eb01204938a928c73fdd791edaac5129a2bcb9d58a9bc36e3be00d9d705080bc3ebf056f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'haf3f19d9e2cb73fc1c39d24f0cdf9c76c9c8836add4118e4e9d9feba7d9ae19236c3451a2f41e135a5a703008f;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h156a6e09f53b66e3dfa8126e4f0c2432d284c36163fdb8da6b5424c05c6764492ca7b60e2e48d33dc92ead1594d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h164ed685b29d39764ccd413c18a3f82e29af4cf5d2583dde8a26e982e62586e9da7752449c53c2d2c724c2ed9b8;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h5f5bb993c4f3df3c46efb0831ccd8bb6abf4eab9c6f43e0acb2dd65e9e701c4983e405f8cb4c94c90dd87da02b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h10c13f30002a6f21d123e2a3058aa0662fe50a08e426bfefc59b1218e4abbb15b44976c74ec5525554a7b2616f2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h150a64b17ad61c8fa2e6fce0c4f7370761ab7c3d37a3d343a7c682aa7ecce368a69224036df6afff64857a16863;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1c27f2a1e0ca67c52a765bbf2bc86fccaa2200d3f5e061dfa60fc3fedab16c2ca5de3e98f648d88b6f1ebb62a07;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa1329efbe89c5dad87f97de4634c634c1e47118b8be600c96da8d0291238f3f89db778df223ba3e192d34b581;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h3f232ad9f5138f36c87411bd7b263c73d58c1a9971d9d5e3ab9141589a9bd1c892144f812fc998bf5ed947f839;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h13ac31c3cd86511fed87e05b775f34ea32b7e2ba19bcee5b25a44275a7e3638fe2c132a7efc009dd3d66f2b530d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15a7afffc942ba7c786c67f905fe1c38b25253db14987ddf2f92ee099147dd2168e976af1cf40e744ab23fc7c90;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1cd4d2e7089d88b4d4b94a1c59d540d03f453d81bb3d5b2e9985e8bc343759d8acccb888ebfc841e54394f5c7fc;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h199bd1901f336cd40fe953e376d7b60dffd4353116889a287c0e5f3f87de18cb5bb0ff7908f5f97438ca9287a25;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h137dc2561ce7e03efb277099a14d9414bca3fdabec3358b5398882c44f9cd51bc94c80586918c4e426e9ce816a1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc80359bc4c58b2170119ea4403d3ead21aeb1cb7777e5de27c2c556427654852d26317547953c269e830143c2b;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h45beecdf40968d6ead0712d17db9a13929fb72ddf88a7567fff17ef58766a2471b60147e9e642ebd16f498399d;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1ed5e14939aee1918f68420d581a40b4bd93b20ae7cedcc96f4f3ecda46934b50a23342ba67b239ef347af88f3;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h101d5920884e05051b94fef3523d41ad5ad39f5cbc5a353ea2e672c1670cf5a484bc31b98a91bd15e8e164bf6b6;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1aa2c9bfb05d92c96b322368992c3818cacf98f2eadf6933022fb6ba70609aced2237fb3d8e8edd7413a723c899;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h11e5d5df9e10af128a8eb7ddba9ea5fb127973392e6ec25a640b19bbe0ee6abdecc16d9234a85a5ebf5335b6137;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h40216b05f8d0e177307a1353e2d923295ad97baaf53bb63e75471621e8c008d7801fccf1346fb55d6a250a97d1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h15b6f8e41ea39e35cad6ee6cc0c295d2853671e4ff380744cce6a051d0a3389fd7344467d8abb422b713a9bb2ca;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1e143133db325b4c2edddbc223af23bf588ad76d9ad809562481225f37b9c44af3066a756a6c6f0af8156afdfc2;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h7329e0df2dc1e7cfcdee94c4e3a9d9837a627a007366230e46c67338709926afe49389578596ae9565438958c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a99c26a58a6a2f3b15ce9978e74994756902d8b082bf66b4886187fafea3ed9108b94569c41d3c9ddd81fed628;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h193f2e36aab74a60b53ebda976f8f1a4ed6312601258ab654093dfe362ae2cd328a4b4898fff00198f9c76c348;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17dbf6b04cec566921f089ef03a357f425a133d3cd420fb5048727d604fb204e6d7b166d6b304dd5aae7d862c47;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h122ae7b2e6741eb1f6eaf23b131b17f7d0fe680d504d734f473a2662dd4afdbc6cd59d5f980f6058696792f01bb;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'hc7db9b8b0f0761f966645e78042bb6b0fbbb0fe6873b143278d83901413da9d98c91923f5ee9a9b48c40375678;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h16716acc32a02764c60a670a0f201ed43d8009d25995be024f083ad88f64e1975ea3b11ae1a9370e6061966030c;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h153266ca4fdfa875ffd6ae002007a617656d686b2f4b0016047c265ea0cd92b676c5292f6aac3e7181558c47298;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1a3ba930c3cee6bcd30759cc083daf2185ea768d687191c0e415a58ddb2e2977760ba9bc49782988f8109a44d26;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h17906c026d00c2fc93e118ef7e34f96fd4384645af23f02a8894db85843916260d2541548de4900fa0ab2055eaa;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h1f76184309a571f8409b1d6e0cba59feee9aa4ca5e38237f51fe1a2d71c54e7f3ab5daa4287bde5b1cfe0714ca1;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h117497cac008bab746adb53aa8cfe8be6c643f2c730c44350bda078e277b68882132ba153fc1898d9eb32bba075;
        #1
        {src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 361'h307e896450d19ba5b7df2cfd2b296e6db8861ce66c8ee06cb7726a8e5e07bbf693235566fbbe2eab107a413aee;
        #1
        $finish();
    end
endmodule
