module testbench();
    reg [10:0] src0;
    reg [10:0] src1;
    reg [10:0] src2;
    reg [10:0] src3;
    reg [10:0] src4;
    reg [10:0] src5;
    reg [10:0] src6;
    reg [10:0] src7;
    reg [10:0] src8;
    reg [10:0] src9;
    reg [10:0] src10;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [14:0] srcsum;
    wire [14:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ffffffffffffffffffffffffffffff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14738f87b56943364dfdb6600d2be27;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h190fb43de3d274fabbcd9ad9ecff569;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16b925f711daa9f2647023c967b8bcf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d17eab8afb96ab6f06c687a77cce3a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc5caa56e2b25889d6d7f9e4dd74769;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1760e36b9d8092f1189ead732a0e6e7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h156e4655c65df12a8290b58dffd04ea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19cc70075dcacf4a385cfc5dfc037b9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c089829473a6c345af753be260096e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d00308335e5d08f4ddaeab0e8afb0e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h158a55314066b45dd171c5d9d73696b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6a228d1768c6a0b38ddbcd9e068226;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h170320e7dedbc7961e49d1377f17e05;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6e9ad3a76eef507048cd58114e08fe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b05d4448e01c589d58366f327080aa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14589f90cb20972ed6c6e1161c2baf0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16b433b635fc69b3c2e7980746d6543;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h174488866a0059a17cee89d9f367579;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14bf5953cb3325dfb5cfd40c0d5df17;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11fa2b9d54d36c5a5830993d9e27b1c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb6979de350f98e6d3f6529e6952c19;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf95cb246d6b01bf8bc314fd11e0e83;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb8d08aad981a085ee72fb94c9048ce;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c7cbdb6556cf40d0d12c77bd169056;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f24cce0ac70cefe2376477f53b5240;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1df44394ed3335bdfa45a3d3f28e616;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ce99060ab905fa89543b04fab0ce1c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hba2fa22443156b10d73cb3ee1b8d05;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1978bac35b9453363056269fdea7ad2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1827dc7e1f4f876132db07d24243fba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd2a37229f7a0ffeb0270bde67a2873;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c774a33007305936407a3fe74e6f7a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h148f1b248cf093f35714b01b695eb16;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcbf5cfe85285b85d2715ab62e0c4e3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f1056d47f0bb1c1cee1bd66f9c1ff9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9377e9ab10f4c45ccc65ec9d8702db;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16a8f72683143a7eaa3c10051f8564c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a0bb68b95249ae5cbd9bf5612e677c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd2f37214bdbc1134a4207bee2eeef1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc96e81f489723928d0072b55c7fb45;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h184dd8a35aad3fe1c9dc1edadf58178;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h542b6719cedcfa94a7e80c63318600;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fe1dc423d467b180dd3aa1db8a295c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he1e793d685ccaf0eb2c6f17f487a19;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h127b9478a44783b080a25ee9e238e95;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hebcfffb8e7e0fe5786fd63a4e8d670;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a6ec56b353952b0dcc7c6e21a0e607;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc30ff04b09c474439052fab1c74da9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb0ddd91285f5276e09777cd83bb81f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h164594cfa29ea281aeeb51da6aad808;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13fbee90b810970dec7839666e3d829;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e4221c6c078fcfddf9c3698ffcf298;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h553742aea7365b34be1ce87e0b9bb6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15bf5f6a19da32a59f35737613c9ec6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he6c5ce4da3b75bd06f4ee8b0086a6f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11657ef69245412ead0c7e8f6bb21cb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19184c677701986ca224d4ba0d8d231;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h74f11817e5eb27e193219a515a546e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfb110f167a18eec131d446acf6d30e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha5a110a934ccb01ac685a4265b786b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h129f3121b4c6b9ff3e36b057bfe9f5d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e948cfd4362ccf9c9b949cc34b3265;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1746e33260abc208eab969e0b01c5f4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1009b3b4adee2bb1fe13f15cc44cb2f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14e71af34a6287905ef1b895ac4ad8c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h24c287fe74db590c7f16e2f230c047;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h92c1ffda6ed1c09df951fe00d00f0b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcc7590cdfd368f2404c124b67fea82;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eedcb53f2cdefd4df494df8bb60ae4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7d0504071bd26bb6167a9cc9689a63;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4c48699632ef9432c9d6ea4d2632fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h459b4cf3535f273e91648d8f408175;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10890403c0b1df19bcb117e0c80f919;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16e864d9bd9d8be878d98db63b2721e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5a0af41016017fbc61533f71679cf1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1120e12fb71e3dc04e6ad9c0408fab5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c7ba8eb896301e2bde5b36f8e22fc4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15b1f6b6320779e215890815b96ba53;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb997f5f228359d42ee6fb7bc53b862;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13091d117499450a3f72bbdc12c9384;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e2d5ac44c33779623e6e4209d3492b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h344727db6277f3071714035c41b270;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f79800ef33f621f0e1c79ee360757d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bffd8b3dc4fb98de02a137a8a21c5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1da95e29ce1bade1b8c37562a477220;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbcfe4608b9a443d8179b9dea7cee6f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he431dca356389ccc5482a55911f86e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e6dd94884fecd0ba555a92ae1c80a6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hde5036ae596bff6280a0e282ad636a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he41dafb4fdc8b248969e8955b093d2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hae89a7c2398d9d9e1cce52c0596779;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7c2041bd45474b99a2581b55d81997;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h125db58326539ad411d02c6e7275109;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b0ef667ab21f27e811aefad819eb9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5dc7030575a42a1741ac07d931913f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h142612de6b5faaeefa19a3294413772;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h134b20e0a69e74f60ff56e30b49d135;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h287f721e7d3e8790c75d558ccbd86f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1098b76a3bd301449a7d8a7b6dc2ee1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bf5fe821e232f459fa151025605100;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h321384c76bc746ccafea13449b3039;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13cef303c7301beeb8c5759ccbe38f4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18e37afb5bb3529305f33619fb3f4a4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf9bee37ae5e8f54553f73b8246e0ab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1000be6d477e753410eebb773cf6dd2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd675fdccad411339338b220243e145;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he7e2a54cea3bd1ba18719e01f7d8a7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h106ba1dc59fea3c4374c2fd4a18f594;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1061efdac0ae79f4250fefc3fc9e3fa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d29ca6a523d5d659e93829f4e46bd8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dda3552241f20c3e1b5d40d09dd27e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2a61800dd1d8ad1c48f485c5187530;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h254ebab8ff29d792735e1e749c3111;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h28aab1ead2a71d386fe999a3d8d828;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d8a44430800a84efc8f8835173de0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4bd03449d65271e884a199b81bc3f7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h100636922330e8623a5f7ca503b2ad1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h186600965e462702d0a2dddbf18528a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h545975c26915b1a882621eb8172c43;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h158fd1f0ef65c3e6de847f94c497de0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbe0dc7a3f5e943ed88822e5ccde78f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9c0b2a0c8aca5092599b4291cf7c5a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dd4530b1d71230bd2362185344dafa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2b442f8380d16f6825c10cbca54ad6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h20709985c85d6888cb616ef969101d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12eb9efc39c8dd72f5abf739812a8ed;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h112dfcf1d9b50be119114d5d230d8a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ae3d6434f36c929fd0f08990514eb8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he6d90d07f2bce1ce40bced0391eb83;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4587c5c5f7bdb3cd5e3a13275a994d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h45d4310ce345f260f503bc07fff906;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h79965d79ef55c345a5dabab3ffb962;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h166855427d8ae70b89f79afa50aa5fe;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10ef673eb80ebe1b491d35e5cc6dece;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c03f2a87fd84e5238522d42ff0dcb3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf096060f04f9b90c05879a1a3ad721;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h138ef5f641c03eaf902827b8e940582;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10cae2db029dddb3d39c0d4706159d8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdfba78a9d1be9f09d8fe197e67d410;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haa2493729feebf1337305deae7e702;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c43b3f6e4bd064b0172a028f58366b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1628a5c1a4f0b69d8375839f521bb15;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17620da06173b42182c7a6a4af506ec;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1969ec4cb3898d560ac86645fe38576;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dc446887ff04a4e6026a697dd3af62;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1deaeaad4dc59b6ce97d4d5a1e76695;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5af9210388aeafbc58eaf81bd943bd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c1e48c3ee295b88aa1ef6e915c80d0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf95efca6d90893a04b1a9fe2b481ec;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8e479b7c38a213764d07d30c1cfda8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13cfbe96d484093030c81a52e78b4fd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2d0ff087793b60c5f743b686d7983e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h427e6a9279b665e558692d43f57967;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8160e4a3c28ecb55f1ccf2e6018d8c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3f10c22d31a009d0756939f485cd9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hca65e8f66ef1086130ed50ec1f7218;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16a6e992f62cbd8c1b64ff066044f26;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dbdd691710fb06cdfe1123103e1e7f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e1b5808729290fa6d3891d56bfa877;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ac836f016ba0efef36e471dcf66f0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1df8895a4257198be95fd393a9bd84b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h148d055d491bdd936fa6b2d572b3dd6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha3c728ad3bb0f9f141c10b52c67e49;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf9bd595e5e457ae332c3ebce695b35;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h127fad868ef179326a176092acd43cb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13ace35665c9c801091dd819ac50fc3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h63b4896c8acb627fc804ffa48bd2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haeeafc648a89708c2b8d10202adffa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h828de2b874598ceccc3c7da60decaf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1276da19e021787584a5a2470a0deb3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11582d4a2593e51df6f8f4f5a0ad18a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1095c14224c27da9fab7f1728c723ca;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb96f2805e1c6cdae62bc1d42d09cbc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1461c2a3e4e982a94bb26e3981e2805;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h193d7b1b171b72d4c42e6e22c0b01f0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h42f24c47d458bd4e2419c739478677;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hca6ad84231d04c49ea067e6dde2a7a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19df13bf24688d80e8f116d05efe9bb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h602f0dbf121f4efffccfa71ac33ade;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha8a3df9775174fd2b0f2293571e854;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e153dea908e5df99c7c669f2172bd9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1270063aaa2096b2de12fd1faef94f7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h27be7ded3609a41aa5dd640d3dfd59;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'heaed2106a99a5214b3465d0e04578b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10679099a2660fc065615fbae804952;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12753b283a4cdd4ffeb32bea02a5263;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hce706ccb5dab6909821005b6f923c1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10ecfab967f551ab187de16587b8a87;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd14eca42d389ffc98e00f7877a781;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12bdb738e683628d63e57c68520f7dd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7ca27ef4ceafc24ecf408131cf1c40;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a85d3f3d276231f5cc944efd61ed04;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha9c1ff9b0b2bdfd7cd17e8ffa72bf0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f9abb22f3f0778152c040a0a127429;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h148ed1d141d86f5f4b9ccde4f3f54d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e4ef5a5fb00b998e6817eaa0441f92;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h78b0cf5df31619d3f94a6262abc58a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15c8771e15fdb9694a70a9dc44df80d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12f5295ae3e44ceb977a8ea7665d358;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc94c2decfe97d15f1be8da27ac182a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h174f5be8f261fca83eebb63b31f4cbc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h31065e47399e23936c12b827609040;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1285c23920be69d0aa9ee380f2b27e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7dbdfe5a0f32a33b902b1b10fafa35;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbb8825058f0b36aceee0b2a85b0119;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a5ceeeee9c40e14917878631c6fde9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe57ba471cb349aea5398de3d09d0e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eb89eac6527bcb039f0a312a9a5826;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbda35f9314c4dff40e053594467245;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h118f08bb14d992f14ef91b445aaa25d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16d44b843d4943626dc35a7adfe70ae;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5845f42a4b9c51d00743ede19185c6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h112ef8d0d405f1c19f0f7bba518591c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc5ce63e66a02bdd98af6b2e969db15;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h160f4e51167f4908f9508e6964e3712;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c4e4b582562897e17e1594d9cce29b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11828e8a97ea7fad6e344fd68673f83;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13bcd1675436250805e1a8283cac959;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h767da0eb621816b39ffc0c8ee78e4d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ff11be6675970bb2da7d0a93c843c3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe549bfc08cca21ed497c19b7ce4e3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h583387b1396388a64b934515141d64;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bf27d2613ccb555d4256d572616a53;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h998cc4f4107816890fe1481158e01a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h86e0ce7afca1838c133f2ae71d6f95;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4aff647c1356f472cd801bf48220bd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11f63d82d08d6edf4194daeaed42bce;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha597c5073565f2f01ac1efd365d543;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc4ff39bef66dd92514e53142118164;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1530426084fed253fa1d9b91932bd0a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h110e3c10baa33f007fb17472d4282d4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb73a64e5cbfce174dc826ba7d75ac9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf14a2e2ba692c080b0618feb01b86b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12f245d54db2b1de8f86c1bc3c20f8a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bc80ebe7f8b247be65d5e2ddf87df1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fabe72f040246acece9d03541f53f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4ce8ee53d991f02e3d07fc53fe517f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17d08b2ca52f054f1ee7ad2323516fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1435277991795c353a367821b060448;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c0a2321721bf9460eb6a1b4cc49af2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc47c13a6bd6510852a6270ed75c32e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12a7df943a55d38dcbb4208f5e40ca4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haaf5c096f7de7f5900a33b2d7e50e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1321fbaa6b7f1b3976f7a2d8b22b78f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d0ad13a58eb2f1713cbc3e527021f7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h46bf790435e6cdb7005bcff2639aba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1be927030f9ae9144061dd4d25b1931;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h933062d8b160bd432d7612012494be;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6a730cb0ac7cf108caa6c2d75924b4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb0fb8483fd337150a115a01bc9223d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8380536d7e525fbe35e4d94b601b02;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c7b4f761350c36ab299f80e7f44df2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16ae6f4893d3fc9e2cb8659bc0fecfa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c3df4251a122ae933e2d2e1d2a4f03;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b84198870c1c2b0e694af53415b5b7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3433dbfd66d51f28ef84c4734d228;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h654e9d0df59b6c4028be86c65db481;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5de9cc1fa6b6b063e73e2c75f9f773;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h117a6b8ec88b337a97a135b66db2679;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10ea2215dd352862f18b19516404b8c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d94c8e3b0e98f1b252ed673813ad9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h43e30f6bb31d08d215b76745b92549;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h933cbff2dda3efdfcff79be97f1fb6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11ab1fafe1bb639b90b8741978c0461;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h50688fbf555ba6e8930ede227f0c5d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbd1e389218cfd6c5b5748bd4d95243;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h145b00f50efabb7f8da13d8621d52dc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he9220cecf09196ff1d593840c97dff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b51b83f76b4448ed9e7eb46ba39f11;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c7a12410b867cad4b3df84b6571971;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1574651bf08e30e563a4027f48ff90;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12652d20e18edcd18d5e9c169ab7e36;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h148642b325104f323560096dc3cf47f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cefd53f0a0660c6efc45f3690fcbb5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7809b7ea1cd7c144f3ddb3e504c347;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12ad65450f96fe51ecfba846cb2f058;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbbeb6a55fad8c589b9581457920dc1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h101f9fc5d6eb8f7d9960ec4abeb0101;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb19e95900eb9cb28a0504ec5229471;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b2c263bf3a0f14657fb17415b3cd3f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9db2fdd903b86af944de59a0f62ce7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hde99367635ef2f18a2621e4b34e4b0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3834f7c743c54058ff913a7c1a24d5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h24b75547a53173dad63feeac60cc06;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10ebb78ff24d657d2f311f381588d26;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h459e65660d2475c3fba8bae24a1817;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7f829eae43e35be451c58c745b3d64;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19cd446c2a4ab3ef51b83724b8b47bf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13766ceaf9bbc8320f87cd34976ba50;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hee8e20db87175b78c2dc720f2530c0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf63790ec8dde75d364846b295730c7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19059d69f0b1119bdd21ea8d75902ab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1409b5a5c5302e4ede77e1a01807dca;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13c7ee7784efa6e611e4035a999a46a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbac10092feb3dc91b8ef4ce4ab1816;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15474516a41e20c3ec522f3f67d4168;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a9cecf01ca68f43144e88e5922aa55;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ce3e11f241bfd6b3e34865884d9038;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12b64b8c77313a5043ac66ff9cdb5f6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdbdc9f700bdac133025415b7a9353c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4f710844f433260de27021209be444;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4028de72b3415d68103d19052f98df;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9ccd277280fd4bb163600d0fb31ec5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1238ebe10e6cc653de73751883f0550;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9635d76d68cbf438fc3212620412c1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10181133589fa5257fe12288c0f1e09;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9fae3c6f57fdbfd0a85d6f2292e74d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h84fea7406a4a4ec25d25d4495a5b31;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc316cecbfc131f683b0153ef5a3f43;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fd7b3efb09d8b0f8a52be5f9f29d73;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c6f61e0ae3447a38e0da821c84dd13;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14d61ecaece101faa37042033886e9e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10cbe3bc40c7288923db57987db41f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha5188f856747ead734654ada675651;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1539f5a745b31b10d6395546e8a9ef5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1558530d1b5bbe1925f0d91f81523ea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h140302e193d24d7b90ceb45f1b2ce7b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf075b5af6e04d099cbb637a346c5a1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c546f450e75af61c27ebc70eed7dcc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf9ccef77065a3658901fb164686ea2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2928fd30f4ec6f5f63c2741ea46a61;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haf2f1db77f533ba271cca199f4b745;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h870c2178176db977d7a18361975542;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15b611291478a89a50b99bd3575b50e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd4dd56c4c0eba19be350caad02cba8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15bdb2b96f0e2860894ce3a16590c15;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he764b7b756c6ebbe40ca98e67da168;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h105b57da01aba91f4fe92b5dbc871ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12c9a4a9edcdc691b672c0de185e24e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18f4d6e2b9347250168725b97d1a43e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d9469357370b02d40ad68aa32ae5a5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2a20517deb6830ad6f8a7973bd9648;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ac4f88f4f1373fddbeee3c10b90ac7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18cc9a3a6487dadc5fcedbaa7079f34;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7a69253a8f7970065eb3259fbfc747;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13fdc385979cb447d59c34142d69f90;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2f9fbc2a1b419a2b98d32c0613983e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f1afcb81839dc463c9690608b5c49;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hab22aeb72bf3f03e3eb96812eee97c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6d21162ae139e03a6e6e8ec13ce057;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha847772815163a788d7112fbc003a0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10838acb63b6ccfa71dc7ffa53e3bbd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1110fb9baae1bf2f6d7e5052de18e1f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h76b15e8e611e8b6ceb892c49696fa9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7407805cc3a3ff4aef05de1ce9a26;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12b91420932a081628f6a8dbe0f5221;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d93a343ae2047973db565336d9cd43;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4a741a5c183e6e81a4237565aee35f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h111d205a5401dd7983355516eb43fa9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a12c4dd31a1ba9b08a6e39a3d3e87;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c8fe32034c282ab2ea383a2cc59702;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11918cd335ae4ff81662fd7eeb5c33b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5849fd5571d9cd82d35e0828ecc064;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14dd8f577512aec5fee78d4219ac477;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h91a4eae37127bc9ce8bfa7a772acf3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb493142f12e704f2f83392102d76d5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ca64e9e309cdbe65a042991538b5b7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he52396a39cb3c02a378c9c13029bc4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18f814ace84320609d2e0ad9874d350;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ca551da118128460080d35e4ac252a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfbf5e0033133a70c5a5baf78931e69;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13b939b6515002aae670cc2976262bd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a834462883a0244360b13497bea889;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1032763da46bafd0b1a4bf135c25e38;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h123a30aa4cb9bc07e2b645c87da7a6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c28eeaf7ceed4594533cfa7fe5e386;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18bb3a4958aa040d338f6b9a743e423;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b711dcb0a4b80cb1020c850b3f49d3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17c2df5a3472e2e6ac5ebc794a8963d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h77f466379fb393b1b5efaa09e94fe4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15f4aff2f591133b6c2cf50c0199e56;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h52e693c4c43b10c17af055e72554a8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a34f24c2fcf161b11369f82286f4bb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1caef28010e1e190eeb53d99fc140b7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6a7af22f87748f4865d01133d39fb9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hec83c5fb67eeb4aa9fc307815c4c75;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c9145fbc4509e5c48844bdeae1cc84;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h138885c96fd539a1df529c8102ddae4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ae9081190c5f63a39a5f68105fb8cd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h180b70c2a1b00d6bcf8eb4869de46dd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdd06789fcdb497076acaeb137aa875;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h525569365a308fee73ae65f64281d0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hacf5aae7a040434661cb6897c541ff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h77f50b6e5202e9d32bb7476b318830;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ae159e20827c3ccc4e873071a4baa5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a4ef5049a472eb2e9bdf48cfa448fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e66cb983b9e02621de5a453e82e279;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d454931c9a4a6f262715630ead1664;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ec6d8697426208f11a05a38c5cc426;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1353a2fe2f10e3ac124269df90a5e62;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc76a5c6e01a76eb3b09d5f5e8f6e7f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13232421737abe671d5bbecf3a20688;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11990f9bc4d0bd418bb68f0be5f6eac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h35b88d83be998c4618f37b2c43505e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7d885acef82cbfddb1ffa69bf91f63;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfccc0b82cb59fdfad4b7ad1d911c7d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h30b64a7c296f1ae9eeeaeeaaa9e709;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b0d4869413992477d6d9570bbdd249;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf143d0667d8ab6f8c9f6f2dfac4ecf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13fccc1129840dea091d09940d6f439;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hefe65274b79be19ea9c82f23f66818;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16114616c96e0cba62fcf1fb0f0e9ff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18cf18c561849d808e9c69d440db4e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha158c9448912f36bd357517bc7329c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha922abd532f76df1cbb837d246e0dc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h54b3c24e6a064cfa8554de2fb29c7f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12933ff7b9298a9efa76e429c1c6fb4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e0ae1c5b97be4b144bae116c6e408d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7078488d31e98e84aed52b18582894;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9bf7c1ad08bb1312c77ef74b285356;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15b05476fd4df2d7664449287350f96;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h748bb93c17516c68266ab87ef6b412;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h112af51be32e6a0cff2f7c624ab1ca1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8f5f42f213f50cfd4b5e1cd2dbfb0c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h161198f062c593d0fb5e111635c0d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb00d69cfb7ce47bb805f557e6985ec;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1236ab66505e9a8838e7f370524bb4c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1765849468c95a749c5626692f60840;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h33bed59351ffbeaab6cd57e232fb0d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha241fd13b36814f7e14b586ab2bcef;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3110441cc71e6ef1c22beea2bee198;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4177b73dae58acc26ef1ca99711613;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a10189ff3930b9bd7c1a6255ca481f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd5aa4c3ccbc3d9f00d248f809b7e19;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7ff2a312a4f47b9af0634b240be736;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10594abff5c55ff4a1a77a8f0734f8a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11d33d824f89c0a9e0bb9c827e07bc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ac49629d917e830da8fa0a78e3098b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc4dbade1a352c73a5b6b427a2c9a89;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc5205bd7cfc2c11693b1b8aa1bc464;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h823f2d51cad6a065a3468bba28b8d2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h52a99ab3fcaa3d1cb9860a80f21e99;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8acfd37587d9b3823c1323de4b422d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c2f3fadef462288a5483c44f829856;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6e1c07e462ae19d0233fe79b319f63;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7d5b27a54cd256b5160e3078574373;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dfd809f218409d22047e028df4a542;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8167773fd08367fd2852025dc62d7d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1013d72db68b710acfae3d4a6d677e9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha94f556a2a6ac53bff83341b8eef8d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16705ae5c59811cbe459d4fc88e0548;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19fc4ef8a37740318ecc28c067fb25;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hac735c1b8768e5cb1ec3d2f8f92eb7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bf493dcdbfa6732c95fae70b84d2df;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd3da8a4c2340aea52b2cc3f4610e08;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1701c5ee23db34c2c4340a1f7a04d7f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11b18a8b2faa71673182411f15ba291;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h121bc4f9fd578bf6f1b4b6cf6f9852c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h163c8b3ad5f393427afa88c83430659;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h152c9375943856aa77bbaa9f84efe27;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bca9cdc0672af88fd66cade75f975d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h833236e52a8fb979209ed6fe59f52b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3d1299d489aa550ee7c22ab0c189fc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f5301b5e178fc2f13c9f298ffd68a1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3a2868adb2d9d225ec6047782ba3bd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he0c4ebf5efe5db335d74f2d42d383f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10ee1bd0fc5741c68ec63e0491874b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14f2767f63658eb7225089a986d66ba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ae67c380f53ca113b8618e104e2a15;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf408b60a1c1e6396a764a587456e75;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5b6d1d35c47baa776a626340ad90e1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1acb543c490c59f77d53c927ad0d489;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1964bdd70db7ca4974a1ac7433e445d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f25874fe6e3304890f2a371cc7e212;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3f960251cb69631de299aea1c7c343;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12c9717b9fa3fe8d6c5dbf542ed9f9c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbf64ad7330078eab7185bdee2c99a4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3913d8494a8faec20ab1729148a549;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8797ac7d0a0a78ba550e03ae5be74d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a87778eac64dd4b6d798aaf16493c4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h119ab626ea3fd6e84f9318aa45fbdf1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h123bc640f410a426ecc63d5885c2713;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h89d225471708e6898392b1047fe034;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb4300a14189384dd0edee8d4682107;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h94113c54429bd6e4316c388bfc9f81;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb5b77e078517a1b62a2549bfe1b928;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h828a90b4b2085b48a60cadc03f60bf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf32756b8a6a5d030e69a46d9130621;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5b60ab4dbb4d8621793d593e59d84d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdb87d17285ebdc5ed179bcb4277557;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19d1d18eb834ff639023f17c6f7b834;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1607416f6e76463c3dc39a23a0d4efb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc6d10fa009f44ed71a97abb245e49;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h169f15bfe074f1e3324e90a0d89872d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5a6608aab5989a02728b88693789b6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17d7eb7f55b98a0336114ec83bfc0a6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h280e908f71b854868a8740ddda91b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7091ffa01489d1e1af9c5618ef3bdb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h154ea0de7ed21198c1a8ed6a859235d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1461aed1b7c40bb4f719ac872183776;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbae6786282d277827a94146dba5eea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1307b653577420936edecf05cf01254;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dc598e25e1d9aceac29bb7798cc99d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h72ecc9451262d6802f9ec92961f277;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10c7d16594cef4aa203bb2b95c12a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fdc8c390a1d6cd7352eb326ce51034;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18a2dd522f91300c385e3480522bcac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6792d11055bec8de6fe94a7413f829;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13b17c0bcb13571648188de1db61395;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h859351ffb8a9fcb555f4c342cacf0e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h109dcb2672e8fabe7e26cba1b8593e9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc59db46b0a2737197438913fe643b2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h853e22064e41eb3ad3e9a546d7431b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h254acd10393ecf314909edcbc5e6c0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd15092798c03b197c562f99b25b606;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h842631b5047bf4a2595622535a30f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fad65f9d129c1d653b249cb0016e60;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h154478d9a4b09a13facf34cfd6f92a7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf2260be31e405ca4fc6ca8d9af3a06;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10c1a7305c309e5c0811922a6b034b9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7c5f0877918e42c7350c151fc3450;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf0543451e3d9aa127c85b2569d114;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a2db6c3a637872e40ef178029ae8c7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h23b32788ce62b268b27649e16b48d1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11ae737848202ccc32fdfbcf5dd380c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d50a7fc6b63f9d60a939852b06f7a8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fc7e7d51e3f67b91ed4d3b23e61cdc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b0dee74396661423220dbad8f2097a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcded6b3738a8bd2bf7e3bad2690650;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f6e5d0469dd1b6d9ce8de08c066092;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he67fff9da7b7efec0d8e42da629317;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b4b064c99e50e96b760cd85ac30255;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h33417f236aec9624b381c3432d89c0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4e34c16032c9aa7676d7e4dd5933f6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h131ff846cf90a829069b2c9a1f10d89;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf43186054e570f52d4d408719fad31;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d1be0274cfab19c886d00772c8a03d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he50f12c7d5aeb226f38ca4da075ce4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb20ed1bfe4e8ff46d33a6cd87b73ba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h75b7c31c5efccd4f1c698b3dc02a74;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17110a2e303c936da1e4a25897355da;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d241eb12a370932a316b4b1d939856;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd7f79958a817e9c2ed660552b411f4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6ab68abe8053c99dce5c6714630cfc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2bce875c8bc24a05b233620ff49cc9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb4e7f0336f7884562eeb093c13bdc6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15923dd2ee118872124c80c9c35060c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14dbb25e6c8941576013a9011432871;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e89ba54d6d6d6bf4ff959a2cef1824;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bac2fb3267cf4dbcb5303d5786fe2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7da9ba9acadf2a628a6ad4a4c38539;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha18cd9d39e43cfac62e575924183e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7ff754dc95d79d468e6b802f2e9e1a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haeb7784a313089e509ab32a3d0b686;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h123f2544e5f6c917050f9e9b3f35745;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6acaf4b1c22ed590bb4ba36ec616d2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hff31553014c01a49587530905f4f4a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f477581777170212299c3b789b8918;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4dfd538515da68f0f4431eb6312424;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf8c3a5c28928fdb33b3acb68578d49;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c3e839f3c70f2ab8f3b4f12981911e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17131360c05b4ce993edf68186b47bd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b0c2135d2a6a829ee4c4e8a71fb497;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h84fc1eaa29e9c0e381f3b6bb72ec63;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfe0131418fa5c5d329a35cc73c495;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12933f5ca45c0ddae821df45007b003;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16064a271bb7c7577d65d7dd94ff4ac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h66b567a860f1178e55e9296077270;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ee33bc9944531a6e667cd1dd483108;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd1aee723f0b93ebdac3a8225b18682;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h148bef994766daa4a30079ea7f2ea12;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10b5f8c7590dd5c03150cb33df7e0c3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h28ca8f487d01c998cf01431548412f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18a52c173b8426c89afc695579fbfe2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h104bde2b5c6dfe5f763c31b9b2ba6b5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dc6f9129cef27130bc49fa729d94d4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hee02dd0dcbf94aae5caf6e7d17d3f4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he4d1fa86f7fc04bbfb194bd417aa1c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e26d2ad4615eb99f209d682af83ace;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h111505997963873c9c67ea0e972ba18;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha08517bc3d368e4a2f7afb45a669ff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd71c0fe58f7c7cc56fc08e720dc233;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h167a1ea5f4dfa58cfea37cc073a72f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9fae9eb6f222a9d9aea70bd7c4d73f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h147d99d81929295de057e61c860f7e6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc5d002aaa1e7307dd7517e5cc4f563;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9120d454b8ec4296012e67bd23b553;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a7bc97a5ef965d3bc09e4acf78723d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e15cfd50e22589f7b1b1d785e354a8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h180f3e572688c2b67a82306bdbbd7dd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h94618490017ed90107c5b8da4863ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h140b18ffc79e5a0987363d04fe09ea9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16c1759f723f834a20189d9fceae35e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1df021cb18f261fa926722f84686b9d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdbee29024c1cafbbd51c49a78ab534;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9ee3d30d1290e5c2ac8fb00635f70e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1faf2130bc1e6e0fd7702d1529e7b30;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bb643190a19c040c5376a6571c98f9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2629949bafcb8be4705f86ec9441cf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16cdf45b5d331465fb942190ea2e174;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h169d9fd4740a42425e6c78d8e16725;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17956496bc5d808a63c9258c4c86b08;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h618ad2dc7a12d94aafefa8bae54f43;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf4995fb367ec9f006f0027a0cf18bc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a44963691cb47333b064c6744fcd40;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha8d9cf7e953f6cc2d733a16f4523a1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12f075115c92b10885b0b33e4fb9955;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18fe03d4ed4b26e84925be76ffe6c27;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bfc406a538ea40acc6fbc5befdd62;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haf395809d3aa7eba0c3c3b84ca15b8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10f7d60fcf8bac858c7edb002f0f70c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16d030101c3e52952d18ee561508981;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10afcff719e5fff317ce6b53d353492;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h101f292253525d2c15096a01f067ff6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he4e6c13a035480047459ad94ae9fa9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9a30e267cd99f50fb228d0f4f2f17e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h198daac6b435021467c16bafef78582;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h814c91629bdcda20597095865e77a7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h141d483fdac174356a45e34b57d38f5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17b8cb2b6350e27abb3266978a01297;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb2cbcf8a07c2093a6e413acfe63340;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h407e5e5627d90e83d5ba61e9dbd078;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ed5fec875192957ea1f66977f30517;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h781ef51e67980f7d4ebc79ac1512de;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbf2e27077127ab6ad09a3281cf2821;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2e6602579a25ff773ec8c26b1fb3c1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h32ce989bc780d99e9d328e865806fb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h194b296ba7f28a89a8cd009f8045422;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h113b080ccfae9fb89e2598864b1045d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbbb1cbb6bdf92e7cccc9a9e3d47b33;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6fa596f7d98dced68ca902ade6a54;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf2ee9883bcc6c0600661b78ed7c737;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3b6c0900e37dc9d64acb7dc13fe76d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcf5cbc69d22c91bafe50a3608c3687;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4ceaa5eaae7b87eb4818d26e1c1d03;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h978d3ff4c0a3271fe1794771a469c0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5a32d8380f6631f5fa94f477cb4ac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf1739bf0a3d2e7f110e0be32e3c9d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12876dfe4ee2c4d5724c5cf8a743144;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13bf8772882808d758a962935e503e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1309c39661529ef914b2219cea77b0b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b6f8a09bf0c575125ded19914736ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h277b39eb19ebb5ea2fccdbab446ba8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13e3c9af1a6195914556e263d9d7b6a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18afa945f40761a5212db1775f35010;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1274cf74a70874e17f608863013382b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dca900382bce76b66be0a2f227f46c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dce8caf64bb207bbdf9eec7b4ce310;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19694d4f1b3f2b9975227d904e3d925;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7027b7c37c5c4622daf5dfdefa8e9e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbf123f3c6fa7cf0831ee167ce87af4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcfdccd4455b0d36ef79166e63ee34;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4ec286f89ec5f46c7c08499a8ec34a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16bd6ab8e68aa50970cab6971197665;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haa6bf9a2af7cb1ccb5ca5a00e0c292;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6a0a608be2b64bf6b1d2e546e344af;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf56c3a260225a10902401dd91c54f3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e34414f5a3aea7fb2951ef1b3ae077;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hefa3932f53dab21e1aedeb9088b56d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h160de7666350995f3432176ec6c5968;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5d1622ac8950ed82e22ee56c4b2004;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14df811a9d1c326cc3ec12b0f0847da;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1954ac093d4caf997028d79c97a2b5f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e3e936665f3d4b637165e33e549ed8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h71f99e6062c5c1049ec5ad735f62f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb160597029406a17d5b13c13dedc5b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17cfb091db6e66c50a3f14ea816128b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1db2fe0dfa5f47606d46998c43175d0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4c077bac55401cb8803ffaf6309cc6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f35feaf1852a33bedfae0a68ec3f3e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4061e49258fd1747c47d9541972cdf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb3a8a01755305899a275128fec32f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c4aed37a673243eca65a6cd7eb8ef8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1631b3d3d3b24fd8de102f424d3f61e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c5b6a510e822fc577a261dc82e396c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9d5aa552543bd6990d6022f53c96c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha5dfdefcdbd5ae95cd854302b4fbad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15a6faf9c00d2f9f61c6203b6b50bd6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12820504890a13a855d15f86a09dca9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h138093bb09906797d923c0f8430b55b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d88bd1e455e703640e6d5e3fa9e93;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8eef8f615c004f9b992ebe73bfd246;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a2c7e922d3d6cf930246b7f2ada51b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12288aceefce5a96265a394c557fa3f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1980d1bd1c346e9c446c7395c936566;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b04be15ac1103a18e62a4771c78875;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18b38df77ae59e426745a629db33a3a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h139be3b3220111780d06ce30d9fa926;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h163fda391153bbb9b0085172fa5a587;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15cabd38649a6d915112a84fedc387;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15a36f02d3f02777754aa8ee5f6e6b5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc2d1290f3f75194a4ab6ddb6fa07e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fc0112e3e3bfffb75e9ebee80145db;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd68cdc9d2231bcc93d96b74b007e3c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h159ba664dfc392cd168e7d31e8d984e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h715bb6eecc43e7d9bff2d62f6d1b7b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1712fd534d4dbd87edfbc8715f7009d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha5dba2600c3a48a822a2ed60705cc0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cf22a994f60a035c5775dde9599fb3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h180c31b68dc82f715f75b02376757a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfcb4b39b848b6f299bcf75f7d9957e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3e3cd416b49ff642ef402fde62d85f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c8715abb2417fb1ad9cf66400bcbf7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eb9885a13f24e21270917e3e810437;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17a3b08488983c0e8298cf870ada951;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a3932b9f15b6484b1d181dad974aed;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h185f27f2961d9bbe2316b75841d82f1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he2a806efaa14adb8d37128a7c87db2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he75b645c44e9d62e5b86d81c722280;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12cbb9bc451ec23ee5774755d006655;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aa386c6e8af9ada73449c6ce98d0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fe4f9ed654d7778c167ded523c3cee;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e8269692b9b07e55f4e2165a9f7262;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ddaaf122183478b81d197962a3a450;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aea8b09477a75d3d909813ce91101;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hde46355684c9d95ac43151d3641cd4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1277abcc75e0accc615dcbe291beb47;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16209951d7d3c5672dabc8e0a314955;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e645c7922c83744fab6526e8a76a62;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hac9a31239e0d2f52fe5a3e9853458;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h16d2b518f4f46f02225e618e26d4fbb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cd499e02f9c1425c61be2d1fd6601a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1341011589d37c7a381db2b89dc5fa8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3bb791adcbd4d938d1a615e98b8068;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd11a10b767f3a1726f8353c99340ce;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h189bba02b48ee4c839676bd6daa0bbf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h143ffb483af77a32e73cd1a24d0c1df;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1111cecbb07b26f7855185f77347c50;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h120c4243bbe25f2945e3ceeffcc3557;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1373ba27b937beda70cec1451f30976;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h198afa91c69a8ba65d366ff483068cd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h175a11302c065145f65aae198d756e7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18a06be8e1060d27fd8c26c87a1c68a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17c62d4220603790b4a0c7f69e1ba6f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h71d547df31c4cb3d2c7c6a66ef21b4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h155acf7e94667f0f18e3dcd4e3dced8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h24431a9b1dc4c65b786610b6fdf498;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haaef95fd533291a2de14ba41d1bd7d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd2e02b1a22fb042e5adb84a7bf99;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h133f5dfb37361a5cc2f4570fc48d36;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h60d6e449405952697613982d38cabc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h47cc948f41693e3dd012fb56db9781;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f6f37775a923c64655d6cf20f738e7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd6f81d459e47d0dccf56704b82b725;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hef88904fd88ac45042ff7e12cc9d96;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14d66cd06e08edbde535f6471242cb3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbb09cb06f0afd7cd9e3d457a41aeb2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h130032f389c9cbb7938dfa72b5d2706;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1857dc12ae7b101eadfc999be9dd620;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h107ba71fc1fb669e786c39cd41176eb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc1e474cf5ca7eddab66ee818ddb34b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hfc3476e4a08dab1b82298e2ab5b248;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a45c01fb74cb9d9fab241afd5d8184;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5b733a0ed665cddc547c875d9516d0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h171af46a44ac376106894a0ed622ebb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf1a6efd1bcf5bfc4f7d97f21d30014;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h95cfb327a528601c17cf0af59a15ea;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19aafbc82726b56a411de68c216bc79;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdb3d61453360a9b979e2259b11ca8e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h182914a389f0ad352b734f20c409cd8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7a4915a185c0d17b3bd64002ebe2e8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc486db2500ed3c95f478778f47627f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15f5b168cf99328929df28354d89073;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6111b87b29a597e0b31e16722073a5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h273e4148730b48604c7992dc467698;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf53814810b7c244015bba08e8e5579;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1756bba973167986085009940de9364;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h533c27d5a4804503355f94cd88a826;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11280b7dba975097f6dca1d962f73f2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h157693c69b3eda1743e1a0f87767ca6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haad4b0a83942fd4440338b1cee1cc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1339fd0aea49adf28290dbdbdb88de4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1eef59c849369428aee7716cedb777d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15a97b0e230a33a085a655856404012;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19a55f0cc4342b4f2cfcf73f6e5d502;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1323a4d831b0f064fe2ff17580db3f5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h91b0ca20fff87ea74cce5e73d7f7f4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f3b34ec605973cdc62cc534500c09e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h178661c0ecc080d6ea7e6bad67d2ab8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b6ee2e0777f70497278edbc57ed987;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3d4a3ecc47c17f02420e985f25e797;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8692d999eb82cd2641a97a5d4ae3a3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb74b4be5b84509f25827d75fd75ae5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fb80c213c3fa8ca66515b741e9d5f5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h197bcbaffdcd6e1ee1c601faa3f7bb6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h72855a91df5ed346d991a6f777cb43;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17f1465432f26772fff8b100ff297a3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h142c3e42d18088447e03cd8b74c64d7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h23a0e8a14b5b0cced52e72e223a503;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10b4bc37be5b3e4076d5f1df1eca5e7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h125f8a598b39c6a6d866ae4dec1c98;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e679472b9c024cc966921d8dcd3712;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14b4d38dffcef8c73b82fab24e219ac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h538ebba287ddde11a5cc7c173b768;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d375ae451e01881b94ba6b5e62531a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h49bc49eff524ca50d3c917cad6f10f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e3686bbaf02145bf3f6362d616472f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h96afeb7e649e7a18850136cba61ea0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdf00041eeec601124f0de5e6c7ca7e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h764c49ad05d316c21ea2ba1d8c36b7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6191c8bbbc8070140f042f311136a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc9f153c699c81a39b43d79c3186426;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15dd749c0027ecefca50b6b0004aeb0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3b5d06fbf2a2c4c183b124cb2b5d70;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf7b0650cabd2835bac86e0c2e9fd38;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he496823165b2a6ad5ef4723a97dd23;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he49f6b18ee07791c7d782898baad21;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h873231d5f42412f3852566b43a2b4b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b330430b910a1c1eb3f860821af4b9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18229e9d8b3494c28e11e7e579b07e7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b9e9aa9eda3f1d79826970296addb5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12dcc4bd795da58a75c94791ede32eb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b2e321536c85bac3b3b16483b51e10;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h146ea00eba0cd65ae147cb1ed16b738;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1cdb4e2946a16ba20e30281c60e5095;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1878680bbd4703424d35f49ce8f5aee;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb1e60856e179e6fd738f44fa600a7f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3f4c0d60c734dcc40cb03eea351710;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13093c82c303d3719c6d7c8909a0d85;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4ff5ac9f87d917fbc8677e3886d424;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd9a4adaf3df82b4d7577199366b5f3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12d705774cdeccf1e9cfaac63e652f6;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h122487e699ca87abf99d471a754e33c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a322267824145453159b79aeef27d2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2a01b8e2e90e89f73db19bec7e3c07;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h91e691a8494179fec50e689416224a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc0e9b36c37a613fd8f301425e59d3c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h192806766b5e9c4aa8c24aded2a7bda;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1dd2b51067a539858332a2fa2b16264;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1212850b9824fd70339f506efb0e3ff;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17c601ff2ce8173325bb4d0574112b0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h106416b1e8702c97b7195650658b96e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8d501dbf988a7456269132d9c89f10;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2284f6f12a674cc41b19580e048bdd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8cdf7e014a357cd3c3acc1b95ea6f4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2192f4eee81a1c401a40ab8d228af5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3489b28884d77bedaf62b227f35a00;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h126f25bea008e0381581bd46069042f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6e7126efafc3dd051feee3e986abf8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3d723af88bb955d08c8e73b915b93e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15f136a74a0e795abb7789414d2c20c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc8674e6b4876e9d1f94f2707a3dd51;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1020a6007634b0df647953bb904164;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1216ca627d2e7c0a18e58cf0747b15f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h93cadb898c73553281c1b597036edf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h157cca249a33aefc686ef93d792669e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd1728f2baefdd7ead81aae6d31961e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h178f37dcc5eecdb3bae54e250aea14f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h159a5725c14afbe00cf03531695a426;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h138d69d8a02e0e6e767c48426a59bfc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h114b7773ae151f13ce08ffe106ef43c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1341e9a656f1da3a190404844cfb15;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13628b375babdbecbbd620b2d3d35a4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1255cdc675a6c7accf492a44c2f1ebc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9d25fc88b7533c316ef41f1cfe093b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1aee09bdae6592a4dc78e45fd950124;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f9156bb54040e8ff794dff7fad31cf;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h142e8af13f1cb8377625929f0a41f0c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7b392d03b8798e5db6d03694770643;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h66985575656102ba0f16df0fd05cdc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1303bf22d6158ce5754dede4b86684c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1fccf2eaa9f2171162f3677494a8cd3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h486ab0beb4d66044ffaa28f2e44b8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha71e0d18b07e8186ac1fa75b36bd22;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haef0de26a054bf83b8ae085eb2686e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h83cdeca52131effe74cc9cf99ea6d8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11c5f61954dbd2999051938a096ee1a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3b5aede53d55b61450c378d95b9d47;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he87ade01ceb8bcf315a56fca166c02;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbbd443dee50263fd2bf7598d030689;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb98e436279cd75d06595bcf8bbd21c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hab114a7cf23a5046308a5c93d29c2d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11426a5ae37f3e8df82b275f9be13cc;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1de02ffd9fb4d40f76cd505ccba3a3f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h5fa8affbda9d63c979982e578776fa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha96633505271f8dfe5e3eb8df9f0c7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ebbe63b486a3433466f78721f7a6a1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haaf2252c48edd1a38dec8364fb44ec;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h54f1a0a1a39a9e558296e101251814;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd68e0b07a61bc46e0348a270fb4633;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4ada59c2c64a5c03589904a7ed072a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcdb4c5f9180380bdaf4edcdb6fb833;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha81d71d69f8473c0f4f54ebb378a38;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f89cd6d6cb686245cd7817988d0a7b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1589a95ccfa23eb5d524bd76ab4858f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c0680060f2afb59b2f62fc42fcfbec;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h575ec459961667d12a4150a058b53d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb9ab4ec090f3f424b9dc90d9b23772;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f4266080eccf1fa925e66b66a7a939;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c4fb83a6a7f7e656e18229c0d83ba0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12d42d185d202e34aab843c3c4a88b2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hde0a6d50eb9be5c4bafd22c532561c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h7cfc2ac2df6b220cca790640451134;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13cb89f60246359541e3ba0ae464b8b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12f9ee39da257b5461abf1e698248fb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb75f193449728d95d5e63046bbe996;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6603a90d3c1702e888f7f5f1bc842f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d97ae485c1b69deb47a654b6b24e44;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1901e8dfd4b95ac1db4505c4c0923ad;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3f5be30584c89ed7bc891f8020eff2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19b3b13f3524cf777dbe8d58e0fee1f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hba83aaa055ca20126dbaa2c940054e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h573f75ad285d8bbaaee50e723ebe18;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f48f61f4fdc85bfb129055c52b4196;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1036fa379af495ec59af66f8c7dbbcb;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a2b72243b5c2abe0fa8203cfa76080;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e15b51baa764a6c857e1998120bc9c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he08b636c72edf09ff27df8a9cd449e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h73fbc3f36e49d96f9bddbb516db3cd;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd703a8a8eaff273d89b623924529d8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h63005be66e0d877acb843611e3c16e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10596e6bcb04abd425a18f8aa91da9b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h160994f35c4fb03f9a44b5b07fcb359;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f837d28058b05e05a7bd42433b808e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4170d36ab648f48db38ab86b2a4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13cf36fa3e8c09a733292081680ed48;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h133a0c02eadd35c90fc77006f94cb17;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h11d769ff326202cafa25b10414b3754;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h170f77b8ae52b5da6aa7397405403b2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hebdeeab2e92610ab4bd564866f45e8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12ca4d23f001ef5d73bc5c0fea36333;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12933019e7c5c42ea45b18d600227a8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdb29d4cfdd877024a7a8e98c10fed3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1d90725fa10e6f0e217f14b78ce2ac4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12566d3fc64b3e66292dfce9650338f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h18fcb926a4b7106a573e7f71a84dd7f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f94b96920e4974abbfee558e631134;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd3885fc4df3a315516b3730be0413c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h151278ed9f32fba8865e97782e54d46;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h133e46a39cc198a1936760fb329ce4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd7f7a83c5a234af553832f416289c5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h110b872b5eff664eb5d05020afa1369;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hbb0723974db22654d03bdbe4152ea7;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2c481729fe05d991b4ccf2d067a64e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h928288b535a5129674ec4c6648f952;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1faea42a942ced0c5ac828f40bed2d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f02ecb5119d78f04b3f54ab5dfa215;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a3be70b2b1f73d80175b3e3e026904;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb163e75af250d7ad586cee4bef022f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h46497c590976e2a45758807deb6b60;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ac9e9a1c15093e65cb56d066e0c85f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h522a88b49f4cddfa95342dcb5d83e8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1edc480953418832c1e799cd654550b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6c6a42541af7d3ee5b7403f55cf4e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h2f8701354a22b2bba0a6d360e8d090;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf13173a1c72698243663f5ecb07b81;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc9ea495c7769aede7dcb5ec0998e39;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hcabe6142bc72680e0ece38a522b95c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h501c4dbdb31c9f16d7195877ff1030;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f3034227227eba37dc2c2053c18d4c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1510b5c83f525ee9dc4117fc0171fc4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h475052eee3653f5ece8e02ed20c4fa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12c45c51df31d8be4029bfe0e49cf09;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he7ff28bb0bb6ed9444f2c420e22c44;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f0b63e331847966f3234aed60afa78;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf159eb730b8871db432381a3865ee5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he64b620cf3984a4e2c250a313561b2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13778b58816060e5cb033361ed557d9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hb79efed5ca5b85c83581fe4fe359a9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd1b3ef2d7177125f6fccfa4d29f613;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10dd79a1ba004ba26373a18e4af36e4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15e2cebba1c0f7329d6216118abe31f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h64b6c2db1e74bcaf191564e4aa3f88;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc9a117c138e906af8d5034de663f6f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdee4786bca15f4da8cfec4efde16ab;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h49b803f2761bb3806fa42d33933780;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h8fafc13756a5ad594218fd71acb16a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha01db334d342fdef4e2b7753f4ee96;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1ba21a11115c758e2233f20fc89ece0;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a22573c18263abeb0f71f6b1d01a42;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1738e2bca4fc040fcc5306197601418;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c49bde1e3d0217cba99c1339ad8b30;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hdbe5c6c0f790cc599e67a76c2cb4b9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h4ce20b778227adc52b0fcd68e2d958;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h36a762870cefc9509470614abdb960;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc4f50b645a76926004bddb5c203701;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19f9fec60f8b2d0d4405e620e6040f2;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b9ef5c8745ceb657733b7786d8b130;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19ca67c2425c0814142fa166910b8b5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h291b81e14cca3ac718fa96808a99d8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'haf15f9e724205d8b82a1f81fc00f8d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha137834a784f3a6deec5401e68c0a4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6b7e9281eb35ec693f11de86611d8f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h61cb41044adc2ff34c0c5776bcc479;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'ha3b97e04e2d4432b7e8f0e962b6309;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h9af642b7a56ad5562035e3f66378b4;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h17c5d31a04281aae2144500063042d9;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h658598273c99f268d47593c72b1991;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h85375a18058ad0064871fa90366620;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a79238c893c3a5c0dd1d7d58d8c186;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1be32be6f8569dd364a35e0783835af;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd409198020e310c885fa342456038b;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1722642d1e4fbca8a51dca077564b53;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1843197d2647a494309344a45404412;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hc7c667fe792702b6903523b17c7ba5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h187abc28867ac76f47a1c19f7c81420;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1588c22351b0e16cb2770771e03d34d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h6737b850386977ffe5c5b62a24f050;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10660cc8b2fd14bf08bdbcd0e184071;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h19ee9c83660ba3182e5e2637218e5ee;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1599cdd7af15fbbc05cad2d6d4ca66e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1e2779294546aa94b24750a1851b77d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1b5ec0717b661099d37924679cd490d;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h927f45dc0ca87b56cfac1e48877e1a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h3681e9f1f1e4ba0195370ff940d126;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1197079174bfceb5ba47c90885cd334;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h405a955acca6f3572f21f0eebda540;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h13ebec9b558f282349e6c1b606b79e3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c95e2b774adba81737468c41cb516a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hff0df25c2abf88abfabf53191d8273;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1a1dd430e9a06c55f761b95c236d8ac;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h161f8d73c23becf07c47cee881b78d3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14f0f46427cf1cc83c971d243de7bba;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h30138f5b8e3c2e84d9bf3c373633e1;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h565645b42fa23c4c971b97699c300a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1bd64ccb3f890ca352e82c6038a56fa;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h15160a7918da2d2bdfc427b8139d26e;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'he4262d611f0a5210fa805215c39fc3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hee9ead227841137a9870122ac92992;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hd916d36ecdac365f8b709889b58259;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14f210b5943346183e5c819dd709f7f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f887632eb2386ccf99b31549c9214c;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h182f22bf0b3e90795b8e2ae66438b02;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h808ec49ed228ab2eedfff15779dfa3;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h10b43d512227dc1ffe27fe18faf2a24;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'hf6143ae213be0c6e15066a7f24563a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h12135d1a3f841899963c511238e01e5;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1f4c193cb16abe7aaaa539bbcf3595f;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h14c32524547fb2136042ff5540f4c0a;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1443c9a5143c9758c3d3fe1920ca519;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h124b0f0db89a40a14772dcaff366c63;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h111a44ccd8035e892a23f3984d90bd8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1c7ed88f0a4d5bcf81fa795ee95d5f8;
        #1
        {src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 121'h1040496991631ca949cef60e489b097;
        #1
        $finish();
    end
endmodule
