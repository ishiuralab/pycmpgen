module testbench();
    reg [13:0] src0;
    reg [13:0] src1;
    reg [13:0] src2;
    reg [13:0] src3;
    reg [13:0] src4;
    reg [13:0] src5;
    reg [13:0] src6;
    reg [13:0] src7;
    reg [13:0] src8;
    reg [13:0] src9;
    reg [13:0] src10;
    reg [13:0] src11;
    reg [13:0] src12;
    reg [13:0] src13;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [17:0] srcsum;
    wire [17:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d1d4c578ed5de1c0d1e55ee9a0f6b083390589b4d1bbcd56;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h382802bd87432ff2982a94bdd996072ffb5c75f9c89ba2f7a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h253110ab549e65a92f3119898991becd31c79ab9e320e9aad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19420ffb2dcc90495f8c37bdd9279e9e4db91216b7d014c8d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hca6c77c3df28462bb2df20c8ce8ddeda355b2afddc094a878;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa10ec367180034863aa5fd805b763e5dd633475c62d6311f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae7cc899c3981557c5a218bfffdffb5a54e2fef6a4d9b1063;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d3bf1cc3e7972af493e5932a47ad7ba94b1b9c3f57fb73fd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8dc2b5532e3b0f93f5fb9bd02c33b8a967f8675d90528397;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h568b3987c85094bb3491d823f85545d58ac88f0df8d098156;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee98d99ee983b6f2240037cdca3593388d0fcc629847593ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62d7b2b7ba0dc2646b31e95a7ff640155e551d25f1ef90d1d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h730e0c6d8709f1f8fbe5bca605dc7ec50fe0feb6ce9e5b284;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he540c48ae62fe79a2e27eef270e62ee25ed42f3b50ca889c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f63b20426627a16fdca1ec217a44787cf6e3da5867dce847;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8393f4f612f6b473aaa87af7d8d084a74b190ad342285c5c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7eff9c0c84413fa660098e8a46040136ae8e0b0293d45e24;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e9bcffde7c4aef9f45c53179163fec6964c7dc298691a1a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6fa2d1e9ccf330ac0f79caea55491fca0f892e6953aebc7f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h38019a70806ddbc4a87e599945bb0becac6be7df94f1a573d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e62d6210aeb647f7ff7b7320ea3687bb02fa600583412fd3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea1abbda7079d9f8f7718b23d25914b01528a00c44e8c8789;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e828472731645aaf32b8070590debe6eb7e8c8b9b977db37;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d569ca105c9211f92a36a2a1ad27bdba2cc6ec061fec08c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h792708070a9db1c4373724940234e8df7ebc0fd761dc288cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd63bec007590500a1710137b7acd19830c0f6098f5e4e98bd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd37d8839181a0a5db20477039ee0bf8af16285378d6dddd8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h82e6ec8be00f5530ff13131c21d1cbdec85a2ddf213e604c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6a7d7abed9da8700bf3f4c0f527711f3cc0e11a41e02c496;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12592abefab0c005f9940a5241a25728cd95f16e2f078c8d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7185a64dfafe06f89a8b8d2e88fa37fcd6b44ea163a1190b2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c5afa3b2bde3b3658423ad7392909e3a0dbd7b7805da15e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf9dcfe4d5ebdb8e3641dca546d5eb1b99e07f02553d54598;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46a4610815d62c9a0b29bcf44d8d13429531e856a689b226a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdfd462208428f1d28168e3081cfbfdc96ced46aa7b72af8db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f6b20faa7cb6431e42896811668447e5c4e6cd96fd72fbbe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e2d9ddda57b6a0f6540aa336c1b12af7cc7db3b88264efaa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h500f5795b74d8afd8ca2f899ca2a44a7cd81fb7aaf8531435;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26827908a60d0f6df6130986ae755348efbb0570ffb6d7609;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h897fc856c87f7b546ce6324ed0ed8d7d8664ce3f84771211d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a9b7070fdd0d581edfafb8ae1323f9b8ca1b2bfbe08f53fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29f7b13d43508cd6d1687048bf3a3b8d148903f3a0ff46e31;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h823223fc531210a6aa62e6caa493a404c3a9b5b6a3d64ad29;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbad0de586f5ad4f0c232fdbd0e8070ddfa886aa7f15ab1186;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f1a51b21a1a96cdd53057046d5391501be9021ae14e69995;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heed35d410d045f863c0b469350ac7711d1feeab283ba0e57e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50c9c620f0c8c2a436d9035f110c8dcca8a6734115096f156;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1bb82a44674c2eeff53d96442391a0bec814440fbd70945c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53a3eafedbe4d8ee1cfd9c1dd1a3a2a9f4861d7d1bc647920;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5eb092cecdd0660a928de30ae3dfb129101ba03424aeed41;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h372a117e287fd10dc5a197d7311e19708b6a94fa774f9414b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he1d95c102c8dcfc3649f21dfdaa2a82efb4147d4e5aa7a799;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb107896171db7299bb047b11ac7c68dbfb1a8571c29f8c0a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96ede661352891e149e760e0145d116bab10a6ab1a63a49e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h188b1d91caab61c4489d61c3f10438d205fd8d9c4c2086d07;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6aad6208fbff380e4dbe9b2734bc8956aadd3c7155943a33;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab0450caf8afa761f6be920a7f6c9160d4b39cd4c8da7d011;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h990d7b77c6c5312dfbd5902e34d0039f64df6d75df1198be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd7518f1db17e8c5ea8ff8fc9b1b900c3a87d7013e2ca40e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h574d2eae6bc394e1a906f92c66bfd1050b85019536f108212;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb9d0518d5360c97bc693115cae6ee41fa731ef0c581ca59b3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2886b839ebb60a6c245c5389efb08633b540e880b10eaf8d5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c0d179cd25b46ff8b0844dd84927ba740fd6adaf337c7d5a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d20acf172fd8184fc2ef229f90e2f16bc7c939b22e1870be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0e8e0cc7be7acafbf259d40aca0d7232904bbe3ded90ba69;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2606f607e434cb3238f1c688cdc38ea5e790cbedb6ba9b858;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f16003d1d42acd1c5c8b51b8b05ea89ac8e3636424a957d9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h825b0106f890d57708753ba9a2bf65f4dcac15866b090bead;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h91fe11676b28458e1e60ec940470bafaa0c835b7f7234ac73;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he40922c0cbe63ab8457c2b47217134636420ac380ef997bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f58eda0f0670cd549ff8ff48d89251c9e9ba947ea090d1e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd46695aca0d5057690b61e98ea0f68c2e048c744b013e225b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a8107e182f09fbf7ccef9443a73e73bd705d7e83fb653330;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdde68e4c69a2b27f3d48e31928803191dbae7c1902c992b49;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e289858e30c4080325d36cdef97df7bf7b54bdc690c83605;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8449f03a1e0d2bedea51cd742d83ea303fc96a59789962de;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha4c1cc062ad4565231e509442bed4836457cccf5f96c98020;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdead2f49a04ef82f1b3a292f271fcc161971bc199534f60c0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9e6535b5d0cd01ad79b5e26bd5ce335b1c854f616efe8698;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8850e6fd4ce46e40753bf255627c6023dd6396061f3a74e89;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h392985d50d4887cc8a8f1f8a5adb6ffd01a4d20ea2629db4c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb280e59495b1e7118e8fd796d030f86bd16e6068dadb24abb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34f42909d14198154f63200ed26cde4715be1d3636af0e2ae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcaa4f73265f37e89dce905910453c15cec428c9b345e8f33;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b628ecfbefebb201f4344afa3e6079369cd94c1f30df42e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde5daa3367bd15573d5133480bf02ce53f62f735cd1ce5fa7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb98bced6eb991e3a6492a84ac534067af94f7db1e0b0a339d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3c51275ba292b7af803769075572fbbfca51cd1239009d55;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68174925694186b4ea22edfabc1081eac7fbd895ef13d442;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f9abc1f176890709ea0a1d00e4257170b00c1db2347a79bd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6b5962889d2d76ee557af9f1afdf54a58f6183c1c3ce39a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e14b1eafa4d0a6e5eaeda56ae7c1f0373ebfaa6a70efc0b8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70289e501a45abe3e53991d73edd01185b586d28d133abda;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had1a3e9c43c8e39a9071eda76e67d807d54fcc31123f497d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hddee194f4f7f0887a4874d28d2373fdbc244817053a446af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ce04bb45e143e2bf8666f476b42a47f48d37cc7da37aef59;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba4314e9ec38f8abb7963c2aecbe43da4201e5d20814cb179;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75804914b0f532e43bae9f37bee334082b24739a50ef244ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12c57e9f291d7d41bbaa053ca2f5babc60829baae24ee4117;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0fa3e3707cade94dccdbe03d608cf4f6cd06045d78035a1e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h349e64822d5a1c17c834b271ce9f8d09d5d743b5d1e8aa3e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3103eea26eafce6619495097109a3ec83cd72b78466c5222d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3472f8badd56f1bdad0622c516b508356cc9c7539d261e11;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3056880b2bc706f3f4296c9adce843dcd021f7a818359aa82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc34c3357b98a921862e52ebccfcbc00d3dbd063b56b7bbc0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7134092a9659a73f177d24654c301778aabfde2f57cf5f063;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d2d99141d3109a2359c6c05c6af4c61a5300a8c0fc889d2c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b7e9cf642849cfe08d25e738f51db39427d73430a9e2ad7a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9909f97d860a18fc66fa0b32ff4b5cae44704710eae1746f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c08debe3ecc87e43ec972e279621ea4a0d2f0aee215c92a8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41fea1e0562d6c7d7d98ad3de30cdba0f552cfa5a2e75d142;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a3f80c0f97ab6a6596c5aab78dc530e48f78d5d58f385366;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d9c41155a5fd6aba727e63aa15d03490dfef907462297462;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34947e06c99e847c57233a17a40cea24fc31220339b40d0ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf38a0342d8c90dac0744dd64e8bf50c1c138ddfcf98ba020;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86b8de29e77f939d2158fe3bb776bc209436e28e3a5171924;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h15821f4a6923f25e6129e2254eabfc2cf6f83790d46915fc4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb231a20a921e02badbccb1085cf227979ce6aad8dd1435dad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ab2a2cfbeddbaf09c306e7da174041cbaed304c026c382f2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed7945d7a5a4a5bb39d40fd6eea28045ae77ae519a4dab6f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a0e482f4594bd863f38e140fcb6c559b6b18f0c5921fa754;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h918d97c915d6be4e27a844f49295eb50db6b7886d7acc1fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h544c2a8edd3107da9b78d151c5f7fea7c571b7a413193cf6f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h289cbdaccf1bb969d683212cde602dce0f5ec935379c889c0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1057dc68d9fb38f8188d2b2a2c2d50f364ffbf03aed34435a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72459545be6e92ce2c35fc72536ac6bb4b30eb163b2f0e3fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18c51b71303bad301fc63eaffaf2ba1b8359e1502648a0c66;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h364a07d61e6a3141eb62c44263471906748db468424db4a7e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd122e05c555d319cc168642e0e19b186c02069c948faa539;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52bb6ee386bcd7626bc8ecbd997c056199633805a7c88f0dd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86d16c0c380cce773c45fdfcf9a4510d25d8b816b34142064;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb789a35931cf877b680e80abc7abe9959a0415be63350db3c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4297b8060b59bc010769ec4a15b3fcf65b781bd4dba928feb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc487ab8af6b14d64a606ace053cdffa9737385cbf4532dd98;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfefce7d20449a5b05e54a02c66b635cf4017874ea5a6ec2ae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd385281fdcf428638417a2ac00c1b8f8cdb6f9764e0ff128;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6af961b92cb35dd769fa0070f02bb2dc1d0ad9a1e7ab86acc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb65372622607d9f636b4b5e457fce043c5654a9586a616301;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h85c51ef77d0d26026e44924baaf677b637cacb38952dba9fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42bd3a9c1be7aff37e78d6f909fd06be0480076b7cfc5f03;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2bcaad19b846fbfc00dcbfa53bc353cbadfbac62a51484a2a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h97bfbfddfa9f0582b7c615f612be15151ad2ee7ea5d5e9d9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd849071ca1f59ffefa619b37c5b0ef6a3eedd7ec0b19ef47c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e04f7be9ed2d8c72082564e8d9aef3422d6ea392c87ee80a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h363c50ae8008e06518847c8f5d0a80766aa5f7104e3b85602;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13822349fd4eb6b57f8cbf4df59ae88293070b580ee95c32d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35983ae9e427312ff0f251d1a5213b443328056fb314760de;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b6c67bbb44c5d0b835ada63c6861afac0ab1ae7037efe036;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50e49b1bd1a9c212012843d208d1bb082041a3314eafeae62;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78c52d3185b31f6b9894c98d75c3a85b45bfdd6d0d69174d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3fef6a9db8b475c86af71102e8a0bc4761e2d3736cb7aae4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8cca7dee292937c0168be03cffcbc54c926c2973c39ceb26;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef6e07a84f91e5bc27a495d7ce0d3de0e9717f66adc2273d1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6cd4c5a2cdf670e7134f00bb31808226a5236405220d9de3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f61ea48c3cfec8dd6f64b7d53447ea3422a112096f35b07a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h995ace3d84713e7d39f6fe9551c4199fc6e6de2966b8e7525;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a6a1dcfc222f7707e0c4c719c374c5b642e6b05c8eae43fa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c16448106720f974ab758f50fff01e5cdca91d8bec29fc4b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd502ccb4d748c33d67a97cf407ced56dbcfb4cac6d01c289a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60cf8ebe0212431633ffc07f1526eb61d751ebf5f4b95cd3d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98e4a7986e8cee9a8613ecf5941e0d067c2a9b9eac7ae13f3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56844ad44eb424f6dcc0e412b924813d70ec473de16bc03fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha621868eeb3344d6f543924a6bbdcc43f01f50cd32130e3e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24c6e3bf54843bfcb7b3efda3b7b9ae75dcaaf94f5f6b7b86;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96cc804b371144cf3ac224de2a013a7a2785f5e779d1f4aa3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ece7545f76191178291aeac6b0338c4bb557b4f2e3f522c0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19dc2178ee8c7bc625a10fc96e37c346dec2394042b12e946;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7cc80a67c91d927d94379d06c5dd47261d3e4d0dd3027b388;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1953e0133b1d8fae3a68c5af7b8a3f55753975c8f20fd4f42;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51f011ac24795cdd8817033cdba219e09b4a0bc4d492a61c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he705023e2289c9c00cddb2d7058fa85faaa9bcf22566157b6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7b73eecd60831e2d13f758458d45be274ba7eb89e7333be8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb08221d9391beddea45d0bb4e78f05679c9e4c89f7e55bd1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e4bd66680da541cd3de3b7086a15f466c261f17dbe746ef5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16201988fc3708957cd21034b15adea55eb8796542b7ab632;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7080990ad3bac110fa2b0514f4b3425b267fcbef9c4e6982b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he45f3e2396c111ed045c78f4ccbe7af532b455f6be2264371;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha370d6a2fd808291c48f0e0e10c37d1cc862b2bfc88563f3c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73fa0a9e8748c579c491f076720c0abf6c9d26af49ec81302;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4177309ba5490f750804a56377079ca2b07c3f252d2921c41;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20f96dd2682e9f99c4ac2fb51a3163b024fe9c7d28ea553b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h621eeb984637d7ab8c9741bfd0b585dd5cec452e1ec9be5b5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4874a776d83a0d07c3d21b4c3d224917d960bf9270e5e890;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8477924ec83b4751feb5e4d9886e1be77254cf69472562ea5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6e963bcf0ca98517891999ae5a52f030928e0796b26233e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10f3ff933f85a65dcbc2e00ad7b670cf81eff183888802990;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f8d60f99a4fa69ab5557d998a0c063e97e5c74242c3b02fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8952c5ac181a8eff2f49d2584fbea35f3a3a56148e934797e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h81ecf8bea61dd18e4315ecb28b4594dc38bb5fcac294672a8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7784f4632534205b0e248a6fc7c241728a250681bb9012726;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4c8545182b23b1d1d34e8778cf2f899542d911fd2f090a12;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcfaca9ecaceac515e8e8127b9ca1595537db594066040db4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hafc595e01a5f4467220fc216d73552b10ce89522bb8d21b8f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h894f871b9266f4b320c305e08fdca0f515001104b949143d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7596717826132f40ee88b7e8e3780df60a9fb36f341ae6220;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a74b2a5ac39eeb931068694a83ca04d54a75a77dacfd2609;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e4b469c58daa22e8ea414aa6060e8ec0d2e72a6fef71e83c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f3bbb384256db25b73834d7c0180bf4d7a2a37d23938c957;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37c6f9334429976ded9d266784691510c60c0e9d6cc50cfc3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6d423f10ffa75fd8cad028cab6e6fb37afb5999eab7e3776;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1810c7673bed98a28a6d30fb46732b575311a352b3aa73c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1c8fa380db19a1a1746c69bc867de36da928f2f3004defbb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8390e2cea878c451017142eb54fa0fa2b2c0c05213011131a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93dc611068462a9f6bca12568c5a5e3d53b64570fefdfc837;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd45f65bb0d575dc0530f1c3a1f42c92c2d047983c9b583acf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2693b80244eb49ffec4ba1563b6712cd23d621540f23d9203;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a2153d46d8cc9d44b14b5175d85956019c7405c52622a28f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb239b04d44180c44fa6a39f3761d3ecde1214eca1109ff6e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5ac0efabd60d6217070349efb94a8994abcc2545112123af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h677134ecf99a84fb3cbb3b61984cedf81870715bf7566320a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f886c30e7bdec4f47c03ef62e8593dfc7103d7b42df7f68;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf6725c925cdfe3c17012ead39523e59447cee7cc3fbc3676;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h925a31f714c50d795a1cb84a3f2951eb31392fdcae1d52c8a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8390aed5df54dfef4b9ea3ab4925eaa9ee8d0580106b455a6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd535f467984e078d86712e24150c9656873dbb13c9889671c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29400e15b74331476b15cda230882ede9246472529e4b9da4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93a0b2a3194c9d73048bb73e37fd53c801ec0e34495390041;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc31f7a59cc5509b10bfb5af926eac2725833ed4564bbacee8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87df17621af2c1111570d53d0c05b992733201f48e965de2b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65b9e82a8b96a11ae0514c87c9873aed12728cb4fe3091e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7fddf106d480a10069749d69da42da497787021730903dd79;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbac778b75f268319094afce3f31c40fbb77c1817c72b9ca83;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbad06df033849364db5046f8baea165ba5ec2df7074aa1076;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee00aeae1201ff816662ceae73c6394d195f1f3ca6dd54ba0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b5a696ed59cb2fdb3cd75473073e79cdda565a9316678c3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f031652024bce985428f9cd64277e1ab8617e693850e3d2b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16732b83b23dd3f45e7dd477c0f600defb4087216d02c01c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4122dfea405c63ea0dfe3cf9974b74dc064e346f55729d5b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8788f485cfcc6c33b6acb45f3774332d866f225c33258ef0d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c03767c252f220c0504d90bd394a7db868f1b272ca34a614;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had7f9cd575a859db0c0f699286fd7523d6ff6d432c021e977;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heaa4b800f5e2f4b9d2316dbcc5beb4fb6404440f3c7b97fd9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc141a139ffc44ed249aee95bb0eb48133205f1c83249b4306;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h266b726227b603e412edd70689a5ca654fb4ec54df0d6d6eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6d2df75bb7ba3bab58086bfea6d1cd7576627cd59211a113;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1497392fd5a7812d8826e618868d91bb63fd2e4751e1a6841;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb69cade9e6a0f01b92e79f60e86b4d3554ac7792fc431e513;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf353cb0198e52ad7cc5163ab150735b3997080802934bea3e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9494999a8bc8ed95d4c9b01fc8f83488a3508bb22031742c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5d2778978cd36e86a7ed163631ca5e054be169d7a10d00b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1f3c94487e7a15876a56fd92c495c302fee0e2e379f1b9d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h349b41bd5f3956cf13cf837caa0f4b92d55d786b3e55171ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c2401ff4fc695c162248ff85aa3d83cf2074ab8cf8229458;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb71f4a5f025fd265e6849af6549cc60831361b88d425bf68e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f1c530816412b46ea16dccd939ee13aa175f03c287664f4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e7975b2578af1a5357e0e2cd6206e33ca005d2149056ccc0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde99e8ee5b543632cc4163a689f686ddc461137cc0c5234f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42f82296714b6dbce36b54c653cc48f96548798c2c1cee97f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67d6e1edd9ae13fa307134a0236915396d0b7908cd8738f12;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26bf8cbdbda1128c24f8fb9740b93b196616b2084bcc979d4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d02db19c9a72ceace5b208451e412b8d7ea386f39a0dc519;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e6ad6a82017d987aaa173b53fbf89c316c84587298fd8b25;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4e3bc42804654cfe789fd76339e28921b7d149c99fbfafae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbab7879aa8b6ff32f16c94baa8c44caabc963d2d99aaa6767;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a64db2af19cce63276ea1e9cad9fb381360fd5264f683c17;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha4aa8389863dc8f0d1a9b3adc912f3cff7e350a36e8d52caa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5265b4d57dbe95b3a4182539c6834142daf2064ea3ac4dbd4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2acc89687227e60ad1e1699b53d09ea9cacf2be60e2f758e5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34766033a26d05b3db15349174d97a8fc389c9c5bd114e3e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d8693caba34222e72cf98b75add8fa2e92e8cdc7055aa6af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf03333a4d92665169d6719690b8410ae746fa339066e9793e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4b4dc0f42efc2572df762b4feffbe30c0d80f4564dd66154;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e1ace9f494fd457c1f7758c6611cf7b908f46b70a3ca9432;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ad1c510a46f0b22fd2ef168cab358cf3d25feac37fef6c69;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6389d795763bb625d2b13a0fba139bb2bbd8817c649b8bba8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16a9d9c7ed402d23604726440b3c79a2affb3ead6aef2ff42;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha90e59a7551c5ac75e65de3b78eaaa0ef092435dfd0f047f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7327b114f0d576d3c5fab558a3fa7e93e38896b04dd99c862;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d49034cab0b27a890f2dae563c8bf36bb4e7439714e9c514;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae2b85072c32a4ba0389e9e3f0355621e8dd9a11a1e34567f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd73f6c0ac00efc1c49295965af2f4b17dd2a74cbca0468d46;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4aec4bc065c8b7e705bf3923b48773d72c8ea06b04aba73d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd31cac9404fe19684bccea1c1fb96ce83645982a3f2eed13;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ef6de019b5b4e77777a756156e651feff6bbb25f21c4fcb5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hacce722f3278e3d7746a4957256c6cd24095458cc9c1c47eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h428c92ec302585682e8639796a3fd7a2ae9d9d703f5fc8df8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heded7d0645461ae3d0972c316db7d30ca9a6c51ff1aa24e1f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h64ab1d8dc25330b9a9d8eef9b1bc2b22c91ba6fa8b0722ac8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf102af28809a20cf805803dea18caca2856f9bafde133dc8b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbbc441270465a4c229a47162772722b8a0e8e807c5de0eac8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d1d9b995ddef87ba44f34725aa14a8eac48cd46050b30d36;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5511ad9f0c1fe2d786628a901247dfc4ede17f48ad2a4505;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd435550c2a91a4b8c2cc6461707109f60dbb60586658c2cb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8980844908897b62253978861b0a68605252e36689203d322;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb76f1d26808aaf5b9cfda6685dce9123f75e8db093211ad3d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1dea185a47fd3303782da8f6bb3152f5076e14b06215ae44a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88e29832e40c18d4ce8e1a56c8021916a8b808c0a96af38db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d82cb10ba58b0d95ecd6b92683430bc6f9d020f6aac6c959;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff576593bc2226685156304c17e149eccd0c8234d0a9b63fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he961561ab4e09f2d111ae5f927058560e0ae944620735fce5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4b4a051dc884238b999cbe92aa42449630515905844b2a8c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb972a7cff33c43f262490897af97a95e3559cbe31fae34667;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd74045252fda2f884b5a53a95d87d9ddf4bfbc439a37383f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb3d09e2850eea1f71fd8f72335309e72976fb9f059b154358;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd7e00a65db6303afa1db567ff8956ddb6f758899a02df5dc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hacf42504280cf354eecaba31bce4f0bb3d90a34199d1474c8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93646c8d646feedef975d7260446ab3b5b5df1d8441065f7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2f29bbd74a01e947383e5622c696272afcc62cdee98c69b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d1d5a287e89eef7f42da218edeafdd864bddafb6f742f269;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13dc27836315621de930c1036c8ca31a296d7f996c779a6bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7150d97e8801f3e3fc377226499e5c2f3928361e8887dfda5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he92af0e196ae065fba320423080e247200b201b2e8419861a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc01754f9d2a071bf96a1400357361dd6e8a44fa5f8e9da5b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8569f72dc8a4fec2bdf9555dc16b88a0225b99098252e4ce9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5fc200784e2391e9599f453c45d4a9fc4f5fdc0fe275b48bd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdef62c1b9f8ef48fbad00d364ab7f834a3771eb5347a18418;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d41c998bf0a0dcfdbe3b6b4e856248c9aed47a798ff1e8fa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d4fc376eb4762d3defbb830918937e297b3d982b8990ca51;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65dbf21703231f49115e4dfcaa3e1b56eeea8499fe162c85b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfbb1760e8d263288c8eda9274ae573af2fcff5b929e2b61e6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2cbc0d04198fd12bd18069f7f5e745c3a96beb9e346bdfd2a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53af7a966623f73994c49d716f2e242b62cdae6d38c9fefc4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h439a2d32e4dd1f9d27a29a08d4e87dbe09449b2ff54d85e27;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ba5b3ac5b047ca7a02639dda2994f9c2f1f3467d6a25f806;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfef96b863058ae6a57bb384ca08999f04eb57a25469af64dd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a61954a189322a0047df231a4ae2f3ef62da9bcb20198341;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f9b93c903b07629e1992dd0a61505d52f087a7acb67779f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6fc1bf5c0334144fd74bab758ba64e6c5515e6db18f64ccbf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3cb49f982bf9d8b789bbcdc68345107eca1af0efc61b9ea76;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h566a6f661607c181271f347124b8a0f8dfa5b149b95432b25;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52722cfbe4f54d622421345f9246663f74fd074e98037ba5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d1c94481071816441e4d1055fa2cee3543035eb7baf73c3a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ce211505c1a2b5feffa9da26b8f4941228ff03d23034d445;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb920a0713bb2d215a2caeaf8b10cae464e899989edb85a11b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c589de15c33c2361f6b428c2b450f32f844c94b9c247cc63;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11c8560f76045e5ff87fc9506364695649c213d4604e72b47;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d20449362f972b8d5f38f1fd21fbe102d86ee3e8d27fbc2a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf31b8fc8f63476d3b43baa2bb82a57db3256ab9086b13e23;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hecfe7d959b1dbff001d2c8c13c919993770dbb4501143e133;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff6154f4bc4dc23e7595c91ad93bbcdb707ffd852696709c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc114e86e8aa7bd6f13ad64b4175acb03ad1621588c5f31e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3154886ff925c028b5184aa9146c94a3edde0d90da8944ff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hffbacfe28d6eeccf6e1eb2c10bf31a83d15ae7d20a1489316;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5d9930ff57f125844ec109c7c030827c7a15335a0f28b5cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba09b9e8aaf1d1962b180dba93df48e47a438eb3838ffec6a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd6d1834c93a45fc48eb5892d20d22616971979fa3faac8a8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfdba874135a84db0c6da678da38968fde0615144d32c9fd6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h342eeeb4eaee7bb36e919b7a192f973f03bfbc9d278746a1a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78c32272bf6fe0fb988582b27d53c857ed9e96228e674b248;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3cb6b31860943a28619c708afd45bc9dc5c747ed23613d8d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d70aa076110eb7289880dcee5daf5cddf7025d7abd3e4c2a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd114627672b69305b5cc39d657e444bd92415e0e200209bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41a1d37afff00d4ad0955882ca54c3d5e09b7f32492044c6e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1c3e9273caedf07f23a798a94e5700267b5e02aa97ef708f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h675d52ed1544d3ba98e256fba1fea3d33674bc768582ae087;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e109f009623def785383e41a0aad2cd61ef182cb0aa7fe3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde602f3502526ae56719f93e5235d51db432f3f2bcd5df2b8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbd1404dca1569847cf88f966160ae57d431f672c2df52891;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22103fc3ace32fc24226f67b89b7b919def1d0406ac4c984;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h531e50f1f38b5c3382079c73c244d99c1a272ebcde0b2ecab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed7429a0ef230d2bbf30d76023029903f81cd82b304f28d7c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5283ff3515edef6e69bafccf8f7e0b8ced8a09e1fa1c0a5b5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35b1b613647f235cc3a95644b6939990a47cd0008eab312a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74acef23bfb36a92cb0409f404c89293555a6b36198de3145;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ab16a124c6daf73c9695b578d86481e92c16c3d63cdd628f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h116ac5f82576dea2f4f1dcc09d52e90db910c27b4e10d078b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5dad64192a1ab254d5bc5d66968dec6b9effaa25efee42b93;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95e937f450d7cf10ad6e830dc0d4e09ac0801ec12a9f2adab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcfa1975c937ac362c1ca5c40e1c19609d37cf93fc41a9a4ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3e01643f2da4843fc3a2f40e3d46da252fe7b90ecfbbd41c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21e078fd7650fac8193a164a854ace37d5da70e48faddd65f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47ddaffd1e742d6c8ed867085e2e5055878a5f873a71c02b3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22b020820bcda3c5591d7a87e06e93c2da8dd0a2b7d4c84a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7014c49df1faa921233aba7608199aa7672613815cf9e04f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff24693eb5bb007f7097fd94abda6eb95471b94b034dd6674;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32ca842b9e526241834501674d2d7bea9ff1b49cae6a7a5f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8719b08878c8524735495c8163eb894271cd152c2a080f196;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71f0bcc83a10d897f2fce7a70539ee6fcf16c3ba01ae52eec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he2508562ec43651c29ae408f4c47e0e89f2728ae5bfaa7e89;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6262f8ffd2c610550cbe62323f91887bbced64b807aa59b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62b8a87e2499fa8fe40a6cb1ef1f3e25a50d43c88bfbd5f3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf57805a984cebe2a9baaee8df8ebd446e0434075824ad3c8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had2d91bc20ed564e6943ebf3191d03a9c3e220065d48efa63;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9430a898543bc1e9547c245a0c05764a97bbf5db11c47831c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h278b06d1495309d2a120eb149cad3fa66fd8a7296f566362f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c8236d94bdc8bf32926826c92d13f2510bae2e38d7a53284;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcea59f35d0c49011cb00506b38f661fbb143a8533c01e35b9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h736302dd0985e34afe33d95bd6f648cbe5e36d045d68ff254;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6638b37ecec2bff00fbf169232ae81fe5c9379c1815cda76;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd491972c140f3b481bc507703bc29f2da6fb1ac260b3ced94;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf19995edb74185dc35dc689311b93c609d070ead13025f7d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c8ad44f582b4ae963e22639f435554f40512849f94849c58;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2978be295013254bc88bed9d605fe7946fdd9d646d594d02f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf5f447dd8e2243c7d5adc6e0a56c22094f40614e474de18f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5f154f3c7e8d23feb2f18c84b05c3511c3eb6fa2d9b3b062;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9000040bc2aebf94f01e409a7522fbe2cc17686cbaf20990d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b8a5df7f74e85fecd815ba440044538765941862cd154181;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d788129fe2ad4c18ae2b5190ed05f482416361bb36cb3ca1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6be4d52067ea9bbe271a935fdb55610f5fdfd15f0e6ca82ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5fbb03a14fba46e078ed47f596f5db03d9b869c1a32bb51a3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcbeb9c6cdf574e3ccb19cab7de2b2d22f02efcc8404b8e7e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ce5908437f2a8dba9b1cd063dc8072207fc01c57387c71bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd866cc11fe76b72d8d49bc919c89af70999da875128da9f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h576e830cabaa657acbc2646decceea1679f7f2f1136b47445;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0a2faf4bdd69da7c96ef9ca3ae42e82c0249fb46b1ebff15;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd67bd825165a1c39a5aa5c0ae8991bf2b5ce4e37356d1a8a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18ff699fa355a8fb6062854945ccd6d57bd348684105d9aad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec8520f956c871aa6348b77eb28630369ed27b842d2aebec4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d2991a067eb334030bd0e66bda62f60f398b19cd10728f23;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he27e97538c3f0fdf5abcbf38754ac74fc032a72dbbb576f80;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d409b28d86636f14845db011ad16622e782b2f31fab0fb82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea989e48de8d0b55c89bb9c557a3db91b190041961d32fddd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ff8a60e861bab7c8f20c92a8bf792d284b7fd08160b4924c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h149302b9636806072ae97f4f1b428d2b8b3bfd4bb82baa264;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79082b7edccba7f93961ba0ec24c433fdda7ca5d9b3478d83;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f2606c560d94907017803c3b99c448c1f75d764fb02caf24;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb8c9298e61d48d25a234fc2df674cba5b42b5d765f8ceb70;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c87a6c9cada6db5646af77e0308cc7fdae797840c88062c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h15c96324310bb15308ca9023c2f4c43b83f4a52d983309083;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h85b3bd3bf9b705c726e527727e00a0b1c258c19c7c696b592;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbace81adba8b5e1f53ed8ad713695914d9cc7a59a606e003c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f8e9bc4004232eb87b2352b326dfd0f0f84f02c5ac1892f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h492839a72da58597bcc53650902979a2407ae348994b76461;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6c7e6db3247235a348fcf7f512e43bda1fefea24417927a4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h39c1a8f7db70406d4b1c1617976851bb9fe2dab5fe00eda9a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f42262673eff6658f7e7c900d4bef21ea1ac7d9efed4c25e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ed858ac00c3ff5d14342c0b843e6532c93ca3486fd9f6e2f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h925b1c840f2c5d59bc44ce7df884b8abd14a85a06cfd578c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84a6fdbc577e966df8b7c3816aa62dd4f0d0063df21f1da73;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd362b98f0c465f7ec0c201e33a065eaed7e50de08caf265bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f171789f80979dcb61b41472015ef90e7ec5d76906fcc9df;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had1866fb5347d98380c906a4077b23e7f3f747c6257d3a4bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed2bdeddb89072ce4dff640fa7c1b3827ec69672041051670;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40ac9b424896d637ea946a0535d46db2c509c67ae0e91fec3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d44d23ff7f68cbdbcf508dae88bb5927c4431ff874c8074a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6ed8b628b00737a05b52f98cb55ac98a529f002f0aa49009;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba9ea577653b0d06a520314074d3321c30d413f47fac407f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfbc3acb8bdfed64ba541e8ca922e41bcbb872439816c129d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4791be841599724f509b809dd7053282fdd1113d0110330c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5fcc6a136e64664d1b3a96e24b61856d6a2e78dcb744cf4cf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c54a3953da73208a880a2231e09e4cb3d91b2d08c6807d65;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1555fc26b8355cad4707739404941c3576fed06d674609b50;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d9391d820089f70891fbd54d14783a65a7080cc3fd248f10;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hefdb7506e388bda8dc59e97ff92e3896d3eb57f181652e0ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c956b8de5a63005bd66543e53b5b00ddaec6eada9a4af22b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h704f507de368a397e76df884a8ff194ec4e01c95db9d6f587;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4e79260041592ae5bb5de56a33dd3f64a6df3fc06fffa80c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34d9443147602e5b10e12c1cd50d490c0960cbc2f66d933c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae579ef8622d0cf335f1470399eceda0093ffe6028685f9fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb24f46859f594d7b977d0ccdc29961194959d945f45d30926;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf33f3953feabb421965ac9fda671a9ca4d360bec90c578230;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcb033f9e18871f4600081da7aea96be1d302806df999eb3cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc41629fe7f4667dc03ff6498b5ab7f6b546c9e91453422426;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2adb3e60a5369f9eb2816456b4ca9fdb537931ebe7acdcc7f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2cdf79f796ad515829941479a8000e9cee20bbe6a45e91f34;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hafc35755a182a61901c5573951c5177f091b35e6fbd3ba67a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f5675921fd046e14c560a22f549b387c8f62e52a0b04bf9e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5293bb252afad3b3008139eb8abb3e683d49d867b73dfced4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77626e555d22bd43a65220915a8495a895ed8e7babcfc3bff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26c0219ffe769d89c09711f1d5724905664b40408dfd6c6f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc9a0736981b7cf35254a81a72d2a156a85578cbb5f52290d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf65f89c492a0e11d18d50ecd8edfaa42c56a10d30784c60db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd820de53b429322788331aa51dc7584f6acce3c9ce09b6ba0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4c930589b0bb131278af50a75c953ca01377a6b4e85bbfd9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1e7e19cad8ca44d3d38d6e9309b423f50961c48de03d180a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hca8943f6db3744f69dfafa36093f100ad41aca1df654737e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbcdb5f9c074395ddb0a50b754d0a15db6e61335d99bad66de;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4fe7ff6b544adac21aa9881f2befee14bc9d4357ccee9e6ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb190e8f842fce313f56ff44cd4e8b0ea1da111447baf953ab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb8d50680a77e63aabfb2595f1f6e4ab80eb036f875e3aad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h64608876cacfe32754ba08527bce207bb09d338986f7b8414;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8e739b74d81fc86e2d3deaf6c7c1fb1d3c81f725be564979;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27ab9b8ba5f530bfac38cf370955f055e10d06d6c15f860d6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h161e17820701b26fb7bc64ad9c2eaf52444d66cc4dac5e839;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35d424d02552d8d64d3998498c1d8c921b94a4fe48072cf80;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28c6d44a99a28efda9d9fd0c8c33bad5b407e39d2ea390a73;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf7c16856e1114d5e625db707633d9a5bb4feace242611ef2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef03785dfaa20c0720bd96920fd1ec210dedcc8d39c0057e6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13ee9d7e2c5d2c4c1dc09fed70d067c5872f91b646825877f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4cc490497d4e7cef897ca3b4c0430c46e45a8b3b4dd65224;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb678c52084b4dffd1c01f700a26fde20d7bf19c0d3491ad6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4cc708554ea06ddecb24bea0ca0a4d798722dbccb0fd35357;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96cd69a88a838d6dc657f464eafe53cf049340872cbecc295;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26331f5ca20ef3313f77bfcc9439c17aca71b5f6789c935a6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7203be5863207721f094e1221f07df431f17a06dcfcdc259;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d6446e2e6b3640223eb9ec8a77f36908b9679275633abab0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h398494af891fa0027c38c4df35deb32b7af3f512050bcbf8c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h442906bca45f2b4d0d4ab60714a4df758ba53c25af7b9969e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3db49f7933daf26ec3df9086223f7ab4c221ca4054d4d4fd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe47ed98e549ed86ea38df8f0762a2492d47bd686eda111a6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hccd4a07c5c3b516dee28b1fba544bd283c0609f624fbfedaa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h23221b4e0d4f7ec1e89d261807fa79912791cf89e0e9f7246;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd19947f16bf42b5084a20b62c59e7787d9a49db499514044f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9652c4c9e6b62789286a58dc67d88be21dc0ae5aa0e6330be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c7fbfcdc39281688fb8207f5d9ef1b1ce427e438737e782;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45a11694aa48ad5d77f3aab470a7523e0e6434ab917b22df1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3c69b4312888a3f92863014e9d753aafe043e1a006965bd4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcadd00291e3209f55c6502cc8d642ac2509d4d3311cdaafd5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e6774dca10c69aac5b39ca4e53d71da5f5843305f1772cfb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hafc1714bb87878a59447f1bcc6d18a23486c2210346a2a6b5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34cdb919d05cb4c17a5d8e30a35b190fbaee2bd1e82f4afcd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2af53aaa2dfc07aa123bbd098902f49235f7ad74b33432f75;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he0cb2b1d4e312d0fdda826c7418c72986c34d02a0c9fc1c50;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h659ad1c7298cec8053cb1d3a1af4f0b62a9539b4de943834;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe3bbca21d09571d8297c61994544d393259d0d5c3c63b64a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hddcab0c7f1b2ff512954f0cbc5a8a2a2b6a3132cc06ecb13a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9396e51d2278e1c03c50d0e7ba57fb264fe93a4fe3a5e285;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d0359efa8aa7edb21fd9eb9e83fe0234b237abce54d5c0bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf83eba7338e5cc08ee219a5a6cb5d1f7cce20f2c29aa49c53;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52405f032d26110ba30bee985ca2c4fbc96ad6b0268ba3731;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3529e379a91fbd5d7aac4a53a23d93e547ad46f644eb85cc1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35d6e56045b1f677c5d28e5cf5b3b640d89473275836423d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbea7e5e5fc00f7a073ccb4f3b64c276be3a2fb22a4a1936a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17f722527392ab133ae660adec164a7b36be9adae49559b77;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf574bb010c697e938e4aeca294474bc8c5b620ac0eeb5a0ac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hea84639d40da0fda373fd628eddb7c720f29c53bd349eac0f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35bbddfbf074f1822df02fbd20ca998e0a04dfa5ae595a909;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf96a63a7c6295e033ac8a0b216f77af6304f0fd50d4a9d4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha671d5eb01f6863303bcbe5e49fb79f26c7ca742119b589f9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd95ee1728cf74da5a00e442f08ed8651519b51060493a45e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5cf6db3a4b6265f567da69b40557a71035f3148b28cf91f4f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7af05c18e6edab944091a54b2364a76bbf8a10d6490444bb6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he551b11b211826ec5d85f964fd40e8b5f0be4aaf49a509aa3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c83f81a8b7a87ca63f8f41ec861ee819e2b8c5330afa6565;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc79dcc397aba8953886433405c6df064d884637f7bd50302;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44feffbae01b24dfb6d351455e961062b68aaf919c4c1a1f3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e3d0db24248cc482a2f22a2a3daf0833eb98d520586518c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1a17d302e8cb19abe320e6d179ad463d803d7d956a4d93fa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42af5bf7f96a737debed3cfd78989c74aae7fdc00473ba63f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53a540ce94e09e64c86703f0a096d402c4d10af9cf4a4829c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef605831716789e7c7c303c1d730aa0b96d47fbedf11abf9d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33200c35bf49ff4ab31e51233b82779fee247b17a17fb446d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4781fe05d3c45c8a1767b6dba5f08fcb66fb9b61dad6c69d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc0e2ce1602562d48094246dcd137664fe3bd33ade9007eab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6016adb9490bd41b79e09823c05949d4676a794655e557eb8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f1a7609b919b7231168bef4a23a6c997edc9980348700e98;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79cab8cc549707ae8abb4b5c2b629144a0307395fe783418f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heaa1cfe32b8ee966a273c0335dccad19ead39edf5376803;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2722b61f610f3077d774cd7c5510d40190c6dbe5fdab646f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hffd66dc2edaa35517fcfa1f6b9210aca8cac6049b58230b78;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b4fe0e4c13c4d6c0e41992595d06816a501ce979499d9f20;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52776d3b5a94c0ffbec714d3b3b59477b364286d61e435670;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c6286b4310fffbe4a568c16beabb6c4f7752832aa2276c92;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d9f6b3d923959551e38011128fb4e2902ba22bf6e26765c1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heeb2a9cf89e3028d2a47caa8484e02182b0ca5bff65ebd181;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89b08d613e040444a17e5033b985e9d4ad094f8b27d8d9e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f6ceab82ed78d0b7cc58e07bba85580e55924e12a627d679;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0a1de06436214d4d2e4713d8e43f7eaa34a41099b5a65355;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b8bf798466b1c140ea32ce9774daf18f932e79671d1fe9bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h105fd72975e61f2e3d145665330a228419d79df1b19a7722a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf5cac552d175f9f5b599d5425e11f1c9acb24881f958ca49;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f1fba50406b3ad25a1bdc82483fee1e9adc6b59fddf9b41c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3cf4493fa12af44ce3ddf923032c606d1ef18e4825b8f5990;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9963259b337250be755b2caed113af9cdbad57b66cab504be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7c1461fa4b3b673908f776de3ecece899e6aa4f4ee83c5d5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5261c690cceb9fa3a04698d4046d9f4120d2fc708cad892ab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc5312a8fda3a03ac80f9455158b7f4184490f4c8029a6e1bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h414c47bf07b1f4e1566d159c4f74836e8bfb007dfe4dc6ad9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a081a8384701bba9ff3d5d16763175f9bc25d5e0c1b2c322;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h801959ad280e064e49570c1440ffcc5d5603a610fa823ce4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h732650aec4325ff5561cf4714c8a760a73c694b9c1b519033;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5b1ad31325021cc2be357fdf02023901d62090e377358981;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5affd3bdb78de4b2a2d67e87d42bfea950945b3f9e2cbc870;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h768f91a42213b713248499b1cb623e304e01cbf5a7b522980;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3404bfff83140ee1815412849e789209168e165671a586815;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d6b842d654b6fdac42adedb8b1a9ba89a1567d21dab075b9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc216e535e21a4a01589af435adcdc31605cfaadef2c2ef4ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd44d1f7833b1664ecaf4dfeb9d3c900254f09929cb36c58d5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha39de623c1a2b1e39b1a200db0b0ebf8156c82d66fd5ea2ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4371f963e40bb0a8663817185cd274909f703cd1b3a2a8d85;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c179c5b104f0518691193f24c40ad9511808e915db9aaa81;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c751d2a2827110ebc18ad46ff791af408b2b6e66de61ee45;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3bf75a77e441fe85d166731e3141777a1d2446f6d96dbd6c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcce4691a1d8a7a410436ec1577c97b6e272918bf7284bdc6d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b4fb8a3bdf876d13ce6bbe8f97bb20e15fa4efdb6a383e9c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc26e6c9f2dc369a2ae7c393b40921290ec24cf2b72108cc9b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h207f28743ad406330dc88c94c6662917fb54cf839330d5cde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7718a883995205075efb125d01cde5e792e1e3603481576da;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68da1a0d7f443c387591edebc8518b930225f02f53232df56;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed3d36129ec1f9fb315d92712ef4e49e9dc607d48145d88b5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h798ce712365cdb2a330f45cda57c480740703d9641d9c7780;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h824bb475a08dfad6c346b4413eb7b00b7f45455e5ce508525;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99c30f7bd757dcc552bc0daa2c2199c4aaf7907e743c0b982;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd102c03cee1e34da580fe7e4b42de076bf3ce9e98d29b89b5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf43104eacc4a412bf4acaaccb53e339e6e814b17a656443a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3615eac6567752efda0b67d7a41de7d4ea03e81404b560de5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54b8cd3075be3e71077dc94beb84a91a032dd48bfb792866a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45bbf935308fdc154ac994acb5b5bceeed6eeffffdaef613a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd8c4171efb7c00f02b14b61a7da75a9ae1af198067c978ac3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc37c776e4d80acb8c284fbae3c444353129159d723f2bb827;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he729933c9f6078977df4a81c5e3d3388ebd0d574a922409fd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he06384b5c0dca41573e2152735912af9a15c3162ce94836bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda36dec2011f07233bb55760f84711907bb4e94c8392bc3db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7bc39813eac7ad60f3a2d50b27d74a5b847497227703dfd50;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd8022fb915f6b9c7e2a23ece2181c12bc3a6301edc629d8d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8faec1360c17337dbb38c9269ade59d82519b8d1d981ff331;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12126d6d93ea12281f1b1572f26e83866b659090a7acbb182;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfecca0e2c973fd7bb962d14311f28dd7c12b8da54d17d8711;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff441731bbecd5ca102464ab3c538caf98a8720098445e026;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h781f1f33f2eab302b2be516f37f9597057881ed1c3c27717f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71edf0c740b6af30f402c2dc3c4bff3eb765e06c7f5ec3b7a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2ad0209cc31ece96a5d58984d817bb5cb5634740307d7985b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5592837212e3c4da64cecbf2c11c4e547915282a6f689db33;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32ad17cadd37e9b2038bb3fe324795d9a4b113d5a61a24e14;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31b19af524c417fe273a41a2b75e2b18a11a8e731680a7e09;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f027e0618ce176c40d9653a7c5427919ad53e327b009a3d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c78bbe91b3e74dd117f95edb78ab0ff6dd61da4d3914a96d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52ac552207d49fb0c96e824491ab07a5492b2d8b139c6a0a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22af6c679a72de7de2402cdabea32a3c74c0dff4a78fa846c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb70f505b2caa05081ff49fe7952fe1a26ed4fc42e3ab57c24;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef55b3ee0bbeddafa0fca6940830d7620b7faca5280dddafd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2576701ea8b785dd513339cf59a9fbafe9450dec100c1bba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb25bdf4176d69948242a818517f7016deed1b74243a92fde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33168bbc11ca7d909101a834b97b03df717a6afc0479eed78;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53ee1545a8936ced77c1e748705bc233ffb9184e9b72a132e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h97ca04948aa0faf5625fb3c0786ffbf6eff4db0fb60b98e2a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb25f48fb94cc76a2c6ed3c81b65684bde9c11e57039717836;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbdf8ac68650b9d7805234c0bf8e137301e3daae05feabb116;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5248a213968eb4d427be5101e66b40ad73e0ec6be0c17f2ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7a303e4d5ce6e65f33aecbd3f77165d3fca149023fab6b8b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d76b222755b8ccf43b4f95b18fd22de42bb4136529548c73;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9dad75d466bf8cfcf37fbb90c67f44aec43ed5f6855ba8d6d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed5262b7974856f838417338dc8134cc561e2cbb1aa2693ff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59ed13f1829bbfd4e52435f6745bfb180819934a995d13faa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72e1bb58bf6fbf77660712efedd8fe035f9945d6a554bf56d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd3c00756a438cb309f5728996602dcc8ff3ac001e8a91fe6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf29ce7677a0ffe580a0af8f9a2caf853c94cd8bee88ed7e00;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86939ff502bef8f83c3dd4c11fcb950ce37484cc65089701;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf015cd05923992f1a5b4609d8ab17288ac65de919c829e413;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2b4d26f9551dc61136874230a36bcc29e643eda368ab6cf0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc2057fc7c3df6761029ab73bd2b953a9c2df96b6b061b0c7b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4926085180bb4be39e42b8dcc7349732f5059435366f3cd1d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ba399d2ae704e4a7f2ad25b5ec8cdecaaeb218b6eca7f716;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff56705dbf0d74433f6b33d6cf4df753142ca25f217bd932a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h425e07d975bb9ffdd0ab6c4347ae081c2c8549ec8e496ac3c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd74eb50ec6e35b52b509da5049a71260d52b2ee2db3631c8a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d157ee91d6aaa1f9a2a960b52db5bab12eee6bcb94333870;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h580104bbe926fc3190b68234a72ed5981960868c3f2a0dd60;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ab1bdfc19da694bafdc67e2f52b5123fb1c111471418dcc4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87bfb19d518c61db45a98825682fbcb32cc2d620682be855a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ab9c78b01c073eada5f150156d1d5f6f46a01f84fb44619d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d29c9d99d413639155aa32e32d05a049df10300f915ffa9e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha12d4c1e1f4e190fb5f61aa04e359d85fb68272d7e8ee236a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h682ecd06496bff1e3fb0888fbb7448170d7c1cdd8a65ab602;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ecb3ec660cba3c517e4140f3dbc59d6497de04fb5e485f7b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba1d69472b5095661d3226c79877f3ae349527b161e5c2410;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce5959665199331d51a2966f3d6133711cfe338ad989f9315;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec7704954df4561d86623cbd4ded254571a2b8243ddc9e544;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe61123dbb80c9cea030230d3d31ea4fff70c2bfe34aca5cb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5cd17ea5b53ebbaf3e3158e9c788dfe109374ce0c06c6c594;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h78bf476c52101f35fb9c345e61169218fb723edda391982b9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3668ed4557037617908ac80568fe1bbdf4bb7aa2895940bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd14c0683dba63abbdba30883b6f6d3ac2be53981c255a8731;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22acddbd9f95b8a4f37e77b25a207a32bc9e9615854ae04bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd48754800a67e5f4e3b6a3756940205fbd68e80d5540631ac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52f46245a5a7e41133d02ae29c5e0f9f2a510f4872c7af8b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75f66d36139c1e5bb4c980c774b0305a6e498a4f5b5950aec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hded2651ba59d534bc0d33ebed96e67fd9156242fc992b61d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h615834e2b6f7c22bba9988d554cd9cd00deed1e830242b7d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5aaa3279562045dc54e035529e42023dc6404851a6feb506c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf49c3b67435d07e13210fb1859c77c68c761834256f248cdc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha36bb668d2337d21fca8ae91efa7f8628543adecf0c8f1ccf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf50320308738d1c66042a16f18aa73fdadbc20ff9d04192ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9f0b1aca3d368a0083adaa19430adae9877948204bd6e04ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4391c9e271a1d90c934e61fba90399fa847c0f0c141f6943b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he2960d0e4554f3de33cb828b307978bce9dd453b7ba3933cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7891d3890508b7f2f56c206d7155a0823f7a2dca0ac05b2fd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f34eb749e6e7c4562742bbfdc62879246127f5599c7ba62e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h64a37855f16d9c51e784b877396a5ec4a38ec155e4180d9e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h653a9d06f5296391bb4c4d7d756d4cebbf4fe5aee546e5745;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d7c27bf2255c03794fee31440db090dfbec1f490565a246e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he8489c3ad17612011ddbb2fa19904f2c9481ace8bc53c2ce5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a23c7130d9cda67448b31171e4e8af400c5083ebfb087f4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9076b78e52dbda442402c457815ecde533ae88074ef6bcb5c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf6c108764c3be4812287d6057a887cc57ae2bd0e945fade7c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79299565bd5fe4ad651132f8b561612d7c0e8e0cf9de18953;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7983815e623daf2d1005d22a3d74cc25b59ad4be6d0bef8b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hddaf364ef9780090851d4a86d014459f34eecc67c2a48b9ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c67cbac27d1e4871df655e8e05a0b8ee467d7e051e9713b6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he59c2ed79bbae4782bd76618cc6a101cd1e6e62ac47f8ee94;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc19c0da1118ea1abf90ee2c3fab191cec1e5e00f896172e8b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72f01d65d2c979595daa7134dab857709f3aa3574d52c7fe7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8425500a55ad958781a206905de22c1a01881886cc9e2afe0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae016ef3a77814a8ce6435f55b7bec148e5a6f8fbd1f82bc1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6707f26bf582b1cb14306e0ca0b77b6b837781c15f28235ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92bf1d98a2b23ed4b57b17c67582b2d764f2b739403afa4f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc1cb7b063a0ac1d0e3b3613b4dda11d69bceb1e69035d658;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he40163dfeeb2c22652adfcb62839a548fab0d55b62999ed97;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h191096c764e6f5da2eab2df36aebc701b3bedd1cf594b645d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3a6e9b36c8076f6381568c4f3c90f60dc1a20f93cb9a9007;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha18f06b3353851a17bcc562720afda80e9803dada0a9f71b9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbdeed7b16ff27003b3843c0b0c31739881415fa3bdb01a844;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h271270f4567bba325ca2fd3c998715cf05f8021924d50baf6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he1b1ff0de65ca6e786ed50a080537c603b63e0e86e65ce16d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40dfb8a7cf1e12eefc2b5e6b28b621b4f3f3bd1649a0dd9f3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5769991f6cdfd1eb1d9fa3ecb09ae8db5e7085f31af225e47;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3edd4aec3eb2653d686bff7b90bab786c4791a35cbeec40bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h269fba1ae9fd54c4442e894d29569c65d40ce596be398dfc5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb998fea77120342237f0369f5e7c6f58de5ee2c5261656be1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c8a2d0e6ad8cd2104ec6b9c32c9568fe97c2c2de7699b72e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h716705a3ba5da4402dfa46d330f34fc4a5b7117432e9af089;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb636adb1397354403f06032ce3a85325421f4e35426a8f74e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1f96228c8a7f38cb2afb69ae666f6c9953381053fdb94f8d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2204f0fdc95049ee5f0c00324b9cfdb937d62ba945c416cb1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50fc1b632c0a74991773341add0d3f068eaa30924efab10a9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3969254e82b8c216cd6da0930ccb7e19c3caae043a9a2a1f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h707a54512a7fce69f3ff03b449a0db4755bb304c6579e1c85;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b1112bba62bbaa98fe709b6befae9063c7d06c6d21f6f93e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h748e310429834c347197f01306d4db2a48fc66d5839ec7a2d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h336d714a515cb179885aa6b4a39b643ab740fe41cc7cde0ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7119344e6d8d35cb02de14dea587f917370568342db60a1a6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcfff9bbf6ba6e788b9a6b815ba87ab421cb0ebcfbc133ca47;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9080b2d7cb552432215d3e776e03dd47566d79dbe84857ade;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6c359f89c76dc13114a93cc0356bd060224211890d1b674a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69c00f205e87b9c5f80428dde2ab58ba56782ceb1c5e9c983;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62b6832395a11437b456d6c8f8b7fa5d5a05c20a5e27566db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7fb777438a2ac50fc22def564e30d12bb5d609242a46219d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1215e5af426b4d2286547bc6d47c9dd71973518cdf8d5c7dd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5af07c31f2f1e235310f3bf7d56ff17a39faf224961f563f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h330452dea61f94de95cc1285173526c96a251b4ea442652fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ecf126bca3180fb44492ebda682a18d453a9f5d81059e38b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52d70ff441da373e88c58b87136872303125f5f2b057e777d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d6e25fd19900d8a91bec6a48996477d83f783fea671e4d18;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h730c155375ef96c584d0e5385cf0483f71f2c9f1fd882920c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha62e2653c0b5fd7169d3fca0a77030487fd723194b1a109a1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b14539c4901f43f8736294d6c709587675fbd12c5be0c301;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf15347fac0d1fbf58a0eb2b078951fb30da99e0586e20eba1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcdd65d1478d1f0f11e6558fa7acf5e0c884979d9ad8f8f259;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd449721bd1dfcc56fbee129d99706bb1a0c1b7892d316494f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ca543c82bcde9acf8c9cda47993a09ab0b5262a69bc8349e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60dc852d0eda348bf9af7b37e2048a32560835a9fd6c0c52f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha765c598bca61f93cf62f430f5ae69612d289f205bf4fcc6a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h401096bba1538a86f473e021ba5eda309317138a34f684c7d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4fb9eeb57dac962fe1e30385cd0172f37be0b362ea12b431;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h80236c7e06ee484b61d30a1ca7bb7e162d535fe5dc43314c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd115e108515b48e6790e53739b570e4f0b3b0ace45d3e9317;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hffd8c5cf61e58d9ef0de1e089576ac20bade9d874d0f957a1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcfcefb826cd4290435b7d9b70f5de7432925a770c06dc754a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52d48b3967bd99a6416c1e66608f04ffbc283dfc7dc73f690;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31282691791735e5919cef7b0e59649388e93e35254d2a7c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h790207203047b3afa3385c4ec5f6f02c83c46306e66682ead;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h240661998f733df2594a7752fd205ed956ca980a1eb596f9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcee19eb78ca6976bb6bd3939a7be7d36591bbad1d53a0cc3d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6ca81865ee79188d49ec5cbcc1b4a92de0063d1423e32a45;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19d60f218d743641a99e9dc90c158364d1a316b2db47d63e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h803f8e653e42c3f5210850b7692db8f41a10bdccf01dc965b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6980d168da3e42d35210e14ac0261af946dfe31590bcf1b5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed77abb024c78d2fbdbc2c83b531fb31c5d5a91d5a12fa482;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25eb790682018fa73ba2897b98f73f981be28fe886e3ea0c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ecb1d0fef41d404108011ac5799232ed71765a2a453f590f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd2c09de0907ecbb7c3e5d923797cc26317eedf1c09d16fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb27cec94d16f0e7e58794c2d52506463ab1c54fd2730bd16f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'habaff9b0981cf55440baa283bcb5cc94f38c6aef54cb3e5cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha854cb31972403af70c5407643c38ec9b1e0ea796853e5fb1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3de72462860985438402f5844c6a374b1222a852b73c24fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f6b7d0632f67b440f9fc45a46342c07889eea79be08c9a3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6fc1dcf04d248502de3a3238bb5a09893da2f966b42daa109;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8990d3f2e814f674988fb48087841f7148f33c246fddb3913;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e7dad6517231f70095e3602663e0c800b4a444209bfb637;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h83fdc0155f2273af1157d7301d86e476d89e71a0dd3cd3e7d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h506d61678386370c1fb163ee4c4fec49a40735958e4591de;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b01737ec1a4b89fa0696a745b818781154cfd2fd2abaf85f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h177d21985819ee2cb38fbf8815a53b72191566e316f4e0f6b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcea06f462efdb0eeef391e8a423430ab6c5b8bd62d3e79731;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4bb4b1b2fc9604e6d60d262cd7e29e23fd898eb1f0457682a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hefeee76e5fb238da075ae45bbe5cc1453092dcddc2a290c83;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h964e497d7c92d1ae6a2cec6bc5d8f9efb7791f922d2b86b92;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha4fb30c00773520fd71d29854211da47b2df30a95fc99b94;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hca3d5f372074512a1e50474a52f90be6f9ca564d6aee79e55;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdcb0a3bf632762947404294a511801b3c4bdb274604e4d0dc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc2f0cce9831f616d13242b62528b1dc415836a10005e9df38;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0844e34a96346b76e1e98b1c57695a2014c53726ba832f0c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ce5622c4d63822e66e3fab91f70d13eeb044a8c78ab0e1d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8fe3bbaaa11c215646f7165b4bf8e3542bb718ead61f809d6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44ccdba669d172ae4e1ff71728c55bc65a25945bdb2f55eb5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6bc90899eb98ae8c569b4c571422c007cfa87c81b57c35513;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h56020068f94b076d17b3e17dc0f9cc943fc5f43dd1a6f1ca1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf724897ee847f01d6b022f25b608fd174c56104656da88716;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef0b04ac0782514301f9cdcde22f267b572c0758fae08c868;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc319a9fa870795456387572eb1abbe32c5f716068ae1a01a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2799f2d92a8047da12900f35b97c325e614982fe90a4e164;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92a42ac8e55c856c2512fe2aa70e94917bd8c60e7b97908ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc45672852bb4586f9988a26a9315a56ad379dfc0317990ec6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae6b84d6a853835407657443090cf1808610c0ac44769cef8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1e44b8d0dc7cb7d28163164280091fbc56b954ed897da4fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0ce567a65dbc9534736341389b2cb37bb83f600024a24d5f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1cfaaf49e7c7d39c20aec7d55b59a21fcc29c6452054fcb43;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h97f659bb39c42015f788a200e43963dea17fc8b4415a01b22;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24459bf07b2f98cd78a1233863bcb86bfcf10e277afe4b907;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2dc57637058e225b62243a5585d31e6902f9b5f51f461d81f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf56b0ee896227cb454982c3202f05d56c0fb2a59d6cd37cf9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3f7798c8339168bfe1c0fa58b97d2998ad1cfbae4ca561d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60f6ca5995da1bc56980d6c6eff26bd7bfb03e456674d4130;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30500dea90190589956cb40366400fe867be9d34e1dfe4b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17da709302194fe5d1c9e3028e9e9e2d691599094e42bd47c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he90623f8b13a1eb2759d77e7acbb8166765cdb1d941dd1215;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf192f2cff35749119e92ef4bdadd6b10f24052bec1ee1acc1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6458fc59e6237034fd903369482e4422bbd4b25c85ceabdb7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc90b0fded12f561ca2247100ddfbe4cb51bbc5dd3a9f865fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6eba475458d6d5f798308ed483af11903b585e992e80011e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51879d0d5ba5b60f9527d7dfe7adcb95ee3f769591b95663c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h396c78abce979f9fe5833a5b73d6ca602b9e4d8ff2b7bd88c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c71b81e5d13f89dfaf0a9f5ceb7fc6ac444346472d04f084;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'headdb8272a110c717b79846fbd2518134cb458ad8da0f7862;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7a853c14b9eef40d8c1c4bd93fb07638e10d2e669529a2e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c1d654fb40688bf76c0d175b164506848b5ad1430e5144ca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae99af63cde9257c6ca04747078926eb4043d57b6cd990cfe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86fdd6d1ff12d6d16fcd455a3f77238accce6bf5e8ebc866e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f5d29bad8151a046ee0e55c1a940ba104a7aa2763a751274;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9ea4c4b2024b43bdc2295c849878cc19e82fb7ecb046f002f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3f5f2e5d82a115f0b285e98f9207790bf4f6ddbc64680bd9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h81ec5e01cc21a6933977377a44a0f766937831669cc54d0eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3800983f7da2c56c0b14b50509b3798bd4755b68d43cec3a3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h373bf25d5857d9eb62f55d53bcafb2d581c965bb56f0c1ef0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67c13d05f6a0309df7912528651f5b4d7256b49be55e9c4fd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd8fcbc0c851e4858e8fefcb13a0e35f35fe62ce2b98563e20;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h115a2d8927b52f38bc690f379d2eb3137df80ea37d7ae17c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0efb12e1d2ba5d137eafd43b22b1746edfd79a6c22ffa6e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65e7e24050b07cb412e1b956061de7a3c7680055bd076d2f9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5439669e82c15eb6321bee37c5e05d6af7d1ecf4198e3a2e1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd22e1e25bc1d76cc5c71f40d698eef496dc7c15bf163876df;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a1426f2d658007646e3cb7efc987e549e03d9d104f958103;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41a78c457d3de9301f0f252858a454cc6166818148c5a2516;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he05e13734cdb37d9a33e5889c38229d88c9f5ce72feb7a226;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf85e90fc9809997b2fc18d87d75cb3824f538cb5e1fef7e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h62ee0692e41972724769301969c998cf6f996b440c48181bd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h414e6bdae0f785441635c6d73b7cb86e6e7ffc8b775a956b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf706ce63e7982f6d5affbb8bd9da3f54d8c6d886202c8bee4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h232c371de3c5c0bdb8eb769f6bb59431b66aeb2726e0a3875;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb039c657320941008a14709e532f96fadc40c846bbecaeb62;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ac5af91b3a0ac6bc70c7430c38a515b1e26c7837ae58dfc8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee216405fd95e164cd5444f6483bb37c3aa01d48b3d9ed3bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ff8fcd2ec7f98cc2426a35b78cc3229b0e97493f2c915414;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h696727f9f3bcbca79f60ba6c1d69f34f2ea79da5cb5c386e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2be1459ef3f576c2c712a3cfcb72e45d4b7c7646d5e08ce6f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h608d15918b9db45a617b4abdc91a2312e5280b9e9caac5c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h316c821e455aefe9576cd813465745818a85bc7a28100b228;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha240f1ed0d8da4eff7839cb6db3a026f4bca3a06a48360949;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53f72072f5d612ff2172ae9fb199c3238e1979147ed00ee96;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9945792fcc7f73f712c1e6075a29c05dfab618fadf2c344a8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d80d06feefd54bd789aa932c5772305403be5b196512af4b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24bcd004a5f56bc1cddb1374fc7bd296a0da656e072319df8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71449c4e73368f1e3988839b1c22a793afa20735ea11612c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8675ed4e5ebd63347ab0d60fe7f779f5415d22338ea4f5f2c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7307c97339b71fecb997fd8873eea609b846d730e23cef972;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6565c9b820d5bf121405bd5c87ac71fe40cc20892d242b40;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h81044cad224a3e35c31f966a627c57f390852c33af48d84b4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3938cc672748e9d751febf79d918b0572c3bfdd4d254d6dcb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha55424cab66e551235a50cc09ccd97d2cb5ca0d8750832184;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he330178be1ee395f5f32514517892dd6056278cb25cc7be7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb83c100b3caa0ceaff35c1f46f1879e69f834960366278c55;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3de34e3e6266613819cb0bc2367713aec54432701325f243e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14620657f879bc607c028f8fdafabaa9dde4490f081143c45;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f7c9c4772945f06e98f8f8d5fb1116b68ab1b123dd58ca11;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h82c2ea18ccbaa55d2d1c988e2d591a4b67393064816acb4a2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4f08ba03d1ff9ae92d36fc7a77022911924039c3f7a931c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h959948e4fc9b2195b7a01522e18a126d562aa21e8aaa6f28f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c4c375cf7a104816fec754bb64855427416b31eecc0d4d7e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc514fc90ed92e5637c39888fe953509e2ba7575fe90e73a9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60e2873463186e481457cdff7d2f036bd0d3567f1f3a30d39;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc71061cbfbe40c9569d7cb6ab5b17bbc0b4a2f8d77db91aa3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc894b51ceede67de384fb9b1796beb7ca2b88d04bca983e91;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99034f7e8730641f570366e3c595e7ec5785603a4df8feba0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0f1975ea86b22dc8e56c99968e14a2c069143e81107cf8f7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c615acc0b0903834a1acf0806dc159b0d13f437024d61b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h553af9571a30506976971b5a478fb5b12a020985a042f30d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49055c512e9f2a05ec10ed1bbaeea9c2bee308327c2ce8c3a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96341dff9f812cbc752f582760e25b28e2e5913e110de1f5e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3efaec61846aa8521fe7777d2f0f37eebb34b6d037175692d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h79198941359e568514a72f36ef0e3e9809f38e6eb83f9384b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hadbd9e8a96d36858b2d8ea2020826f45e03acb2240e793cb5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6fb15d9ba51e7f95b6892b46caabc54db858530fe99d4761f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe9b54cce2a63681298e4ec2beed3dc74ffa0f21003a8577c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd2307fb96b1539ac07e309d9be6c2d461686e131d9c9a3cc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ac74f57a9fa19eb8dd3978bc610fa8b778f0b83d809d99fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd614cde435eaaf886c0a4e12ef2de7d4dced036c25d41e5b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd593fbc7e517c068d9090cbb4a78944f6e1d274bb085a651a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a600a934a785a7ce872b865f3f2d64bec9eec02af22f4cc0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h173a97a7371a894cdd8d8ef780c9fdbf18aba4923b7c783f2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe2bcf5ae0365a06017c2471ded38dae38b10966fe6f86717;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2b70be06459f8e5c484648386a64247bdd7e894987672a268;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf049951004f3a1a5fcd27bd3e5462113d7b8588166442f777;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb8ab141ccebc34459822c039a225f71030d858b432ddaa4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7fc628db2a155562f53fc182411163ae5ce04befa9cc3aad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51a33de786da930048dc00e3f0d4f581c3125e28a440330c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7d1e49a3faf5ba4295346d0830a5170b3e303f680a7a88d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2e4fc760e40fd353bc8f8f322f0e1266c07866712fe25568;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h53ae840c88a6112ec8b2dc9e42f7509bd43a33345fa65efb2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8cbc23c035c02ca09f5a47db04795d78aa0db643c43cbd1f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfec77da408b695f251024ff214b31c1bef5c8f205ffbab3f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfcc63152fa878c913ced1c14eb32ced68a9ee2a01169ce12f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h730abf8722727a5547247eabc90953e738c1ca3893d9e71df;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ffbcdcb7f30e3a3d864ff688c4b93152fdbe9dbea7f05554;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7aa75c54523749486d51a58da000859ac7f9c36cba7e47237;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3e85d34498b37a21ada333d11ea1c12c95d82fc82d619ffa4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcad936b55778fcb11bace6462e2e63712fda68fb3a679a7ef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31e6b121c56c42e438b6dc68466e40222e46bc8543dc11b27;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hded46ac33c4c2a2df780bea631a27c259e4b1c22ccf11fe04;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd62ed7bd51ee30f752af8ba24fdb0bed42610fb4992cf7fd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86aa6a2fa0704677310f9c546c6c777e831cec683591ccbde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1bb45937d90078401ce1799c7838a0fd06e9a9f91fd2a012a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdca42b9497e03516cccbbc9d118eddbfd9496387f9db429a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71df48d7120d04d86068b46646267e3f97f7d60725f9ffc06;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hefd8b27e23513c8692fded45632c1d9e89d90913ffb54585c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67fa8b2772daa6814c98c20da2ac25c8b11abfa911e9d38cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70133c286a045afed1a59b44303cb2e640255eec47e5a987f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h55006d16ae46f68b90db27de1c1d802fb1ff5ffcd2ad2dff3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ca7e004db628b8f4a36539e375f9bd2b30ca825957222179;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e8e021bd48bc053e0352299239664176cde3cf19dc36671e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ae60c81fa164dbef1ece19cde546273ff79750a353975db3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e132f5694f1eca96fca06a8db9a7671d686a7a2cf72c9942;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h219b95ec8eb19df9062179a71c0a45a0938506a497caa9e47;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6082a747bacee23aa02a3c52e3efc98873f1dc40ee50759a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8d8136902054f678cbeb60b255ac71bbd9f458ed2f89caf3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd7907e8041c15922596b44d919620f8adf367d27c9ef3af6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c98c5642406ca1ff33abc976eeb30c2732bc2c776915d6f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha24e6b6381204f398fa5af0c717a2b63f3a3cdb1e04c58272;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfab31531078325b6e6491f0313e9c069597d1574a221f2ff2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfff0414e7374b7d425b877f89907637c52a732740114060eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha267165536895eb4b9769760665f079f0f9f39c84f7fa7f40;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd15dc87e5046738099697763d46f8748b160e2f255ec4eeeb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3cf0cdd785de5cfa11c1305ebe84f3d8f7842f3e29f80cc7d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92fe2e07b8c4c58de5d69578d5d013788a44985faee3f7b52;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbcc972e3ebca57881116304de61206ce0b1db53e08a888d04;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37970c07e8cd314abfafde0dc1bfaf9d8e794cb365ac4e29b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hccf9948ec021d29e74aa1fd66e190c313c1938ef25b7e6473;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4dff4ef55b7367e5941c3aad30770162653a1daf7291dd993;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35e7433351ffc55ce7783aa987b241ba32963733ad4fbd989;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8122108b56b83760a1086b19c5a31a3e1c8c3f50c9ddbfad2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4953d3971dd78816fd2fdaab49b3cfa64b9bbf102ac423a9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h882c9f9e90bd4f0da99ab3283fcfe5f5fb04874284ff1f58e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b976ded27663f45475d96fa32d9f3bdcf6511b3ab8726960;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20f2f48035b523384b6e2a78b966154496f8ddbe0d1672500;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h72324653401bc1fa9fd7abe7ee24181bd4b66695943d67660;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2aa3ea73063cf19ff2451544fbdfd0fa558d67ad6553ab354;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he92b43b66207459e190f99eea21cec58446d719bdd5017a79;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70baca678841d80b37d3979af593e2e3a461c310befc7c623;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda032e17b68c627329b6e11784c86f9ff0beb65787f9905af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h961db61afe8d5946dabee5b0ecc2190c1df9460faeb70cc35;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8343e196a901762e6db17050003944088f073294977c06b49;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73ff2a6edce58650f6ede217267179f7d8e85954a825981e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4825512604b1880445f0ca9c5016b0a84ab0790b9e2909a16;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84d56663096023b9fb06bef2631c2751100b6c1b5c595ca7c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h958d589ddfb5de2c860885b26aabf644146e6467524d66dc5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b1391f83082ca7fcb6d010889e95306d3a1d788a762c1190;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc94538c3e7ed438483586c6467e285cf2a67d02386a29a006;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6475952a9dfec2ac5a686263897fcd69ece82966896f6216;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbde357a0442315f891690f28285818586b35347aba8eab341;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h373f383a2c5932ce058476ea8c31f7e231d9b2f5aff435890;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hddc01ceedcaa515ab7e572a369f5385280dcd6c1ee945f6f7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h13babdfdefcc5bbbf48cf4d9a513c2c84b18691768137d5b9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h46acee7aae4ae80c0175b0492f005f93d365851f9fab6232a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h91c4680775b343bb92048528711ca879e05aa6546cf8118be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h853ff8aa36438d4c91c646f3a6d67c95333a7d0d98a6e99ee;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b60c1adb2f9d5d29bb1370d2ed1c376dc5ecfba5c069cea5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87d0c5fe6b8adeab0f4ce7e28c7d8cb8c5a3150dd2eb34b49;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9023ac549282091826457e920f11df67348074a35c05359dc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h460a9fae7f5147f0b27f81d4fbedb3e0d1053e01639e1acf1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7af2af5ec3cdc030bbf4bb20349da7fd0085809213750ea78;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he78a6117dcdba752f6ae43bab38802ffa4952990913860f62;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbfa7b07dbdec7c190cf9c020887a51cf4d28017de688b254b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h876421370b2d116a03f5fc8dfd8e5416543aa1114d1f233e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf3143f2e41a371a7d3d2daa481299b2fea8fa15c17dd818a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8aee73a5dbaf11d999782f7e3046f6a54c10315ff316d2855;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb12193ea2afd1fe7d2aa4b7a70daeefef9487de656f8fd124;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7bb0300ead158d9eec9eb772aabb3dde9e7920b7eac9cf01;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4779ae76713a798fe8bab631a88c35a5b8083604e5ad3eef7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb6c761bcbfb38ee1f72b14137cd3da2593da2ef2a79f4f4c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb632bda9a14a9b8e26ff19970defe5b383142981ede170dbc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h703fca93f35019e92b9b9a9c9a6623ffb93d8232457b8bc53;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbcab031d25481c7d8a5475e52de604b6daba4a8e24d02460c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf527fc21397d55c7651e8788eb94d33494f87d24ba2fc732;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b2230c072aeb1002a8cb1078eca780577ac5efa63aa0a5da;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8997a18faa2d77965c01f5b012aac391dedf6895b4cd31fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h596e73689376abed53249f905a1c24de0cd32365d1a059f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec4c81420097159597bdee1e4bc6925c79afae3a9fdcfd3fa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5134ae40d703a617d52b54bdb112df0937b03be9ca2eff91;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hca1c7ea3a6baedb74bd18b75a390a915316b8a0bba9b55a49;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae53d585f74a5f64f42136e9f567834bcc0a5cd8a5ec30c0f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h55d1d310a822294beb1b099aea82c6f094229476911f45657;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h39bbe0cde5406c9c2c96fe8750d28f7e33d7805c0c1937453;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2bbff42e3fd367120c3657d37b3b5f16bcd202cbb76c084d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c4b25e499d67ce419af276ed459257df465f6bba70d33bb0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h932fef3af966c0de9eca7923c3d82ee335bbc6eaa6ee511a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h84384649331eb0cee9cd038728d5c811e487f5a0802ccf364;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h377d5a9a69cf7aa0dac6d2dc9362f0e39bef7f635dffccbf3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h737ec2c3b0cb0ee22889fc7badc2074cef1ede3163d8621df;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ebaa49e50069eb57034f1797cf32fd6a4c8b78b548c17b3c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h624c463bc27392aef819ba68712d30f0bc7999046113d85dc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h963b77d7bd7740895e434cc8c86c7ec21981ef2c04a806e59;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha13b459f90badb20b4750bd052ef33d9248fe7ee70f4d2f82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h12edbed4dfcdf2aa9e0b76359197e4123c90e60f9f67428aa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4289c2a2a8d4a3de20dcd9a9fb28b623ba5c8ccef9a437ee;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41c7a51c90983d7a2d9fb1cf03a530f6df2845f626146c60c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7322ee22cbbaf023415701a086ce3ec298a3f227a9e897c77;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee371b2a4352bc45a92e75e999f74c1dd21cc1ed8cf86efaf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h798b3d787b4205bd8a712ba1ee6fe0a8111dea387c80628a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4ea29cda8b2207507bdfec195b961a6dfed9d60cc5558da7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc57fbdfdc27fe739d486f4c7853a83a1961ace18e52b1f63c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc6604c11addbd0163ea4cfabfe8231eec82dcf5e95d95ad0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf8940e4c477c050e108d50aa91279186bfa1d937bbda5e56;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67fc414d4b799476bff22ca3ebd90fff9cd110be7275965f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h988de925fb396fe736fd77d5121b3f4374a60dbf891423e12;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc798c9e0bc6a3c79d4c827b5857c55550eca20b02b392371;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65f51af2e19ce73a30eec55b3839e1d97000c8c12d26cd160;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h83e28e888d43fde25b1c6574cc5fff45a0473c3a7ed757eb6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2046d6cd4db8fc79434128fbb5bde8818226ca1b8857e540b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6291442e3c970ac017af6685abebe9583e1d76d37fc305c43;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e6437c7162cede629b636a700da7f50f99381583b8deb440;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17e57935e4271bb964a2ea43c79e630bcd015b83b603acd40;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd1b6db58802a997b279a15606d1e6e594c24f7aa9bb98fa6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5f2b6287af09fecb4979e0c3516bb738af4b5dfd463e8b6f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he675c99d97c0461549782ab8d947f898b887a3a8be42b57f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6370d4dfa4c61add15ae7f575748aedf65a5c1502d1e6fd9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18a060574ccd77d6644addcef3832b4f17be9c2114e3e530;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ce8e409b570d613624976e858f21b36ec64d0c77acedf3e4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h81b46279328b4b1583b41fa083f6f9988857af5e6b84629e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he482d3173e6bc2193bde7f91eb61362869ac61ff01d8a310d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ad8960cc958a9bcb0ac42e1c1ead1fd167acc5e50bac57cf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ee29833b7ece5d08526c2dbab2aa520aa28909b68687f89c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b73c0b7d5f41ea2ee24016fb630610cae7d5ab22519688fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26c3a40897b01fadaa585cf80efab769c46f530cadbc86465;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc59ad02145bee5918e2d272372f43e76d2e46b524e83f956;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd4b1f01a073c6b89905312e6b02611b12504d3369c8282;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h958a5d69f9f71856743d2544c12bbcd7ceadd79dda84666fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbde090eeebcf363f591ae892484e4006f2dfd61fbfafa39cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6c7c93e1f2a2bc14547164500e057ecc6c32a45a82be7447;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c8d5c81790133d7736201a4974b7545af490a78085a6a4db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6a5c880ac891996942e7d2e67244c7cc27a967a28bb238f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8669c98313e9a927f66762b18d9e3a31e36ce773445be7a05;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42f4bf32181d33b50cc66377745b1b68316029bb61e3b6603;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47bf5f99da4bef2b2eb587efa8cd48434bdd2c89246aa35e5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74c4107ff0f783f44ed63af8dc84fc29204350773be4e4576;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7284903d7882dc0ebf571dfa2473b0fa7eb57c4702214b20;
        #1
        $finish();
    end
endmodule
