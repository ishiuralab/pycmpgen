module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23);
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    reg [161:0] src12;
    reg [161:0] src13;
    reg [161:0] src14;
    reg [161:0] src15;
    compressor_CLA162_16 compressor_CLA162_16(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23));
    initial begin
        src0 <= 162'h0;
        src1 <= 162'h0;
        src2 <= 162'h0;
        src3 <= 162'h0;
        src4 <= 162'h0;
        src5 <= 162'h0;
        src6 <= 162'h0;
        src7 <= 162'h0;
        src8 <= 162'h0;
        src9 <= 162'h0;
        src10 <= 162'h0;
        src11 <= 162'h0;
        src12 <= 162'h0;
        src13 <= 162'h0;
        src14 <= 162'h0;
        src15 <= 162'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
    end
endmodule
module compressor_CLA162_16(
    input [161:0]src0,
    input [161:0]src1,
    input [161:0]src2,
    input [161:0]src3,
    input [161:0]src4,
    input [161:0]src5,
    input [161:0]src6,
    input [161:0]src7,
    input [161:0]src8,
    input [161:0]src9,
    input [161:0]src10,
    input [161:0]src11,
    input [161:0]src12,
    input [161:0]src13,
    input [161:0]src14,
    input [161:0]src15,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [0:0] comp_out22;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [161:0] src0,
      input wire [161:0] src1,
      input wire [161:0] src2,
      input wire [161:0] src3,
      input wire [161:0] src4,
      input wire [161:0] src5,
      input wire [161:0] src6,
      input wire [161:0] src7,
      input wire [161:0] src8,
      input wire [161:0] src9,
      input wire [161:0] src10,
      input wire [161:0] src11,
      input wire [161:0] src12,
      input wire [161:0] src13,
      input wire [161:0] src14,
      input wire [161:0] src15,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [0:0] dst22);

   wire [161:0] stage0_0;
   wire [161:0] stage0_1;
   wire [161:0] stage0_2;
   wire [161:0] stage0_3;
   wire [161:0] stage0_4;
   wire [161:0] stage0_5;
   wire [161:0] stage0_6;
   wire [161:0] stage0_7;
   wire [161:0] stage0_8;
   wire [161:0] stage0_9;
   wire [161:0] stage0_10;
   wire [161:0] stage0_11;
   wire [161:0] stage0_12;
   wire [161:0] stage0_13;
   wire [161:0] stage0_14;
   wire [161:0] stage0_15;
   wire [32:0] stage1_0;
   wire [47:0] stage1_1;
   wire [63:0] stage1_2;
   wire [91:0] stage1_3;
   wire [74:0] stage1_4;
   wire [70:0] stage1_5;
   wire [59:0] stage1_6;
   wire [53:0] stage1_7;
   wire [89:0] stage1_8;
   wire [82:0] stage1_9;
   wire [60:0] stage1_10;
   wire [57:0] stage1_11;
   wire [72:0] stage1_12;
   wire [77:0] stage1_13;
   wire [77:0] stage1_14;
   wire [53:0] stage1_15;
   wire [48:0] stage1_16;
   wire [27:0] stage1_17;
   wire [10:0] stage2_0;
   wire [29:0] stage2_1;
   wire [15:0] stage2_2;
   wire [36:0] stage2_3;
   wire [29:0] stage2_4;
   wire [29:0] stage2_5;
   wire [29:0] stage2_6;
   wire [38:0] stage2_7;
   wire [29:0] stage2_8;
   wire [51:0] stage2_9;
   wire [25:0] stage2_10;
   wire [28:0] stage2_11;
   wire [33:0] stage2_12;
   wire [26:0] stage2_13;
   wire [29:0] stage2_14;
   wire [50:0] stage2_15;
   wire [17:0] stage2_16;
   wire [34:0] stage2_17;
   wire [8:0] stage2_18;
   wire [0:0] stage2_19;
   wire [6:0] stage3_0;
   wire [4:0] stage3_1;
   wire [18:0] stage3_2;
   wire [13:0] stage3_3;
   wire [14:0] stage3_4;
   wire [11:0] stage3_5;
   wire [10:0] stage3_6;
   wire [13:0] stage3_7;
   wire [16:0] stage3_8;
   wire [19:0] stage3_9;
   wire [14:0] stage3_10;
   wire [12:0] stage3_11;
   wire [15:0] stage3_12;
   wire [15:0] stage3_13;
   wire [9:0] stage3_14;
   wire [17:0] stage3_15;
   wire [14:0] stage3_16;
   wire [10:0] stage3_17;
   wire [10:0] stage3_18;
   wire [7:0] stage3_19;
   wire [0:0] stage3_20;
   wire [6:0] stage4_0;
   wire [4:0] stage4_1;
   wire [10:0] stage4_2;
   wire [5:0] stage4_3;
   wire [4:0] stage4_4;
   wire [3:0] stage4_5;
   wire [6:0] stage4_6;
   wire [7:0] stage4_7;
   wire [6:0] stage4_8;
   wire [6:0] stage4_9;
   wire [9:0] stage4_10;
   wire [11:0] stage4_11;
   wire [6:0] stage4_12;
   wire [5:0] stage4_13;
   wire [7:0] stage4_14;
   wire [5:0] stage4_15;
   wire [5:0] stage4_16;
   wire [9:0] stage4_17;
   wire [3:0] stage4_18;
   wire [4:0] stage4_19;
   wire [3:0] stage4_20;
   wire [0:0] stage4_21;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [5:0] stage5_2;
   wire [1:0] stage5_3;
   wire [6:0] stage5_4;
   wire [4:0] stage5_5;
   wire [2:0] stage5_6;
   wire [1:0] stage5_7;
   wire [2:0] stage5_8;
   wire [4:0] stage5_9;
   wire [3:0] stage5_10;
   wire [3:0] stage5_11;
   wire [5:0] stage5_12;
   wire [3:0] stage5_13;
   wire [4:0] stage5_14;
   wire [2:0] stage5_15;
   wire [1:0] stage5_16;
   wire [5:0] stage5_17;
   wire [5:0] stage5_18;
   wire [5:0] stage5_19;
   wire [3:0] stage5_20;
   wire [0:0] stage5_21;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [1:0] stage6_19;
   wire [1:0] stage6_20;
   wire [1:0] stage6_21;
   wire [0:0] stage6_22;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;
   assign dst20 = stage6_20;
   assign dst21 = stage6_21;
   assign dst22 = stage6_22;

   gpc2135_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4]},
      {stage0_1[0], stage0_1[1], stage0_1[2]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2135_5 gpc1 (
      {stage0_0[5], stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9]},
      {stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc2135_5 gpc2 (
      {stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[6], stage0_1[7], stage0_1[8]},
      {stage0_2[2]},
      {stage0_3[4], stage0_3[5]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc2135_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[3]},
      {stage0_3[6], stage0_3[7]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc2135_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24]},
      {stage0_1[12], stage0_1[13], stage0_1[14]},
      {stage0_2[4]},
      {stage0_3[8], stage0_3[9]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc2135_5 gpc5 (
      {stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[5]},
      {stage0_3[10], stage0_3[11]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc2135_5 gpc6 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[18], stage0_1[19], stage0_1[20]},
      {stage0_2[6]},
      {stage0_3[12], stage0_3[13]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc2135_5 gpc7 (
      {stage0_0[35], stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39]},
      {stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[7]},
      {stage0_3[14], stage0_3[15]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc1163_5 gpc8 (
      {stage0_0[40], stage0_0[41], stage0_0[42]},
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[8]},
      {stage0_3[16]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc1163_5 gpc9 (
      {stage0_0[43], stage0_0[44], stage0_0[45]},
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[9]},
      {stage0_3[17]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc1163_5 gpc10 (
      {stage0_0[46], stage0_0[47], stage0_0[48]},
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[10]},
      {stage0_3[18]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[49], stage0_0[50], stage0_0[51]},
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[11]},
      {stage0_3[19]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[52], stage0_0[53], stage0_0[54]},
      {stage0_1[48], stage0_1[49], stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53]},
      {stage0_2[12]},
      {stage0_3[20]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[55], stage0_0[56], stage0_0[57]},
      {stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59]},
      {stage0_2[13]},
      {stage0_3[21]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[58], stage0_0[59], stage0_0[60], stage0_0[61], stage0_0[62], stage0_0[63]},
      {stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[64], stage0_0[65], stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69]},
      {stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73], stage0_0[74], stage0_0[75]},
      {stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79], stage0_0[80], stage0_0[81]},
      {stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85], stage0_0[86], stage0_0[87]},
      {stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91], stage0_0[92], stage0_0[93]},
      {stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97], stage0_0[98], stage0_0[99]},
      {stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105]},
      {stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110], stage0_0[111]},
      {stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115], stage0_0[116], stage0_0[117]},
      {stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121], stage0_0[122], stage0_0[123]},
      {stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79]},
      {stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[124], stage0_0[125], stage0_0[126], stage0_0[127], stage0_0[128], stage0_0[129]},
      {stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85]},
      {stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[130], stage0_0[131], stage0_0[132], stage0_0[133], stage0_0[134], stage0_0[135]},
      {stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91]},
      {stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[136], stage0_0[137], stage0_0[138], stage0_0[139], stage0_0[140], stage0_0[141]},
      {stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97]},
      {stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[142], stage0_0[143], stage0_0[144], stage0_0[145], stage0_0[146], stage0_0[147]},
      {stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103]},
      {stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[148], stage0_0[149], stage0_0[150], stage0_0[151], stage0_0[152], stage0_0[153]},
      {stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109]},
      {stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_0[154], stage0_0[155], stage0_0[156], stage0_0[157], stage0_0[158], stage0_0[159]},
      {stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115]},
      {stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30],stage1_0[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65]},
      {stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27]},
      {stage1_5[0],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71]},
      {stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33]},
      {stage1_5[1],stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77]},
      {stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37], stage0_3[38], stage0_3[39]},
      {stage1_5[2],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83]},
      {stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45]},
      {stage1_5[3],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89]},
      {stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51]},
      {stage1_5[4],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc606_5 gpc36 (
      {stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95]},
      {stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56], stage0_3[57]},
      {stage1_5[5],stage1_4[36],stage1_3[36],stage1_2[36],stage1_1[36]}
   );
   gpc606_5 gpc37 (
      {stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101]},
      {stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61], stage0_3[62], stage0_3[63]},
      {stage1_5[6],stage1_4[37],stage1_3[37],stage1_2[37],stage1_1[37]}
   );
   gpc606_5 gpc38 (
      {stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107]},
      {stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67], stage0_3[68], stage0_3[69]},
      {stage1_5[7],stage1_4[38],stage1_3[38],stage1_2[38],stage1_1[38]}
   );
   gpc606_5 gpc39 (
      {stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113]},
      {stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75]},
      {stage1_5[8],stage1_4[39],stage1_3[39],stage1_2[39],stage1_1[39]}
   );
   gpc606_5 gpc40 (
      {stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119]},
      {stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81]},
      {stage1_5[9],stage1_4[40],stage1_3[40],stage1_2[40],stage1_1[40]}
   );
   gpc606_5 gpc41 (
      {stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125]},
      {stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86], stage0_3[87]},
      {stage1_5[10],stage1_4[41],stage1_3[41],stage1_2[41],stage1_1[41]}
   );
   gpc606_5 gpc42 (
      {stage0_1[126], stage0_1[127], stage0_1[128], stage0_1[129], stage0_1[130], stage0_1[131]},
      {stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91], stage0_3[92], stage0_3[93]},
      {stage1_5[11],stage1_4[42],stage1_3[42],stage1_2[42],stage1_1[42]}
   );
   gpc606_5 gpc43 (
      {stage0_1[132], stage0_1[133], stage0_1[134], stage0_1[135], stage0_1[136], stage0_1[137]},
      {stage0_3[94], stage0_3[95], stage0_3[96], stage0_3[97], stage0_3[98], stage0_3[99]},
      {stage1_5[12],stage1_4[43],stage1_3[43],stage1_2[43],stage1_1[43]}
   );
   gpc606_5 gpc44 (
      {stage0_1[138], stage0_1[139], stage0_1[140], stage0_1[141], stage0_1[142], stage0_1[143]},
      {stage0_3[100], stage0_3[101], stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105]},
      {stage1_5[13],stage1_4[44],stage1_3[44],stage1_2[44],stage1_1[44]}
   );
   gpc606_5 gpc45 (
      {stage0_1[144], stage0_1[145], stage0_1[146], stage0_1[147], stage0_1[148], stage0_1[149]},
      {stage0_3[106], stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111]},
      {stage1_5[14],stage1_4[45],stage1_3[45],stage1_2[45],stage1_1[45]}
   );
   gpc606_5 gpc46 (
      {stage0_1[150], stage0_1[151], stage0_1[152], stage0_1[153], stage0_1[154], stage0_1[155]},
      {stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116], stage0_3[117]},
      {stage1_5[15],stage1_4[46],stage1_3[46],stage1_2[46],stage1_1[46]}
   );
   gpc606_5 gpc47 (
      {stage0_1[156], stage0_1[157], stage0_1[158], stage0_1[159], stage0_1[160], stage0_1[161]},
      {stage0_3[118], stage0_3[119], stage0_3[120], stage0_3[121], stage0_3[122], stage0_3[123]},
      {stage1_5[16],stage1_4[47],stage1_3[47],stage1_2[47],stage1_1[47]}
   );
   gpc606_5 gpc48 (
      {stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120], stage0_2[121]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[17],stage1_4[48],stage1_3[48],stage1_2[48]}
   );
   gpc606_5 gpc49 (
      {stage0_2[122], stage0_2[123], stage0_2[124], stage0_2[125], stage0_2[126], stage0_2[127]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[18],stage1_4[49],stage1_3[49],stage1_2[49]}
   );
   gpc606_5 gpc50 (
      {stage0_2[128], stage0_2[129], stage0_2[130], stage0_2[131], stage0_2[132], stage0_2[133]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[19],stage1_4[50],stage1_3[50],stage1_2[50]}
   );
   gpc606_5 gpc51 (
      {stage0_2[134], stage0_2[135], stage0_2[136], stage0_2[137], stage0_2[138], stage0_2[139]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[20],stage1_4[51],stage1_3[51],stage1_2[51]}
   );
   gpc606_5 gpc52 (
      {stage0_2[140], stage0_2[141], stage0_2[142], stage0_2[143], stage0_2[144], stage0_2[145]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[21],stage1_4[52],stage1_3[52],stage1_2[52]}
   );
   gpc606_5 gpc53 (
      {stage0_2[146], stage0_2[147], stage0_2[148], stage0_2[149], stage0_2[150], stage0_2[151]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[22],stage1_4[53],stage1_3[53],stage1_2[53]}
   );
   gpc606_5 gpc54 (
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[0],stage1_6[6],stage1_5[23],stage1_4[54]}
   );
   gpc606_5 gpc55 (
      {stage0_4[42], stage0_4[43], stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[1],stage1_6[7],stage1_5[24],stage1_4[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[48], stage0_4[49], stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[2],stage1_6[8],stage1_5[25],stage1_4[56]}
   );
   gpc606_5 gpc57 (
      {stage0_4[54], stage0_4[55], stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[3],stage1_6[9],stage1_5[26],stage1_4[57]}
   );
   gpc606_5 gpc58 (
      {stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[4],stage1_6[10],stage1_5[27],stage1_4[58]}
   );
   gpc606_5 gpc59 (
      {stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[5],stage1_6[11],stage1_5[28],stage1_4[59]}
   );
   gpc606_5 gpc60 (
      {stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[6],stage1_6[12],stage1_5[29],stage1_4[60]}
   );
   gpc606_5 gpc61 (
      {stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[7],stage1_6[13],stage1_5[30],stage1_4[61]}
   );
   gpc606_5 gpc62 (
      {stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[8],stage1_6[14],stage1_5[31],stage1_4[62]}
   );
   gpc606_5 gpc63 (
      {stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[9],stage1_6[15],stage1_5[32],stage1_4[63]}
   );
   gpc606_5 gpc64 (
      {stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[10],stage1_6[16],stage1_5[33],stage1_4[64]}
   );
   gpc606_5 gpc65 (
      {stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[11],stage1_6[17],stage1_5[34],stage1_4[65]}
   );
   gpc606_5 gpc66 (
      {stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113]},
      {stage0_6[72], stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77]},
      {stage1_8[12],stage1_7[12],stage1_6[18],stage1_5[35],stage1_4[66]}
   );
   gpc606_5 gpc67 (
      {stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119]},
      {stage0_6[78], stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83]},
      {stage1_8[13],stage1_7[13],stage1_6[19],stage1_5[36],stage1_4[67]}
   );
   gpc606_5 gpc68 (
      {stage0_4[120], stage0_4[121], stage0_4[122], stage0_4[123], stage0_4[124], stage0_4[125]},
      {stage0_6[84], stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89]},
      {stage1_8[14],stage1_7[14],stage1_6[20],stage1_5[37],stage1_4[68]}
   );
   gpc606_5 gpc69 (
      {stage0_4[126], stage0_4[127], stage0_4[128], stage0_4[129], stage0_4[130], stage0_4[131]},
      {stage0_6[90], stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95]},
      {stage1_8[15],stage1_7[15],stage1_6[21],stage1_5[38],stage1_4[69]}
   );
   gpc606_5 gpc70 (
      {stage0_4[132], stage0_4[133], stage0_4[134], stage0_4[135], stage0_4[136], stage0_4[137]},
      {stage0_6[96], stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101]},
      {stage1_8[16],stage1_7[16],stage1_6[22],stage1_5[39],stage1_4[70]}
   );
   gpc606_5 gpc71 (
      {stage0_4[138], stage0_4[139], stage0_4[140], stage0_4[141], stage0_4[142], stage0_4[143]},
      {stage0_6[102], stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107]},
      {stage1_8[17],stage1_7[17],stage1_6[23],stage1_5[40],stage1_4[71]}
   );
   gpc606_5 gpc72 (
      {stage0_4[144], stage0_4[145], stage0_4[146], stage0_4[147], stage0_4[148], stage0_4[149]},
      {stage0_6[108], stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage1_8[18],stage1_7[18],stage1_6[24],stage1_5[41],stage1_4[72]}
   );
   gpc606_5 gpc73 (
      {stage0_4[150], stage0_4[151], stage0_4[152], stage0_4[153], stage0_4[154], stage0_4[155]},
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118], stage0_6[119]},
      {stage1_8[19],stage1_7[19],stage1_6[25],stage1_5[42],stage1_4[73]}
   );
   gpc606_5 gpc74 (
      {stage0_4[156], stage0_4[157], stage0_4[158], stage0_4[159], stage0_4[160], stage0_4[161]},
      {stage0_6[120], stage0_6[121], stage0_6[122], stage0_6[123], stage0_6[124], stage0_6[125]},
      {stage1_8[20],stage1_7[20],stage1_6[26],stage1_5[43],stage1_4[74]}
   );
   gpc606_5 gpc75 (
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[21],stage1_7[21],stage1_6[27],stage1_5[44]}
   );
   gpc606_5 gpc76 (
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[22],stage1_7[22],stage1_6[28],stage1_5[45]}
   );
   gpc606_5 gpc77 (
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[23],stage1_7[23],stage1_6[29],stage1_5[46]}
   );
   gpc606_5 gpc78 (
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[24],stage1_7[24],stage1_6[30],stage1_5[47]}
   );
   gpc606_5 gpc79 (
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[25],stage1_7[25],stage1_6[31],stage1_5[48]}
   );
   gpc606_5 gpc80 (
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[26],stage1_7[26],stage1_6[32],stage1_5[49]}
   );
   gpc606_5 gpc81 (
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[27],stage1_7[27],stage1_6[33],stage1_5[50]}
   );
   gpc606_5 gpc82 (
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[28],stage1_7[28],stage1_6[34],stage1_5[51]}
   );
   gpc606_5 gpc83 (
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[29],stage1_7[29],stage1_6[35],stage1_5[52]}
   );
   gpc606_5 gpc84 (
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[30],stage1_7[30],stage1_6[36],stage1_5[53]}
   );
   gpc606_5 gpc85 (
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[31],stage1_7[31],stage1_6[37],stage1_5[54]}
   );
   gpc606_5 gpc86 (
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[32],stage1_7[32],stage1_6[38],stage1_5[55]}
   );
   gpc606_5 gpc87 (
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[33],stage1_7[33],stage1_6[39],stage1_5[56]}
   );
   gpc606_5 gpc88 (
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[34],stage1_7[34],stage1_6[40],stage1_5[57]}
   );
   gpc606_5 gpc89 (
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage0_7[84], stage0_7[85], stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89]},
      {stage1_9[14],stage1_8[35],stage1_7[35],stage1_6[41],stage1_5[58]}
   );
   gpc606_5 gpc90 (
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage0_7[90], stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage1_9[15],stage1_8[36],stage1_7[36],stage1_6[42],stage1_5[59]}
   );
   gpc606_5 gpc91 (
      {stage0_5[96], stage0_5[97], stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101]},
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101]},
      {stage1_9[16],stage1_8[37],stage1_7[37],stage1_6[43],stage1_5[60]}
   );
   gpc606_5 gpc92 (
      {stage0_5[102], stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_7[102], stage0_7[103], stage0_7[104], stage0_7[105], stage0_7[106], stage0_7[107]},
      {stage1_9[17],stage1_8[38],stage1_7[38],stage1_6[44],stage1_5[61]}
   );
   gpc606_5 gpc93 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113]},
      {stage0_7[108], stage0_7[109], stage0_7[110], stage0_7[111], stage0_7[112], stage0_7[113]},
      {stage1_9[18],stage1_8[39],stage1_7[39],stage1_6[45],stage1_5[62]}
   );
   gpc606_5 gpc94 (
      {stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117], stage0_5[118], stage0_5[119]},
      {stage0_7[114], stage0_7[115], stage0_7[116], stage0_7[117], stage0_7[118], stage0_7[119]},
      {stage1_9[19],stage1_8[40],stage1_7[40],stage1_6[46],stage1_5[63]}
   );
   gpc606_5 gpc95 (
      {stage0_5[120], stage0_5[121], stage0_5[122], stage0_5[123], stage0_5[124], stage0_5[125]},
      {stage0_7[120], stage0_7[121], stage0_7[122], stage0_7[123], stage0_7[124], stage0_7[125]},
      {stage1_9[20],stage1_8[41],stage1_7[41],stage1_6[47],stage1_5[64]}
   );
   gpc606_5 gpc96 (
      {stage0_5[126], stage0_5[127], stage0_5[128], stage0_5[129], stage0_5[130], stage0_5[131]},
      {stage0_7[126], stage0_7[127], stage0_7[128], stage0_7[129], stage0_7[130], stage0_7[131]},
      {stage1_9[21],stage1_8[42],stage1_7[42],stage1_6[48],stage1_5[65]}
   );
   gpc606_5 gpc97 (
      {stage0_5[132], stage0_5[133], stage0_5[134], stage0_5[135], stage0_5[136], stage0_5[137]},
      {stage0_7[132], stage0_7[133], stage0_7[134], stage0_7[135], stage0_7[136], stage0_7[137]},
      {stage1_9[22],stage1_8[43],stage1_7[43],stage1_6[49],stage1_5[66]}
   );
   gpc606_5 gpc98 (
      {stage0_5[138], stage0_5[139], stage0_5[140], stage0_5[141], stage0_5[142], stage0_5[143]},
      {stage0_7[138], stage0_7[139], stage0_7[140], stage0_7[141], stage0_7[142], stage0_7[143]},
      {stage1_9[23],stage1_8[44],stage1_7[44],stage1_6[50],stage1_5[67]}
   );
   gpc606_5 gpc99 (
      {stage0_5[144], stage0_5[145], stage0_5[146], stage0_5[147], stage0_5[148], stage0_5[149]},
      {stage0_7[144], stage0_7[145], stage0_7[146], stage0_7[147], stage0_7[148], stage0_7[149]},
      {stage1_9[24],stage1_8[45],stage1_7[45],stage1_6[51],stage1_5[68]}
   );
   gpc606_5 gpc100 (
      {stage0_5[150], stage0_5[151], stage0_5[152], stage0_5[153], stage0_5[154], stage0_5[155]},
      {stage0_7[150], stage0_7[151], stage0_7[152], stage0_7[153], stage0_7[154], stage0_7[155]},
      {stage1_9[25],stage1_8[46],stage1_7[46],stage1_6[52],stage1_5[69]}
   );
   gpc606_5 gpc101 (
      {stage0_5[156], stage0_5[157], stage0_5[158], stage0_5[159], stage0_5[160], stage0_5[161]},
      {stage0_7[156], stage0_7[157], stage0_7[158], stage0_7[159], stage0_7[160], stage0_7[161]},
      {stage1_9[26],stage1_8[47],stage1_7[47],stage1_6[53],stage1_5[70]}
   );
   gpc606_5 gpc102 (
      {stage0_6[126], stage0_6[127], stage0_6[128], stage0_6[129], stage0_6[130], stage0_6[131]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[27],stage1_8[48],stage1_7[48],stage1_6[54]}
   );
   gpc606_5 gpc103 (
      {stage0_6[132], stage0_6[133], stage0_6[134], stage0_6[135], stage0_6[136], stage0_6[137]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[28],stage1_8[49],stage1_7[49],stage1_6[55]}
   );
   gpc606_5 gpc104 (
      {stage0_6[138], stage0_6[139], stage0_6[140], stage0_6[141], stage0_6[142], stage0_6[143]},
      {stage0_8[12], stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17]},
      {stage1_10[2],stage1_9[29],stage1_8[50],stage1_7[50],stage1_6[56]}
   );
   gpc606_5 gpc105 (
      {stage0_6[144], stage0_6[145], stage0_6[146], stage0_6[147], stage0_6[148], stage0_6[149]},
      {stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage1_10[3],stage1_9[30],stage1_8[51],stage1_7[51],stage1_6[57]}
   );
   gpc606_5 gpc106 (
      {stage0_6[150], stage0_6[151], stage0_6[152], stage0_6[153], stage0_6[154], stage0_6[155]},
      {stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29]},
      {stage1_10[4],stage1_9[31],stage1_8[52],stage1_7[52],stage1_6[58]}
   );
   gpc606_5 gpc107 (
      {stage0_6[156], stage0_6[157], stage0_6[158], stage0_6[159], stage0_6[160], stage0_6[161]},
      {stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35]},
      {stage1_10[5],stage1_9[32],stage1_8[53],stage1_7[53],stage1_6[59]}
   );
   gpc606_5 gpc108 (
      {stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[0],stage1_10[6],stage1_9[33],stage1_8[54]}
   );
   gpc606_5 gpc109 (
      {stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[1],stage1_10[7],stage1_9[34],stage1_8[55]}
   );
   gpc606_5 gpc110 (
      {stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[2],stage1_10[8],stage1_9[35],stage1_8[56]}
   );
   gpc606_5 gpc111 (
      {stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[3],stage1_10[9],stage1_9[36],stage1_8[57]}
   );
   gpc606_5 gpc112 (
      {stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[4],stage1_10[10],stage1_9[37],stage1_8[58]}
   );
   gpc606_5 gpc113 (
      {stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[5],stage1_10[11],stage1_9[38],stage1_8[59]}
   );
   gpc615_5 gpc114 (
      {stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76]},
      {stage0_9[0]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[6],stage1_10[12],stage1_9[39],stage1_8[60]}
   );
   gpc615_5 gpc115 (
      {stage0_8[77], stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81]},
      {stage0_9[1]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[7],stage1_10[13],stage1_9[40],stage1_8[61]}
   );
   gpc615_5 gpc116 (
      {stage0_8[82], stage0_8[83], stage0_8[84], stage0_8[85], stage0_8[86]},
      {stage0_9[2]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[8],stage1_10[14],stage1_9[41],stage1_8[62]}
   );
   gpc615_5 gpc117 (
      {stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90], stage0_8[91]},
      {stage0_9[3]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[9],stage1_10[15],stage1_9[42],stage1_8[63]}
   );
   gpc615_5 gpc118 (
      {stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96]},
      {stage0_9[4]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[10],stage1_10[16],stage1_9[43],stage1_8[64]}
   );
   gpc615_5 gpc119 (
      {stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101]},
      {stage0_9[5]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[11],stage1_10[17],stage1_9[44],stage1_8[65]}
   );
   gpc615_5 gpc120 (
      {stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106]},
      {stage0_9[6]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[12],stage1_10[18],stage1_9[45],stage1_8[66]}
   );
   gpc615_5 gpc121 (
      {stage0_8[107], stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111]},
      {stage0_9[7]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[13],stage1_10[19],stage1_9[46],stage1_8[67]}
   );
   gpc615_5 gpc122 (
      {stage0_8[112], stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116]},
      {stage0_9[8]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[14],stage1_10[20],stage1_9[47],stage1_8[68]}
   );
   gpc615_5 gpc123 (
      {stage0_8[117], stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121]},
      {stage0_9[9]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[15],stage1_10[21],stage1_9[48],stage1_8[69]}
   );
   gpc615_5 gpc124 (
      {stage0_8[122], stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126]},
      {stage0_9[10]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[16],stage1_10[22],stage1_9[49],stage1_8[70]}
   );
   gpc615_5 gpc125 (
      {stage0_8[127], stage0_8[128], stage0_8[129], stage0_8[130], stage0_8[131]},
      {stage0_9[11]},
      {stage0_10[102], stage0_10[103], stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107]},
      {stage1_12[17],stage1_11[17],stage1_10[23],stage1_9[50],stage1_8[71]}
   );
   gpc615_5 gpc126 (
      {stage0_8[132], stage0_8[133], stage0_8[134], stage0_8[135], stage0_8[136]},
      {stage0_9[12]},
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113]},
      {stage1_12[18],stage1_11[18],stage1_10[24],stage1_9[51],stage1_8[72]}
   );
   gpc615_5 gpc127 (
      {stage0_8[137], stage0_8[138], stage0_8[139], stage0_8[140], stage0_8[141]},
      {stage0_9[13]},
      {stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117], stage0_10[118], stage0_10[119]},
      {stage1_12[19],stage1_11[19],stage1_10[25],stage1_9[52],stage1_8[73]}
   );
   gpc615_5 gpc128 (
      {stage0_8[142], stage0_8[143], stage0_8[144], stage0_8[145], stage0_8[146]},
      {stage0_9[14]},
      {stage0_10[120], stage0_10[121], stage0_10[122], stage0_10[123], stage0_10[124], stage0_10[125]},
      {stage1_12[20],stage1_11[20],stage1_10[26],stage1_9[53],stage1_8[74]}
   );
   gpc606_5 gpc129 (
      {stage0_9[15], stage0_9[16], stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[21],stage1_11[21],stage1_10[27],stage1_9[54]}
   );
   gpc606_5 gpc130 (
      {stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25], stage0_9[26]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[22],stage1_11[22],stage1_10[28],stage1_9[55]}
   );
   gpc606_5 gpc131 (
      {stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31], stage0_9[32]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[23],stage1_11[23],stage1_10[29],stage1_9[56]}
   );
   gpc606_5 gpc132 (
      {stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37], stage0_9[38]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[24],stage1_11[24],stage1_10[30],stage1_9[57]}
   );
   gpc606_5 gpc133 (
      {stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43], stage0_9[44]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[25],stage1_11[25],stage1_10[31],stage1_9[58]}
   );
   gpc606_5 gpc134 (
      {stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49], stage0_9[50]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[26],stage1_11[26],stage1_10[32],stage1_9[59]}
   );
   gpc606_5 gpc135 (
      {stage0_9[51], stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55], stage0_9[56]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[27],stage1_11[27],stage1_10[33],stage1_9[60]}
   );
   gpc606_5 gpc136 (
      {stage0_9[57], stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61], stage0_9[62]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[28],stage1_11[28],stage1_10[34],stage1_9[61]}
   );
   gpc606_5 gpc137 (
      {stage0_9[63], stage0_9[64], stage0_9[65], stage0_9[66], stage0_9[67], stage0_9[68]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[29],stage1_11[29],stage1_10[35],stage1_9[62]}
   );
   gpc606_5 gpc138 (
      {stage0_9[69], stage0_9[70], stage0_9[71], stage0_9[72], stage0_9[73], stage0_9[74]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[30],stage1_11[30],stage1_10[36],stage1_9[63]}
   );
   gpc606_5 gpc139 (
      {stage0_9[75], stage0_9[76], stage0_9[77], stage0_9[78], stage0_9[79], stage0_9[80]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[31],stage1_11[31],stage1_10[37],stage1_9[64]}
   );
   gpc606_5 gpc140 (
      {stage0_9[81], stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85], stage0_9[86]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[32],stage1_11[32],stage1_10[38],stage1_9[65]}
   );
   gpc606_5 gpc141 (
      {stage0_9[87], stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91], stage0_9[92]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[33],stage1_11[33],stage1_10[39],stage1_9[66]}
   );
   gpc606_5 gpc142 (
      {stage0_9[93], stage0_9[94], stage0_9[95], stage0_9[96], stage0_9[97], stage0_9[98]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[34],stage1_11[34],stage1_10[40],stage1_9[67]}
   );
   gpc606_5 gpc143 (
      {stage0_9[99], stage0_9[100], stage0_9[101], stage0_9[102], stage0_9[103], stage0_9[104]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[35],stage1_11[35],stage1_10[41],stage1_9[68]}
   );
   gpc606_5 gpc144 (
      {stage0_9[105], stage0_9[106], stage0_9[107], stage0_9[108], stage0_9[109], stage0_9[110]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[36],stage1_11[36],stage1_10[42],stage1_9[69]}
   );
   gpc606_5 gpc145 (
      {stage0_9[111], stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115], stage0_9[116]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[37],stage1_11[37],stage1_10[43],stage1_9[70]}
   );
   gpc606_5 gpc146 (
      {stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120], stage0_9[121], stage0_9[122]},
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage1_13[17],stage1_12[38],stage1_11[38],stage1_10[44],stage1_9[71]}
   );
   gpc606_5 gpc147 (
      {stage0_9[123], stage0_9[124], stage0_9[125], stage0_9[126], stage0_9[127], stage0_9[128]},
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112], stage0_11[113]},
      {stage1_13[18],stage1_12[39],stage1_11[39],stage1_10[45],stage1_9[72]}
   );
   gpc606_5 gpc148 (
      {stage0_9[129], stage0_9[130], stage0_9[131], stage0_9[132], stage0_9[133], stage0_9[134]},
      {stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117], stage0_11[118], stage0_11[119]},
      {stage1_13[19],stage1_12[40],stage1_11[40],stage1_10[46],stage1_9[73]}
   );
   gpc606_5 gpc149 (
      {stage0_9[135], stage0_9[136], stage0_9[137], stage0_9[138], stage0_9[139], stage0_9[140]},
      {stage0_11[120], stage0_11[121], stage0_11[122], stage0_11[123], stage0_11[124], stage0_11[125]},
      {stage1_13[20],stage1_12[41],stage1_11[41],stage1_10[47],stage1_9[74]}
   );
   gpc606_5 gpc150 (
      {stage0_9[141], stage0_9[142], stage0_9[143], stage0_9[144], stage0_9[145], stage0_9[146]},
      {stage0_11[126], stage0_11[127], stage0_11[128], stage0_11[129], stage0_11[130], stage0_11[131]},
      {stage1_13[21],stage1_12[42],stage1_11[42],stage1_10[48],stage1_9[75]}
   );
   gpc615_5 gpc151 (
      {stage0_9[147], stage0_9[148], stage0_9[149], stage0_9[150], stage0_9[151]},
      {stage0_10[126]},
      {stage0_11[132], stage0_11[133], stage0_11[134], stage0_11[135], stage0_11[136], stage0_11[137]},
      {stage1_13[22],stage1_12[43],stage1_11[43],stage1_10[49],stage1_9[76]}
   );
   gpc615_5 gpc152 (
      {stage0_9[152], stage0_9[153], stage0_9[154], stage0_9[155], stage0_9[156]},
      {stage0_10[127]},
      {stage0_11[138], stage0_11[139], stage0_11[140], stage0_11[141], stage0_11[142], stage0_11[143]},
      {stage1_13[23],stage1_12[44],stage1_11[44],stage1_10[50],stage1_9[77]}
   );
   gpc615_5 gpc153 (
      {stage0_10[128], stage0_10[129], stage0_10[130], stage0_10[131], stage0_10[132]},
      {stage0_11[144]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[24],stage1_12[45],stage1_11[45],stage1_10[51]}
   );
   gpc615_5 gpc154 (
      {stage0_10[133], stage0_10[134], stage0_10[135], stage0_10[136], stage0_10[137]},
      {stage0_11[145]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[25],stage1_12[46],stage1_11[46],stage1_10[52]}
   );
   gpc615_5 gpc155 (
      {stage0_10[138], stage0_10[139], stage0_10[140], stage0_10[141], stage0_10[142]},
      {stage0_11[146]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[26],stage1_12[47],stage1_11[47],stage1_10[53]}
   );
   gpc615_5 gpc156 (
      {stage0_10[143], stage0_10[144], stage0_10[145], stage0_10[146], stage0_10[147]},
      {stage0_11[147]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[27],stage1_12[48],stage1_11[48],stage1_10[54]}
   );
   gpc615_5 gpc157 (
      {stage0_10[148], stage0_10[149], stage0_10[150], stage0_10[151], stage0_10[152]},
      {stage0_11[148]},
      {stage0_12[24], stage0_12[25], stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29]},
      {stage1_14[4],stage1_13[28],stage1_12[49],stage1_11[49],stage1_10[55]}
   );
   gpc615_5 gpc158 (
      {stage0_10[153], stage0_10[154], stage0_10[155], stage0_10[156], stage0_10[157]},
      {stage0_11[149]},
      {stage0_12[30], stage0_12[31], stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35]},
      {stage1_14[5],stage1_13[29],stage1_12[50],stage1_11[50],stage1_10[56]}
   );
   gpc606_5 gpc159 (
      {stage0_11[150], stage0_11[151], stage0_11[152], stage0_11[153], stage0_11[154], stage0_11[155]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[6],stage1_13[30],stage1_12[51],stage1_11[51]}
   );
   gpc606_5 gpc160 (
      {stage0_12[36], stage0_12[37], stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[1],stage1_14[7],stage1_13[31],stage1_12[52]}
   );
   gpc606_5 gpc161 (
      {stage0_12[42], stage0_12[43], stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[2],stage1_14[8],stage1_13[32],stage1_12[53]}
   );
   gpc606_5 gpc162 (
      {stage0_12[48], stage0_12[49], stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[3],stage1_14[9],stage1_13[33],stage1_12[54]}
   );
   gpc606_5 gpc163 (
      {stage0_12[54], stage0_12[55], stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[4],stage1_14[10],stage1_13[34],stage1_12[55]}
   );
   gpc606_5 gpc164 (
      {stage0_12[60], stage0_12[61], stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[5],stage1_14[11],stage1_13[35],stage1_12[56]}
   );
   gpc606_5 gpc165 (
      {stage0_12[66], stage0_12[67], stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[6],stage1_14[12],stage1_13[36],stage1_12[57]}
   );
   gpc606_5 gpc166 (
      {stage0_12[72], stage0_12[73], stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[7],stage1_14[13],stage1_13[37],stage1_12[58]}
   );
   gpc606_5 gpc167 (
      {stage0_12[78], stage0_12[79], stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[8],stage1_14[14],stage1_13[38],stage1_12[59]}
   );
   gpc606_5 gpc168 (
      {stage0_12[84], stage0_12[85], stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[9],stage1_14[15],stage1_13[39],stage1_12[60]}
   );
   gpc606_5 gpc169 (
      {stage0_12[90], stage0_12[91], stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[10],stage1_14[16],stage1_13[40],stage1_12[61]}
   );
   gpc606_5 gpc170 (
      {stage0_12[96], stage0_12[97], stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[11],stage1_14[17],stage1_13[41],stage1_12[62]}
   );
   gpc606_5 gpc171 (
      {stage0_12[102], stage0_12[103], stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[12],stage1_14[18],stage1_13[42],stage1_12[63]}
   );
   gpc606_5 gpc172 (
      {stage0_12[108], stage0_12[109], stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[13],stage1_14[19],stage1_13[43],stage1_12[64]}
   );
   gpc606_5 gpc173 (
      {stage0_12[114], stage0_12[115], stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[14],stage1_14[20],stage1_13[44],stage1_12[65]}
   );
   gpc606_5 gpc174 (
      {stage0_12[120], stage0_12[121], stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[15],stage1_14[21],stage1_13[45],stage1_12[66]}
   );
   gpc606_5 gpc175 (
      {stage0_12[126], stage0_12[127], stage0_12[128], stage0_12[129], stage0_12[130], stage0_12[131]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[16],stage1_14[22],stage1_13[46],stage1_12[67]}
   );
   gpc606_5 gpc176 (
      {stage0_12[132], stage0_12[133], stage0_12[134], stage0_12[135], stage0_12[136], stage0_12[137]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[17],stage1_14[23],stage1_13[47],stage1_12[68]}
   );
   gpc606_5 gpc177 (
      {stage0_12[138], stage0_12[139], stage0_12[140], stage0_12[141], stage0_12[142], stage0_12[143]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[18],stage1_14[24],stage1_13[48],stage1_12[69]}
   );
   gpc606_5 gpc178 (
      {stage0_12[144], stage0_12[145], stage0_12[146], stage0_12[147], stage0_12[148], stage0_12[149]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[19],stage1_14[25],stage1_13[49],stage1_12[70]}
   );
   gpc606_5 gpc179 (
      {stage0_12[150], stage0_12[151], stage0_12[152], stage0_12[153], stage0_12[154], stage0_12[155]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[20],stage1_14[26],stage1_13[50],stage1_12[71]}
   );
   gpc606_5 gpc180 (
      {stage0_12[156], stage0_12[157], stage0_12[158], stage0_12[159], stage0_12[160], stage0_12[161]},
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124], stage0_14[125]},
      {stage1_16[20],stage1_15[21],stage1_14[27],stage1_13[51],stage1_12[72]}
   );
   gpc606_5 gpc181 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[21],stage1_15[22],stage1_14[28],stage1_13[52]}
   );
   gpc606_5 gpc182 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[22],stage1_15[23],stage1_14[29],stage1_13[53]}
   );
   gpc606_5 gpc183 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[23],stage1_15[24],stage1_14[30],stage1_13[54]}
   );
   gpc606_5 gpc184 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[24],stage1_15[25],stage1_14[31],stage1_13[55]}
   );
   gpc606_5 gpc185 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[25],stage1_15[26],stage1_14[32],stage1_13[56]}
   );
   gpc606_5 gpc186 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[26],stage1_15[27],stage1_14[33],stage1_13[57]}
   );
   gpc606_5 gpc187 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[27],stage1_15[28],stage1_14[34],stage1_13[58]}
   );
   gpc606_5 gpc188 (
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[28],stage1_15[29],stage1_14[35],stage1_13[59]}
   );
   gpc606_5 gpc189 (
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[29],stage1_15[30],stage1_14[36],stage1_13[60]}
   );
   gpc606_5 gpc190 (
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[30],stage1_15[31],stage1_14[37],stage1_13[61]}
   );
   gpc606_5 gpc191 (
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[31],stage1_15[32],stage1_14[38],stage1_13[62]}
   );
   gpc606_5 gpc192 (
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[32],stage1_15[33],stage1_14[39],stage1_13[63]}
   );
   gpc606_5 gpc193 (
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[33],stage1_15[34],stage1_14[40],stage1_13[64]}
   );
   gpc606_5 gpc194 (
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[34],stage1_15[35],stage1_14[41],stage1_13[65]}
   );
   gpc606_5 gpc195 (
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[35],stage1_15[36],stage1_14[42],stage1_13[66]}
   );
   gpc606_5 gpc196 (
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[36],stage1_15[37],stage1_14[43],stage1_13[67]}
   );
   gpc606_5 gpc197 (
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[37],stage1_15[38],stage1_14[44],stage1_13[68]}
   );
   gpc606_5 gpc198 (
      {stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[38],stage1_15[39],stage1_14[45],stage1_13[69]}
   );
   gpc606_5 gpc199 (
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[39],stage1_15[40],stage1_14[46],stage1_13[70]}
   );
   gpc606_5 gpc200 (
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage0_15[114], stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage1_17[19],stage1_16[40],stage1_15[41],stage1_14[47],stage1_13[71]}
   );
   gpc606_5 gpc201 (
      {stage0_13[126], stage0_13[127], stage0_13[128], stage0_13[129], stage0_13[130], stage0_13[131]},
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124], stage0_15[125]},
      {stage1_17[20],stage1_16[41],stage1_15[42],stage1_14[48],stage1_13[72]}
   );
   gpc606_5 gpc202 (
      {stage0_13[132], stage0_13[133], stage0_13[134], stage0_13[135], stage0_13[136], stage0_13[137]},
      {stage0_15[126], stage0_15[127], stage0_15[128], stage0_15[129], stage0_15[130], stage0_15[131]},
      {stage1_17[21],stage1_16[42],stage1_15[43],stage1_14[49],stage1_13[73]}
   );
   gpc606_5 gpc203 (
      {stage0_13[138], stage0_13[139], stage0_13[140], stage0_13[141], stage0_13[142], stage0_13[143]},
      {stage0_15[132], stage0_15[133], stage0_15[134], stage0_15[135], stage0_15[136], stage0_15[137]},
      {stage1_17[22],stage1_16[43],stage1_15[44],stage1_14[50],stage1_13[74]}
   );
   gpc606_5 gpc204 (
      {stage0_13[144], stage0_13[145], stage0_13[146], stage0_13[147], stage0_13[148], stage0_13[149]},
      {stage0_15[138], stage0_15[139], stage0_15[140], stage0_15[141], stage0_15[142], stage0_15[143]},
      {stage1_17[23],stage1_16[44],stage1_15[45],stage1_14[51],stage1_13[75]}
   );
   gpc606_5 gpc205 (
      {stage0_13[150], stage0_13[151], stage0_13[152], stage0_13[153], stage0_13[154], stage0_13[155]},
      {stage0_15[144], stage0_15[145], stage0_15[146], stage0_15[147], stage0_15[148], stage0_15[149]},
      {stage1_17[24],stage1_16[45],stage1_15[46],stage1_14[52],stage1_13[76]}
   );
   gpc606_5 gpc206 (
      {stage0_13[156], stage0_13[157], stage0_13[158], stage0_13[159], stage0_13[160], stage0_13[161]},
      {stage0_15[150], stage0_15[151], stage0_15[152], stage0_15[153], stage0_15[154], stage0_15[155]},
      {stage1_17[25],stage1_16[46],stage1_15[47],stage1_14[53],stage1_13[77]}
   );
   gpc117_4 gpc207 (
      {stage0_14[126], stage0_14[127], stage0_14[128], stage0_14[129], stage0_14[130], stage0_14[131], stage0_14[132]},
      {stage0_15[156]},
      {1'b0},
      {stage1_17[26],stage1_16[47],stage1_15[48],stage1_14[54]}
   );
   gpc117_4 gpc208 (
      {stage0_14[133], stage0_14[134], stage0_14[135], stage0_14[136], stage0_14[137], stage0_14[138], stage0_14[139]},
      {stage0_15[157]},
      {1'b0},
      {stage1_17[27],stage1_16[48],stage1_15[49],stage1_14[55]}
   );
   gpc1_1 gpc209 (
      {stage0_0[160]},
      {stage1_0[31]}
   );
   gpc1_1 gpc210 (
      {stage0_0[161]},
      {stage1_0[32]}
   );
   gpc1_1 gpc211 (
      {stage0_2[152]},
      {stage1_2[54]}
   );
   gpc1_1 gpc212 (
      {stage0_2[153]},
      {stage1_2[55]}
   );
   gpc1_1 gpc213 (
      {stage0_2[154]},
      {stage1_2[56]}
   );
   gpc1_1 gpc214 (
      {stage0_2[155]},
      {stage1_2[57]}
   );
   gpc1_1 gpc215 (
      {stage0_2[156]},
      {stage1_2[58]}
   );
   gpc1_1 gpc216 (
      {stage0_2[157]},
      {stage1_2[59]}
   );
   gpc1_1 gpc217 (
      {stage0_2[158]},
      {stage1_2[60]}
   );
   gpc1_1 gpc218 (
      {stage0_2[159]},
      {stage1_2[61]}
   );
   gpc1_1 gpc219 (
      {stage0_2[160]},
      {stage1_2[62]}
   );
   gpc1_1 gpc220 (
      {stage0_2[161]},
      {stage1_2[63]}
   );
   gpc1_1 gpc221 (
      {stage0_3[124]},
      {stage1_3[54]}
   );
   gpc1_1 gpc222 (
      {stage0_3[125]},
      {stage1_3[55]}
   );
   gpc1_1 gpc223 (
      {stage0_3[126]},
      {stage1_3[56]}
   );
   gpc1_1 gpc224 (
      {stage0_3[127]},
      {stage1_3[57]}
   );
   gpc1_1 gpc225 (
      {stage0_3[128]},
      {stage1_3[58]}
   );
   gpc1_1 gpc226 (
      {stage0_3[129]},
      {stage1_3[59]}
   );
   gpc1_1 gpc227 (
      {stage0_3[130]},
      {stage1_3[60]}
   );
   gpc1_1 gpc228 (
      {stage0_3[131]},
      {stage1_3[61]}
   );
   gpc1_1 gpc229 (
      {stage0_3[132]},
      {stage1_3[62]}
   );
   gpc1_1 gpc230 (
      {stage0_3[133]},
      {stage1_3[63]}
   );
   gpc1_1 gpc231 (
      {stage0_3[134]},
      {stage1_3[64]}
   );
   gpc1_1 gpc232 (
      {stage0_3[135]},
      {stage1_3[65]}
   );
   gpc1_1 gpc233 (
      {stage0_3[136]},
      {stage1_3[66]}
   );
   gpc1_1 gpc234 (
      {stage0_3[137]},
      {stage1_3[67]}
   );
   gpc1_1 gpc235 (
      {stage0_3[138]},
      {stage1_3[68]}
   );
   gpc1_1 gpc236 (
      {stage0_3[139]},
      {stage1_3[69]}
   );
   gpc1_1 gpc237 (
      {stage0_3[140]},
      {stage1_3[70]}
   );
   gpc1_1 gpc238 (
      {stage0_3[141]},
      {stage1_3[71]}
   );
   gpc1_1 gpc239 (
      {stage0_3[142]},
      {stage1_3[72]}
   );
   gpc1_1 gpc240 (
      {stage0_3[143]},
      {stage1_3[73]}
   );
   gpc1_1 gpc241 (
      {stage0_3[144]},
      {stage1_3[74]}
   );
   gpc1_1 gpc242 (
      {stage0_3[145]},
      {stage1_3[75]}
   );
   gpc1_1 gpc243 (
      {stage0_3[146]},
      {stage1_3[76]}
   );
   gpc1_1 gpc244 (
      {stage0_3[147]},
      {stage1_3[77]}
   );
   gpc1_1 gpc245 (
      {stage0_3[148]},
      {stage1_3[78]}
   );
   gpc1_1 gpc246 (
      {stage0_3[149]},
      {stage1_3[79]}
   );
   gpc1_1 gpc247 (
      {stage0_3[150]},
      {stage1_3[80]}
   );
   gpc1_1 gpc248 (
      {stage0_3[151]},
      {stage1_3[81]}
   );
   gpc1_1 gpc249 (
      {stage0_3[152]},
      {stage1_3[82]}
   );
   gpc1_1 gpc250 (
      {stage0_3[153]},
      {stage1_3[83]}
   );
   gpc1_1 gpc251 (
      {stage0_3[154]},
      {stage1_3[84]}
   );
   gpc1_1 gpc252 (
      {stage0_3[155]},
      {stage1_3[85]}
   );
   gpc1_1 gpc253 (
      {stage0_3[156]},
      {stage1_3[86]}
   );
   gpc1_1 gpc254 (
      {stage0_3[157]},
      {stage1_3[87]}
   );
   gpc1_1 gpc255 (
      {stage0_3[158]},
      {stage1_3[88]}
   );
   gpc1_1 gpc256 (
      {stage0_3[159]},
      {stage1_3[89]}
   );
   gpc1_1 gpc257 (
      {stage0_3[160]},
      {stage1_3[90]}
   );
   gpc1_1 gpc258 (
      {stage0_3[161]},
      {stage1_3[91]}
   );
   gpc1_1 gpc259 (
      {stage0_8[147]},
      {stage1_8[75]}
   );
   gpc1_1 gpc260 (
      {stage0_8[148]},
      {stage1_8[76]}
   );
   gpc1_1 gpc261 (
      {stage0_8[149]},
      {stage1_8[77]}
   );
   gpc1_1 gpc262 (
      {stage0_8[150]},
      {stage1_8[78]}
   );
   gpc1_1 gpc263 (
      {stage0_8[151]},
      {stage1_8[79]}
   );
   gpc1_1 gpc264 (
      {stage0_8[152]},
      {stage1_8[80]}
   );
   gpc1_1 gpc265 (
      {stage0_8[153]},
      {stage1_8[81]}
   );
   gpc1_1 gpc266 (
      {stage0_8[154]},
      {stage1_8[82]}
   );
   gpc1_1 gpc267 (
      {stage0_8[155]},
      {stage1_8[83]}
   );
   gpc1_1 gpc268 (
      {stage0_8[156]},
      {stage1_8[84]}
   );
   gpc1_1 gpc269 (
      {stage0_8[157]},
      {stage1_8[85]}
   );
   gpc1_1 gpc270 (
      {stage0_8[158]},
      {stage1_8[86]}
   );
   gpc1_1 gpc271 (
      {stage0_8[159]},
      {stage1_8[87]}
   );
   gpc1_1 gpc272 (
      {stage0_8[160]},
      {stage1_8[88]}
   );
   gpc1_1 gpc273 (
      {stage0_8[161]},
      {stage1_8[89]}
   );
   gpc1_1 gpc274 (
      {stage0_9[157]},
      {stage1_9[78]}
   );
   gpc1_1 gpc275 (
      {stage0_9[158]},
      {stage1_9[79]}
   );
   gpc1_1 gpc276 (
      {stage0_9[159]},
      {stage1_9[80]}
   );
   gpc1_1 gpc277 (
      {stage0_9[160]},
      {stage1_9[81]}
   );
   gpc1_1 gpc278 (
      {stage0_9[161]},
      {stage1_9[82]}
   );
   gpc1_1 gpc279 (
      {stage0_10[158]},
      {stage1_10[57]}
   );
   gpc1_1 gpc280 (
      {stage0_10[159]},
      {stage1_10[58]}
   );
   gpc1_1 gpc281 (
      {stage0_10[160]},
      {stage1_10[59]}
   );
   gpc1_1 gpc282 (
      {stage0_10[161]},
      {stage1_10[60]}
   );
   gpc1_1 gpc283 (
      {stage0_11[156]},
      {stage1_11[52]}
   );
   gpc1_1 gpc284 (
      {stage0_11[157]},
      {stage1_11[53]}
   );
   gpc1_1 gpc285 (
      {stage0_11[158]},
      {stage1_11[54]}
   );
   gpc1_1 gpc286 (
      {stage0_11[159]},
      {stage1_11[55]}
   );
   gpc1_1 gpc287 (
      {stage0_11[160]},
      {stage1_11[56]}
   );
   gpc1_1 gpc288 (
      {stage0_11[161]},
      {stage1_11[57]}
   );
   gpc1_1 gpc289 (
      {stage0_14[140]},
      {stage1_14[56]}
   );
   gpc1_1 gpc290 (
      {stage0_14[141]},
      {stage1_14[57]}
   );
   gpc1_1 gpc291 (
      {stage0_14[142]},
      {stage1_14[58]}
   );
   gpc1_1 gpc292 (
      {stage0_14[143]},
      {stage1_14[59]}
   );
   gpc1_1 gpc293 (
      {stage0_14[144]},
      {stage1_14[60]}
   );
   gpc1_1 gpc294 (
      {stage0_14[145]},
      {stage1_14[61]}
   );
   gpc1_1 gpc295 (
      {stage0_14[146]},
      {stage1_14[62]}
   );
   gpc1_1 gpc296 (
      {stage0_14[147]},
      {stage1_14[63]}
   );
   gpc1_1 gpc297 (
      {stage0_14[148]},
      {stage1_14[64]}
   );
   gpc1_1 gpc298 (
      {stage0_14[149]},
      {stage1_14[65]}
   );
   gpc1_1 gpc299 (
      {stage0_14[150]},
      {stage1_14[66]}
   );
   gpc1_1 gpc300 (
      {stage0_14[151]},
      {stage1_14[67]}
   );
   gpc1_1 gpc301 (
      {stage0_14[152]},
      {stage1_14[68]}
   );
   gpc1_1 gpc302 (
      {stage0_14[153]},
      {stage1_14[69]}
   );
   gpc1_1 gpc303 (
      {stage0_14[154]},
      {stage1_14[70]}
   );
   gpc1_1 gpc304 (
      {stage0_14[155]},
      {stage1_14[71]}
   );
   gpc1_1 gpc305 (
      {stage0_14[156]},
      {stage1_14[72]}
   );
   gpc1_1 gpc306 (
      {stage0_14[157]},
      {stage1_14[73]}
   );
   gpc1_1 gpc307 (
      {stage0_14[158]},
      {stage1_14[74]}
   );
   gpc1_1 gpc308 (
      {stage0_14[159]},
      {stage1_14[75]}
   );
   gpc1_1 gpc309 (
      {stage0_14[160]},
      {stage1_14[76]}
   );
   gpc1_1 gpc310 (
      {stage0_14[161]},
      {stage1_14[77]}
   );
   gpc1_1 gpc311 (
      {stage0_15[158]},
      {stage1_15[50]}
   );
   gpc1_1 gpc312 (
      {stage0_15[159]},
      {stage1_15[51]}
   );
   gpc1_1 gpc313 (
      {stage0_15[160]},
      {stage1_15[52]}
   );
   gpc1_1 gpc314 (
      {stage0_15[161]},
      {stage1_15[53]}
   );
   gpc606_5 gpc315 (
      {stage1_0[0], stage1_0[1], stage1_0[2], stage1_0[3], stage1_0[4], stage1_0[5]},
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc606_5 gpc316 (
      {stage1_0[6], stage1_0[7], stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11]},
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc317 (
      {stage1_0[12], stage1_0[13], stage1_0[14], stage1_0[15], stage1_0[16]},
      {stage1_1[0]},
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc615_5 gpc318 (
      {stage1_0[17], stage1_0[18], stage1_0[19], stage1_0[20], stage1_0[21]},
      {stage1_1[1]},
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23]},
      {stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3],stage2_0[3]}
   );
   gpc615_5 gpc319 (
      {stage1_0[22], stage1_0[23], stage1_0[24], stage1_0[25], stage1_0[26]},
      {stage1_1[2]},
      {stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29]},
      {stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4],stage2_0[4]}
   );
   gpc606_5 gpc320 (
      {stage1_1[3], stage1_1[4], stage1_1[5], stage1_1[6], stage1_1[7], stage1_1[8]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5]}
   );
   gpc606_5 gpc321 (
      {stage1_1[9], stage1_1[10], stage1_1[11], stage1_1[12], stage1_1[13], stage1_1[14]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[1],stage2_4[6],stage2_3[6],stage2_2[6],stage2_1[6]}
   );
   gpc606_5 gpc322 (
      {stage1_1[15], stage1_1[16], stage1_1[17], stage1_1[18], stage1_1[19], stage1_1[20]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[2],stage2_4[7],stage2_3[7],stage2_2[7],stage2_1[7]}
   );
   gpc606_5 gpc323 (
      {stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25], stage1_1[26]},
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage2_5[3],stage2_4[8],stage2_3[8],stage2_2[8],stage2_1[8]}
   );
   gpc615_5 gpc324 (
      {stage1_2[30], stage1_2[31], stage1_2[32], stage1_2[33], stage1_2[34]},
      {stage1_3[24]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[4],stage2_4[9],stage2_3[9],stage2_2[9]}
   );
   gpc615_5 gpc325 (
      {stage1_2[35], stage1_2[36], stage1_2[37], stage1_2[38], stage1_2[39]},
      {stage1_3[25]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[5],stage2_4[10],stage2_3[10],stage2_2[10]}
   );
   gpc615_5 gpc326 (
      {stage1_2[40], stage1_2[41], stage1_2[42], stage1_2[43], stage1_2[44]},
      {stage1_3[26]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[6],stage2_4[11],stage2_3[11],stage2_2[11]}
   );
   gpc615_5 gpc327 (
      {stage1_2[45], stage1_2[46], stage1_2[47], stage1_2[48], stage1_2[49]},
      {stage1_3[27]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[7],stage2_4[12],stage2_3[12],stage2_2[12]}
   );
   gpc615_5 gpc328 (
      {stage1_2[50], stage1_2[51], stage1_2[52], stage1_2[53], stage1_2[54]},
      {stage1_3[28]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[8],stage2_4[13],stage2_3[13],stage2_2[13]}
   );
   gpc615_5 gpc329 (
      {stage1_2[55], stage1_2[56], stage1_2[57], stage1_2[58], stage1_2[59]},
      {stage1_3[29]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[9],stage2_4[14],stage2_3[14],stage2_2[14]}
   );
   gpc615_5 gpc330 (
      {stage1_2[60], stage1_2[61], stage1_2[62], stage1_2[63], 1'b0},
      {stage1_3[30]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[10],stage2_4[15],stage2_3[15],stage2_2[15]}
   );
   gpc615_5 gpc331 (
      {stage1_3[31], stage1_3[32], stage1_3[33], stage1_3[34], stage1_3[35]},
      {stage1_4[42]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[7],stage2_5[11],stage2_4[16],stage2_3[16]}
   );
   gpc615_5 gpc332 (
      {stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39], stage1_3[40]},
      {stage1_4[43]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[8],stage2_5[12],stage2_4[17],stage2_3[17]}
   );
   gpc615_5 gpc333 (
      {stage1_3[41], stage1_3[42], stage1_3[43], stage1_3[44], stage1_3[45]},
      {stage1_4[44]},
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage2_7[2],stage2_6[9],stage2_5[13],stage2_4[18],stage2_3[18]}
   );
   gpc615_5 gpc334 (
      {stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49], stage1_3[50]},
      {stage1_4[45]},
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage2_7[3],stage2_6[10],stage2_5[14],stage2_4[19],stage2_3[19]}
   );
   gpc615_5 gpc335 (
      {stage1_3[51], stage1_3[52], stage1_3[53], stage1_3[54], stage1_3[55]},
      {stage1_4[46]},
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage2_7[4],stage2_6[11],stage2_5[15],stage2_4[20],stage2_3[20]}
   );
   gpc615_5 gpc336 (
      {stage1_3[56], stage1_3[57], stage1_3[58], stage1_3[59], stage1_3[60]},
      {stage1_4[47]},
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage2_7[5],stage2_6[12],stage2_5[16],stage2_4[21],stage2_3[21]}
   );
   gpc615_5 gpc337 (
      {stage1_3[61], stage1_3[62], stage1_3[63], stage1_3[64], stage1_3[65]},
      {stage1_4[48]},
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage2_7[6],stage2_6[13],stage2_5[17],stage2_4[22],stage2_3[22]}
   );
   gpc615_5 gpc338 (
      {stage1_3[66], stage1_3[67], stage1_3[68], stage1_3[69], stage1_3[70]},
      {stage1_4[49]},
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage2_7[7],stage2_6[14],stage2_5[18],stage2_4[23],stage2_3[23]}
   );
   gpc615_5 gpc339 (
      {stage1_3[71], stage1_3[72], stage1_3[73], stage1_3[74], stage1_3[75]},
      {stage1_4[50]},
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage2_7[8],stage2_6[15],stage2_5[19],stage2_4[24],stage2_3[24]}
   );
   gpc615_5 gpc340 (
      {stage1_3[76], stage1_3[77], stage1_3[78], stage1_3[79], stage1_3[80]},
      {stage1_4[51]},
      {stage1_5[54], stage1_5[55], stage1_5[56], stage1_5[57], stage1_5[58], stage1_5[59]},
      {stage2_7[9],stage2_6[16],stage2_5[20],stage2_4[25],stage2_3[25]}
   );
   gpc606_5 gpc341 (
      {stage1_4[52], stage1_4[53], stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[10],stage2_6[17],stage2_5[21],stage2_4[26]}
   );
   gpc606_5 gpc342 (
      {stage1_4[58], stage1_4[59], stage1_4[60], stage1_4[61], stage1_4[62], stage1_4[63]},
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage2_8[1],stage2_7[11],stage2_6[18],stage2_5[22],stage2_4[27]}
   );
   gpc606_5 gpc343 (
      {stage1_4[64], stage1_4[65], stage1_4[66], stage1_4[67], stage1_4[68], stage1_4[69]},
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage2_8[2],stage2_7[12],stage2_6[19],stage2_5[23],stage2_4[28]}
   );
   gpc615_5 gpc344 (
      {stage1_4[70], stage1_4[71], stage1_4[72], stage1_4[73], stage1_4[74]},
      {stage1_5[60]},
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23]},
      {stage2_8[3],stage2_7[13],stage2_6[20],stage2_5[24],stage2_4[29]}
   );
   gpc606_5 gpc345 (
      {stage1_5[61], stage1_5[62], stage1_5[63], stage1_5[64], stage1_5[65], stage1_5[66]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[4],stage2_7[14],stage2_6[21],stage2_5[25]}
   );
   gpc606_5 gpc346 (
      {stage1_6[24], stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[1],stage2_8[5],stage2_7[15],stage2_6[22]}
   );
   gpc606_5 gpc347 (
      {stage1_6[30], stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[2],stage2_8[6],stage2_7[16],stage2_6[23]}
   );
   gpc606_5 gpc348 (
      {stage1_6[36], stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[3],stage2_8[7],stage2_7[17],stage2_6[24]}
   );
   gpc606_5 gpc349 (
      {stage1_6[42], stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[4],stage2_8[8],stage2_7[18],stage2_6[25]}
   );
   gpc615_5 gpc350 (
      {stage1_6[48], stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52]},
      {stage1_7[6]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[5],stage2_8[9],stage2_7[19],stage2_6[26]}
   );
   gpc615_5 gpc351 (
      {stage1_6[53], stage1_6[54], stage1_6[55], stage1_6[56], stage1_6[57]},
      {stage1_7[7]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[6],stage2_8[10],stage2_7[20],stage2_6[27]}
   );
   gpc615_5 gpc352 (
      {stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage1_8[36]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[6],stage2_9[7],stage2_8[11],stage2_7[21]}
   );
   gpc615_5 gpc353 (
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage1_8[37]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[7],stage2_9[8],stage2_8[12],stage2_7[22]}
   );
   gpc615_5 gpc354 (
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22]},
      {stage1_8[38]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[8],stage2_9[9],stage2_8[13],stage2_7[23]}
   );
   gpc615_5 gpc355 (
      {stage1_7[23], stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27]},
      {stage1_8[39]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[9],stage2_9[10],stage2_8[14],stage2_7[24]}
   );
   gpc615_5 gpc356 (
      {stage1_7[28], stage1_7[29], stage1_7[30], stage1_7[31], stage1_7[32]},
      {stage1_8[40]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[10],stage2_9[11],stage2_8[15],stage2_7[25]}
   );
   gpc615_5 gpc357 (
      {stage1_7[33], stage1_7[34], stage1_7[35], stage1_7[36], stage1_7[37]},
      {stage1_8[41]},
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage2_11[5],stage2_10[11],stage2_9[12],stage2_8[16],stage2_7[26]}
   );
   gpc615_5 gpc358 (
      {stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41], stage1_7[42]},
      {stage1_8[42]},
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage2_11[6],stage2_10[12],stage2_9[13],stage2_8[17],stage2_7[27]}
   );
   gpc606_5 gpc359 (
      {stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47], stage1_8[48]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[7],stage2_10[13],stage2_9[14],stage2_8[18]}
   );
   gpc606_5 gpc360 (
      {stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53], stage1_8[54]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[8],stage2_10[14],stage2_9[15],stage2_8[19]}
   );
   gpc606_5 gpc361 (
      {stage1_8[55], stage1_8[56], stage1_8[57], stage1_8[58], stage1_8[59], stage1_8[60]},
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage2_12[2],stage2_11[9],stage2_10[15],stage2_9[16],stage2_8[20]}
   );
   gpc606_5 gpc362 (
      {stage1_8[61], stage1_8[62], stage1_8[63], stage1_8[64], stage1_8[65], stage1_8[66]},
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage2_12[3],stage2_11[10],stage2_10[16],stage2_9[17],stage2_8[21]}
   );
   gpc606_5 gpc363 (
      {stage1_8[67], stage1_8[68], stage1_8[69], stage1_8[70], stage1_8[71], stage1_8[72]},
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage2_12[4],stage2_11[11],stage2_10[17],stage2_9[18],stage2_8[22]}
   );
   gpc606_5 gpc364 (
      {stage1_8[73], stage1_8[74], stage1_8[75], stage1_8[76], stage1_8[77], stage1_8[78]},
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage2_12[5],stage2_11[12],stage2_10[18],stage2_9[19],stage2_8[23]}
   );
   gpc606_5 gpc365 (
      {stage1_8[79], stage1_8[80], stage1_8[81], stage1_8[82], stage1_8[83], stage1_8[84]},
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage2_12[6],stage2_11[13],stage2_10[19],stage2_9[20],stage2_8[24]}
   );
   gpc606_5 gpc366 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[7],stage2_11[14],stage2_10[20],stage2_9[21]}
   );
   gpc606_5 gpc367 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[8],stage2_11[15],stage2_10[21],stage2_9[22]}
   );
   gpc615_5 gpc368 (
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46]},
      {stage1_11[12]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[2],stage2_12[9],stage2_11[16],stage2_10[22]}
   );
   gpc615_5 gpc369 (
      {stage1_10[47], stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51]},
      {stage1_11[13]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[3],stage2_12[10],stage2_11[17],stage2_10[23]}
   );
   gpc615_5 gpc370 (
      {stage1_10[52], stage1_10[53], stage1_10[54], stage1_10[55], stage1_10[56]},
      {stage1_11[14]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[4],stage2_12[11],stage2_11[18],stage2_10[24]}
   );
   gpc615_5 gpc371 (
      {stage1_10[57], stage1_10[58], stage1_10[59], stage1_10[60], 1'b0},
      {stage1_11[15]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[5],stage2_12[12],stage2_11[19],stage2_10[25]}
   );
   gpc1343_5 gpc372 (
      {stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27]},
      {stage1_13[0], stage1_13[1], stage1_13[2]},
      {stage1_14[0]},
      {stage2_15[0],stage2_14[4],stage2_13[6],stage2_12[13],stage2_11[20]}
   );
   gpc615_5 gpc373 (
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage1_12[28]},
      {stage1_13[3], stage1_13[4], stage1_13[5], stage1_13[6], stage1_13[7], stage1_13[8]},
      {stage2_15[1],stage2_14[5],stage2_13[7],stage2_12[14],stage2_11[21]}
   );
   gpc615_5 gpc374 (
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28]},
      {stage1_12[29]},
      {stage1_13[9], stage1_13[10], stage1_13[11], stage1_13[12], stage1_13[13], stage1_13[14]},
      {stage2_15[2],stage2_14[6],stage2_13[8],stage2_12[15],stage2_11[22]}
   );
   gpc615_5 gpc375 (
      {stage1_11[29], stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33]},
      {stage1_12[30]},
      {stage1_13[15], stage1_13[16], stage1_13[17], stage1_13[18], stage1_13[19], stage1_13[20]},
      {stage2_15[3],stage2_14[7],stage2_13[9],stage2_12[16],stage2_11[23]}
   );
   gpc615_5 gpc376 (
      {stage1_11[34], stage1_11[35], stage1_11[36], stage1_11[37], stage1_11[38]},
      {stage1_12[31]},
      {stage1_13[21], stage1_13[22], stage1_13[23], stage1_13[24], stage1_13[25], stage1_13[26]},
      {stage2_15[4],stage2_14[8],stage2_13[10],stage2_12[17],stage2_11[24]}
   );
   gpc615_5 gpc377 (
      {stage1_11[39], stage1_11[40], stage1_11[41], stage1_11[42], stage1_11[43]},
      {stage1_12[32]},
      {stage1_13[27], stage1_13[28], stage1_13[29], stage1_13[30], stage1_13[31], stage1_13[32]},
      {stage2_15[5],stage2_14[9],stage2_13[11],stage2_12[18],stage2_11[25]}
   );
   gpc615_5 gpc378 (
      {stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48]},
      {stage1_12[33]},
      {stage1_13[33], stage1_13[34], stage1_13[35], stage1_13[36], stage1_13[37], stage1_13[38]},
      {stage2_15[6],stage2_14[10],stage2_13[12],stage2_12[19],stage2_11[26]}
   );
   gpc615_5 gpc379 (
      {stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage1_12[34]},
      {stage1_13[39], stage1_13[40], stage1_13[41], stage1_13[42], stage1_13[43], stage1_13[44]},
      {stage2_15[7],stage2_14[11],stage2_13[13],stage2_12[20],stage2_11[27]}
   );
   gpc615_5 gpc380 (
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], 1'b0},
      {stage1_12[35]},
      {stage1_13[45], stage1_13[46], stage1_13[47], stage1_13[48], stage1_13[49], stage1_13[50]},
      {stage2_15[8],stage2_14[12],stage2_13[14],stage2_12[21],stage2_11[28]}
   );
   gpc606_5 gpc381 (
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6]},
      {stage2_16[0],stage2_15[9],stage2_14[13],stage2_13[15],stage2_12[22]}
   );
   gpc606_5 gpc382 (
      {stage1_12[42], stage1_12[43], stage1_12[44], stage1_12[45], stage1_12[46], stage1_12[47]},
      {stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12]},
      {stage2_16[1],stage2_15[10],stage2_14[14],stage2_13[16],stage2_12[23]}
   );
   gpc606_5 gpc383 (
      {stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52], stage1_12[53]},
      {stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17], stage1_14[18]},
      {stage2_16[2],stage2_15[11],stage2_14[15],stage2_13[17],stage2_12[24]}
   );
   gpc606_5 gpc384 (
      {stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], stage1_12[58], stage1_12[59]},
      {stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22], stage1_14[23], stage1_14[24]},
      {stage2_16[3],stage2_15[12],stage2_14[16],stage2_13[18],stage2_12[25]}
   );
   gpc606_5 gpc385 (
      {stage1_12[60], stage1_12[61], stage1_12[62], stage1_12[63], stage1_12[64], stage1_12[65]},
      {stage1_14[25], stage1_14[26], stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30]},
      {stage2_16[4],stage2_15[13],stage2_14[17],stage2_13[19],stage2_12[26]}
   );
   gpc606_5 gpc386 (
      {stage1_13[51], stage1_13[52], stage1_13[53], stage1_13[54], stage1_13[55], stage1_13[56]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[5],stage2_15[14],stage2_14[18],stage2_13[20]}
   );
   gpc606_5 gpc387 (
      {stage1_13[57], stage1_13[58], stage1_13[59], stage1_13[60], stage1_13[61], stage1_13[62]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[6],stage2_15[15],stage2_14[19],stage2_13[21]}
   );
   gpc606_5 gpc388 (
      {stage1_13[63], stage1_13[64], stage1_13[65], stage1_13[66], stage1_13[67], stage1_13[68]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[7],stage2_15[16],stage2_14[20],stage2_13[22]}
   );
   gpc606_5 gpc389 (
      {stage1_13[69], stage1_13[70], stage1_13[71], stage1_13[72], stage1_13[73], stage1_13[74]},
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage2_17[3],stage2_16[8],stage2_15[17],stage2_14[21],stage2_13[23]}
   );
   gpc606_5 gpc390 (
      {stage1_14[31], stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[4],stage2_16[9],stage2_15[18],stage2_14[22]}
   );
   gpc606_5 gpc391 (
      {stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41], stage1_14[42]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[5],stage2_16[10],stage2_15[19],stage2_14[23]}
   );
   gpc606_5 gpc392 (
      {stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47], stage1_14[48]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[6],stage2_16[11],stage2_15[20],stage2_14[24]}
   );
   gpc606_5 gpc393 (
      {stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52], stage1_14[53], stage1_14[54]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[7],stage2_16[12],stage2_15[21],stage2_14[25]}
   );
   gpc606_5 gpc394 (
      {stage1_14[55], stage1_14[56], stage1_14[57], stage1_14[58], stage1_14[59], stage1_14[60]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[8],stage2_16[13],stage2_15[22],stage2_14[26]}
   );
   gpc606_5 gpc395 (
      {stage1_14[61], stage1_14[62], stage1_14[63], stage1_14[64], stage1_14[65], stage1_14[66]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[9],stage2_16[14],stage2_15[23],stage2_14[27]}
   );
   gpc606_5 gpc396 (
      {stage1_14[67], stage1_14[68], stage1_14[69], stage1_14[70], stage1_14[71], stage1_14[72]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[10],stage2_16[15],stage2_15[24],stage2_14[28]}
   );
   gpc615_5 gpc397 (
      {stage1_14[73], stage1_14[74], stage1_14[75], stage1_14[76], stage1_14[77]},
      {stage1_15[24]},
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage2_18[7],stage2_17[11],stage2_16[16],stage2_15[25],stage2_14[29]}
   );
   gpc615_5 gpc398 (
      {stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage1_16[48]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[8],stage2_17[12],stage2_16[17],stage2_15[26]}
   );
   gpc1_1 gpc399 (
      {stage1_0[27]},
      {stage2_0[5]}
   );
   gpc1_1 gpc400 (
      {stage1_0[28]},
      {stage2_0[6]}
   );
   gpc1_1 gpc401 (
      {stage1_0[29]},
      {stage2_0[7]}
   );
   gpc1_1 gpc402 (
      {stage1_0[30]},
      {stage2_0[8]}
   );
   gpc1_1 gpc403 (
      {stage1_0[31]},
      {stage2_0[9]}
   );
   gpc1_1 gpc404 (
      {stage1_0[32]},
      {stage2_0[10]}
   );
   gpc1_1 gpc405 (
      {stage1_1[27]},
      {stage2_1[9]}
   );
   gpc1_1 gpc406 (
      {stage1_1[28]},
      {stage2_1[10]}
   );
   gpc1_1 gpc407 (
      {stage1_1[29]},
      {stage2_1[11]}
   );
   gpc1_1 gpc408 (
      {stage1_1[30]},
      {stage2_1[12]}
   );
   gpc1_1 gpc409 (
      {stage1_1[31]},
      {stage2_1[13]}
   );
   gpc1_1 gpc410 (
      {stage1_1[32]},
      {stage2_1[14]}
   );
   gpc1_1 gpc411 (
      {stage1_1[33]},
      {stage2_1[15]}
   );
   gpc1_1 gpc412 (
      {stage1_1[34]},
      {stage2_1[16]}
   );
   gpc1_1 gpc413 (
      {stage1_1[35]},
      {stage2_1[17]}
   );
   gpc1_1 gpc414 (
      {stage1_1[36]},
      {stage2_1[18]}
   );
   gpc1_1 gpc415 (
      {stage1_1[37]},
      {stage2_1[19]}
   );
   gpc1_1 gpc416 (
      {stage1_1[38]},
      {stage2_1[20]}
   );
   gpc1_1 gpc417 (
      {stage1_1[39]},
      {stage2_1[21]}
   );
   gpc1_1 gpc418 (
      {stage1_1[40]},
      {stage2_1[22]}
   );
   gpc1_1 gpc419 (
      {stage1_1[41]},
      {stage2_1[23]}
   );
   gpc1_1 gpc420 (
      {stage1_1[42]},
      {stage2_1[24]}
   );
   gpc1_1 gpc421 (
      {stage1_1[43]},
      {stage2_1[25]}
   );
   gpc1_1 gpc422 (
      {stage1_1[44]},
      {stage2_1[26]}
   );
   gpc1_1 gpc423 (
      {stage1_1[45]},
      {stage2_1[27]}
   );
   gpc1_1 gpc424 (
      {stage1_1[46]},
      {stage2_1[28]}
   );
   gpc1_1 gpc425 (
      {stage1_1[47]},
      {stage2_1[29]}
   );
   gpc1_1 gpc426 (
      {stage1_3[81]},
      {stage2_3[26]}
   );
   gpc1_1 gpc427 (
      {stage1_3[82]},
      {stage2_3[27]}
   );
   gpc1_1 gpc428 (
      {stage1_3[83]},
      {stage2_3[28]}
   );
   gpc1_1 gpc429 (
      {stage1_3[84]},
      {stage2_3[29]}
   );
   gpc1_1 gpc430 (
      {stage1_3[85]},
      {stage2_3[30]}
   );
   gpc1_1 gpc431 (
      {stage1_3[86]},
      {stage2_3[31]}
   );
   gpc1_1 gpc432 (
      {stage1_3[87]},
      {stage2_3[32]}
   );
   gpc1_1 gpc433 (
      {stage1_3[88]},
      {stage2_3[33]}
   );
   gpc1_1 gpc434 (
      {stage1_3[89]},
      {stage2_3[34]}
   );
   gpc1_1 gpc435 (
      {stage1_3[90]},
      {stage2_3[35]}
   );
   gpc1_1 gpc436 (
      {stage1_3[91]},
      {stage2_3[36]}
   );
   gpc1_1 gpc437 (
      {stage1_5[67]},
      {stage2_5[26]}
   );
   gpc1_1 gpc438 (
      {stage1_5[68]},
      {stage2_5[27]}
   );
   gpc1_1 gpc439 (
      {stage1_5[69]},
      {stage2_5[28]}
   );
   gpc1_1 gpc440 (
      {stage1_5[70]},
      {stage2_5[29]}
   );
   gpc1_1 gpc441 (
      {stage1_6[58]},
      {stage2_6[28]}
   );
   gpc1_1 gpc442 (
      {stage1_6[59]},
      {stage2_6[29]}
   );
   gpc1_1 gpc443 (
      {stage1_7[43]},
      {stage2_7[28]}
   );
   gpc1_1 gpc444 (
      {stage1_7[44]},
      {stage2_7[29]}
   );
   gpc1_1 gpc445 (
      {stage1_7[45]},
      {stage2_7[30]}
   );
   gpc1_1 gpc446 (
      {stage1_7[46]},
      {stage2_7[31]}
   );
   gpc1_1 gpc447 (
      {stage1_7[47]},
      {stage2_7[32]}
   );
   gpc1_1 gpc448 (
      {stage1_7[48]},
      {stage2_7[33]}
   );
   gpc1_1 gpc449 (
      {stage1_7[49]},
      {stage2_7[34]}
   );
   gpc1_1 gpc450 (
      {stage1_7[50]},
      {stage2_7[35]}
   );
   gpc1_1 gpc451 (
      {stage1_7[51]},
      {stage2_7[36]}
   );
   gpc1_1 gpc452 (
      {stage1_7[52]},
      {stage2_7[37]}
   );
   gpc1_1 gpc453 (
      {stage1_7[53]},
      {stage2_7[38]}
   );
   gpc1_1 gpc454 (
      {stage1_8[85]},
      {stage2_8[25]}
   );
   gpc1_1 gpc455 (
      {stage1_8[86]},
      {stage2_8[26]}
   );
   gpc1_1 gpc456 (
      {stage1_8[87]},
      {stage2_8[27]}
   );
   gpc1_1 gpc457 (
      {stage1_8[88]},
      {stage2_8[28]}
   );
   gpc1_1 gpc458 (
      {stage1_8[89]},
      {stage2_8[29]}
   );
   gpc1_1 gpc459 (
      {stage1_9[54]},
      {stage2_9[23]}
   );
   gpc1_1 gpc460 (
      {stage1_9[55]},
      {stage2_9[24]}
   );
   gpc1_1 gpc461 (
      {stage1_9[56]},
      {stage2_9[25]}
   );
   gpc1_1 gpc462 (
      {stage1_9[57]},
      {stage2_9[26]}
   );
   gpc1_1 gpc463 (
      {stage1_9[58]},
      {stage2_9[27]}
   );
   gpc1_1 gpc464 (
      {stage1_9[59]},
      {stage2_9[28]}
   );
   gpc1_1 gpc465 (
      {stage1_9[60]},
      {stage2_9[29]}
   );
   gpc1_1 gpc466 (
      {stage1_9[61]},
      {stage2_9[30]}
   );
   gpc1_1 gpc467 (
      {stage1_9[62]},
      {stage2_9[31]}
   );
   gpc1_1 gpc468 (
      {stage1_9[63]},
      {stage2_9[32]}
   );
   gpc1_1 gpc469 (
      {stage1_9[64]},
      {stage2_9[33]}
   );
   gpc1_1 gpc470 (
      {stage1_9[65]},
      {stage2_9[34]}
   );
   gpc1_1 gpc471 (
      {stage1_9[66]},
      {stage2_9[35]}
   );
   gpc1_1 gpc472 (
      {stage1_9[67]},
      {stage2_9[36]}
   );
   gpc1_1 gpc473 (
      {stage1_9[68]},
      {stage2_9[37]}
   );
   gpc1_1 gpc474 (
      {stage1_9[69]},
      {stage2_9[38]}
   );
   gpc1_1 gpc475 (
      {stage1_9[70]},
      {stage2_9[39]}
   );
   gpc1_1 gpc476 (
      {stage1_9[71]},
      {stage2_9[40]}
   );
   gpc1_1 gpc477 (
      {stage1_9[72]},
      {stage2_9[41]}
   );
   gpc1_1 gpc478 (
      {stage1_9[73]},
      {stage2_9[42]}
   );
   gpc1_1 gpc479 (
      {stage1_9[74]},
      {stage2_9[43]}
   );
   gpc1_1 gpc480 (
      {stage1_9[75]},
      {stage2_9[44]}
   );
   gpc1_1 gpc481 (
      {stage1_9[76]},
      {stage2_9[45]}
   );
   gpc1_1 gpc482 (
      {stage1_9[77]},
      {stage2_9[46]}
   );
   gpc1_1 gpc483 (
      {stage1_9[78]},
      {stage2_9[47]}
   );
   gpc1_1 gpc484 (
      {stage1_9[79]},
      {stage2_9[48]}
   );
   gpc1_1 gpc485 (
      {stage1_9[80]},
      {stage2_9[49]}
   );
   gpc1_1 gpc486 (
      {stage1_9[81]},
      {stage2_9[50]}
   );
   gpc1_1 gpc487 (
      {stage1_9[82]},
      {stage2_9[51]}
   );
   gpc1_1 gpc488 (
      {stage1_12[66]},
      {stage2_12[27]}
   );
   gpc1_1 gpc489 (
      {stage1_12[67]},
      {stage2_12[28]}
   );
   gpc1_1 gpc490 (
      {stage1_12[68]},
      {stage2_12[29]}
   );
   gpc1_1 gpc491 (
      {stage1_12[69]},
      {stage2_12[30]}
   );
   gpc1_1 gpc492 (
      {stage1_12[70]},
      {stage2_12[31]}
   );
   gpc1_1 gpc493 (
      {stage1_12[71]},
      {stage2_12[32]}
   );
   gpc1_1 gpc494 (
      {stage1_12[72]},
      {stage2_12[33]}
   );
   gpc1_1 gpc495 (
      {stage1_13[75]},
      {stage2_13[24]}
   );
   gpc1_1 gpc496 (
      {stage1_13[76]},
      {stage2_13[25]}
   );
   gpc1_1 gpc497 (
      {stage1_13[77]},
      {stage2_13[26]}
   );
   gpc1_1 gpc498 (
      {stage1_15[30]},
      {stage2_15[27]}
   );
   gpc1_1 gpc499 (
      {stage1_15[31]},
      {stage2_15[28]}
   );
   gpc1_1 gpc500 (
      {stage1_15[32]},
      {stage2_15[29]}
   );
   gpc1_1 gpc501 (
      {stage1_15[33]},
      {stage2_15[30]}
   );
   gpc1_1 gpc502 (
      {stage1_15[34]},
      {stage2_15[31]}
   );
   gpc1_1 gpc503 (
      {stage1_15[35]},
      {stage2_15[32]}
   );
   gpc1_1 gpc504 (
      {stage1_15[36]},
      {stage2_15[33]}
   );
   gpc1_1 gpc505 (
      {stage1_15[37]},
      {stage2_15[34]}
   );
   gpc1_1 gpc506 (
      {stage1_15[38]},
      {stage2_15[35]}
   );
   gpc1_1 gpc507 (
      {stage1_15[39]},
      {stage2_15[36]}
   );
   gpc1_1 gpc508 (
      {stage1_15[40]},
      {stage2_15[37]}
   );
   gpc1_1 gpc509 (
      {stage1_15[41]},
      {stage2_15[38]}
   );
   gpc1_1 gpc510 (
      {stage1_15[42]},
      {stage2_15[39]}
   );
   gpc1_1 gpc511 (
      {stage1_15[43]},
      {stage2_15[40]}
   );
   gpc1_1 gpc512 (
      {stage1_15[44]},
      {stage2_15[41]}
   );
   gpc1_1 gpc513 (
      {stage1_15[45]},
      {stage2_15[42]}
   );
   gpc1_1 gpc514 (
      {stage1_15[46]},
      {stage2_15[43]}
   );
   gpc1_1 gpc515 (
      {stage1_15[47]},
      {stage2_15[44]}
   );
   gpc1_1 gpc516 (
      {stage1_15[48]},
      {stage2_15[45]}
   );
   gpc1_1 gpc517 (
      {stage1_15[49]},
      {stage2_15[46]}
   );
   gpc1_1 gpc518 (
      {stage1_15[50]},
      {stage2_15[47]}
   );
   gpc1_1 gpc519 (
      {stage1_15[51]},
      {stage2_15[48]}
   );
   gpc1_1 gpc520 (
      {stage1_15[52]},
      {stage2_15[49]}
   );
   gpc1_1 gpc521 (
      {stage1_15[53]},
      {stage2_15[50]}
   );
   gpc1_1 gpc522 (
      {stage1_17[6]},
      {stage2_17[13]}
   );
   gpc1_1 gpc523 (
      {stage1_17[7]},
      {stage2_17[14]}
   );
   gpc1_1 gpc524 (
      {stage1_17[8]},
      {stage2_17[15]}
   );
   gpc1_1 gpc525 (
      {stage1_17[9]},
      {stage2_17[16]}
   );
   gpc1_1 gpc526 (
      {stage1_17[10]},
      {stage2_17[17]}
   );
   gpc1_1 gpc527 (
      {stage1_17[11]},
      {stage2_17[18]}
   );
   gpc1_1 gpc528 (
      {stage1_17[12]},
      {stage2_17[19]}
   );
   gpc1_1 gpc529 (
      {stage1_17[13]},
      {stage2_17[20]}
   );
   gpc1_1 gpc530 (
      {stage1_17[14]},
      {stage2_17[21]}
   );
   gpc1_1 gpc531 (
      {stage1_17[15]},
      {stage2_17[22]}
   );
   gpc1_1 gpc532 (
      {stage1_17[16]},
      {stage2_17[23]}
   );
   gpc1_1 gpc533 (
      {stage1_17[17]},
      {stage2_17[24]}
   );
   gpc1_1 gpc534 (
      {stage1_17[18]},
      {stage2_17[25]}
   );
   gpc1_1 gpc535 (
      {stage1_17[19]},
      {stage2_17[26]}
   );
   gpc1_1 gpc536 (
      {stage1_17[20]},
      {stage2_17[27]}
   );
   gpc1_1 gpc537 (
      {stage1_17[21]},
      {stage2_17[28]}
   );
   gpc1_1 gpc538 (
      {stage1_17[22]},
      {stage2_17[29]}
   );
   gpc1_1 gpc539 (
      {stage1_17[23]},
      {stage2_17[30]}
   );
   gpc1_1 gpc540 (
      {stage1_17[24]},
      {stage2_17[31]}
   );
   gpc1_1 gpc541 (
      {stage1_17[25]},
      {stage2_17[32]}
   );
   gpc1_1 gpc542 (
      {stage1_17[26]},
      {stage2_17[33]}
   );
   gpc1_1 gpc543 (
      {stage1_17[27]},
      {stage2_17[34]}
   );
   gpc1163_5 gpc544 (
      {stage2_0[0], stage2_0[1], stage2_0[2]},
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[0]},
      {stage2_3[0]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc1163_5 gpc545 (
      {stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[1]},
      {stage2_3[1]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc606_5 gpc546 (
      {stage2_1[12], stage2_1[13], stage2_1[14], stage2_1[15], stage2_1[16], stage2_1[17]},
      {stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7]},
      {stage3_5[0],stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2]}
   );
   gpc606_5 gpc547 (
      {stage2_1[18], stage2_1[19], stage2_1[20], stage2_1[21], stage2_1[22], stage2_1[23]},
      {stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12], stage2_3[13]},
      {stage3_5[1],stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3]}
   );
   gpc606_5 gpc548 (
      {stage2_1[24], stage2_1[25], stage2_1[26], stage2_1[27], stage2_1[28], stage2_1[29]},
      {stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18], stage2_3[19]},
      {stage3_5[2],stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4]}
   );
   gpc615_5 gpc549 (
      {stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23], stage2_3[24]},
      {stage2_4[0]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[0],stage3_5[3],stage3_4[5],stage3_3[5]}
   );
   gpc615_5 gpc550 (
      {stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28], stage2_3[29]},
      {stage2_4[1]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[1],stage3_5[4],stage3_4[6],stage3_3[6]}
   );
   gpc606_5 gpc551 (
      {stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5], stage2_4[6], stage2_4[7]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[2],stage3_6[2],stage3_5[5],stage3_4[7]}
   );
   gpc606_5 gpc552 (
      {stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11], stage2_4[12], stage2_4[13]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[3],stage3_6[3],stage3_5[6],stage3_4[8]}
   );
   gpc606_5 gpc553 (
      {stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17], stage2_4[18], stage2_4[19]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[4],stage3_6[4],stage3_5[7],stage3_4[9]}
   );
   gpc606_5 gpc554 (
      {stage2_4[20], stage2_4[21], stage2_4[22], stage2_4[23], stage2_4[24], stage2_4[25]},
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage3_8[3],stage3_7[5],stage3_6[5],stage3_5[8],stage3_4[10]}
   );
   gpc606_5 gpc555 (
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[4],stage3_7[6],stage3_6[6],stage3_5[9]}
   );
   gpc606_5 gpc556 (
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[5],stage3_7[7],stage3_6[7],stage3_5[10]}
   );
   gpc606_5 gpc557 (
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17]},
      {stage3_9[2],stage3_8[6],stage3_7[8],stage3_6[8],stage3_5[11]}
   );
   gpc615_5 gpc558 (
      {stage2_6[24], stage2_6[25], stage2_6[26], stage2_6[27], stage2_6[28]},
      {stage2_7[18]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[3],stage3_8[7],stage3_7[9],stage3_6[9]}
   );
   gpc615_5 gpc559 (
      {stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23]},
      {stage2_8[6]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[1],stage3_9[4],stage3_8[8],stage3_7[10]}
   );
   gpc615_5 gpc560 (
      {stage2_7[24], stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28]},
      {stage2_8[7]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[2],stage3_9[5],stage3_8[9],stage3_7[11]}
   );
   gpc615_5 gpc561 (
      {stage2_7[29], stage2_7[30], stage2_7[31], stage2_7[32], stage2_7[33]},
      {stage2_8[8]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[3],stage3_9[6],stage3_8[10],stage3_7[12]}
   );
   gpc615_5 gpc562 (
      {stage2_7[34], stage2_7[35], stage2_7[36], stage2_7[37], stage2_7[38]},
      {stage2_8[9]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[4],stage3_9[7],stage3_8[11],stage3_7[13]}
   );
   gpc606_5 gpc563 (
      {stage2_8[10], stage2_8[11], stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[4],stage3_10[5],stage3_9[8],stage3_8[12]}
   );
   gpc606_5 gpc564 (
      {stage2_8[16], stage2_8[17], stage2_8[18], stage2_8[19], stage2_8[20], stage2_8[21]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[5],stage3_10[6],stage3_9[9],stage3_8[13]}
   );
   gpc606_5 gpc565 (
      {stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25], stage2_8[26], stage2_8[27]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[6],stage3_10[7],stage3_9[10],stage3_8[14]}
   );
   gpc606_5 gpc566 (
      {stage2_9[24], stage2_9[25], stage2_9[26], stage2_9[27], stage2_9[28], stage2_9[29]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[3],stage3_11[7],stage3_10[8],stage3_9[11]}
   );
   gpc606_5 gpc567 (
      {stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34], stage2_9[35]},
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage3_13[1],stage3_12[4],stage3_11[8],stage3_10[9],stage3_9[12]}
   );
   gpc606_5 gpc568 (
      {stage2_9[36], stage2_9[37], stage2_9[38], stage2_9[39], stage2_9[40], stage2_9[41]},
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16], stage2_11[17]},
      {stage3_13[2],stage3_12[5],stage3_11[9],stage3_10[10],stage3_9[13]}
   );
   gpc615_5 gpc569 (
      {stage2_9[42], stage2_9[43], stage2_9[44], stage2_9[45], stage2_9[46]},
      {stage2_10[18]},
      {stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23]},
      {stage3_13[3],stage3_12[6],stage3_11[10],stage3_10[11],stage3_9[14]}
   );
   gpc615_5 gpc570 (
      {stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage2_11[24]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[4],stage3_12[7],stage3_11[11],stage3_10[12]}
   );
   gpc615_5 gpc571 (
      {stage2_11[25], stage2_11[26], stage2_11[27], stage2_11[28], 1'b0},
      {stage2_12[6]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[1],stage3_13[5],stage3_12[8],stage3_11[12]}
   );
   gpc606_5 gpc572 (
      {stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[1],stage3_14[2],stage3_13[6],stage3_12[9]}
   );
   gpc606_5 gpc573 (
      {stage2_12[13], stage2_12[14], stage2_12[15], stage2_12[16], stage2_12[17], stage2_12[18]},
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage3_16[1],stage3_15[2],stage3_14[3],stage3_13[7],stage3_12[10]}
   );
   gpc606_5 gpc574 (
      {stage2_12[19], stage2_12[20], stage2_12[21], stage2_12[22], stage2_12[23], stage2_12[24]},
      {stage2_14[12], stage2_14[13], stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17]},
      {stage3_16[2],stage3_15[3],stage3_14[4],stage3_13[8],stage3_12[11]}
   );
   gpc606_5 gpc575 (
      {stage2_12[25], stage2_12[26], stage2_12[27], stage2_12[28], stage2_12[29], stage2_12[30]},
      {stage2_14[18], stage2_14[19], stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23]},
      {stage3_16[3],stage3_15[4],stage3_14[5],stage3_13[9],stage3_12[12]}
   );
   gpc606_5 gpc576 (
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5]},
      {stage3_17[0],stage3_16[4],stage3_15[5],stage3_14[6],stage3_13[10]}
   );
   gpc606_5 gpc577 (
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11]},
      {stage3_17[1],stage3_16[5],stage3_15[6],stage3_14[7],stage3_13[11]}
   );
   gpc606_5 gpc578 (
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage2_15[12], stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage3_17[2],stage3_16[6],stage3_15[7],stage3_14[8],stage3_13[12]}
   );
   gpc606_5 gpc579 (
      {stage2_14[24], stage2_14[25], stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[3],stage3_16[7],stage3_15[8],stage3_14[9]}
   );
   gpc615_5 gpc580 (
      {stage2_15[18], stage2_15[19], stage2_15[20], stage2_15[21], stage2_15[22]},
      {stage2_16[6]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[1],stage3_17[4],stage3_16[8],stage3_15[9]}
   );
   gpc615_5 gpc581 (
      {stage2_15[23], stage2_15[24], stage2_15[25], stage2_15[26], stage2_15[27]},
      {stage2_16[7]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[2],stage3_17[5],stage3_16[9],stage3_15[10]}
   );
   gpc615_5 gpc582 (
      {stage2_15[28], stage2_15[29], stage2_15[30], stage2_15[31], stage2_15[32]},
      {stage2_16[8]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[3],stage3_17[6],stage3_16[10],stage3_15[11]}
   );
   gpc615_5 gpc583 (
      {stage2_15[33], stage2_15[34], stage2_15[35], stage2_15[36], stage2_15[37]},
      {stage2_16[9]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[4],stage3_17[7],stage3_16[11],stage3_15[12]}
   );
   gpc615_5 gpc584 (
      {stage2_15[38], stage2_15[39], stage2_15[40], stage2_15[41], stage2_15[42]},
      {stage2_16[10]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[5],stage3_17[8],stage3_16[12],stage3_15[13]}
   );
   gpc615_5 gpc585 (
      {stage2_15[43], stage2_15[44], stage2_15[45], stage2_15[46], stage2_15[47]},
      {stage2_16[11]},
      {stage2_17[30], stage2_17[31], stage2_17[32], stage2_17[33], stage2_17[34], 1'b0},
      {stage3_19[5],stage3_18[6],stage3_17[9],stage3_16[13],stage3_15[14]}
   );
   gpc606_5 gpc586 (
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5]},
      {stage3_20[0],stage3_19[6],stage3_18[7],stage3_17[10],stage3_16[14]}
   );
   gpc1_1 gpc587 (
      {stage2_0[6]},
      {stage3_0[2]}
   );
   gpc1_1 gpc588 (
      {stage2_0[7]},
      {stage3_0[3]}
   );
   gpc1_1 gpc589 (
      {stage2_0[8]},
      {stage3_0[4]}
   );
   gpc1_1 gpc590 (
      {stage2_0[9]},
      {stage3_0[5]}
   );
   gpc1_1 gpc591 (
      {stage2_0[10]},
      {stage3_0[6]}
   );
   gpc1_1 gpc592 (
      {stage2_2[2]},
      {stage3_2[5]}
   );
   gpc1_1 gpc593 (
      {stage2_2[3]},
      {stage3_2[6]}
   );
   gpc1_1 gpc594 (
      {stage2_2[4]},
      {stage3_2[7]}
   );
   gpc1_1 gpc595 (
      {stage2_2[5]},
      {stage3_2[8]}
   );
   gpc1_1 gpc596 (
      {stage2_2[6]},
      {stage3_2[9]}
   );
   gpc1_1 gpc597 (
      {stage2_2[7]},
      {stage3_2[10]}
   );
   gpc1_1 gpc598 (
      {stage2_2[8]},
      {stage3_2[11]}
   );
   gpc1_1 gpc599 (
      {stage2_2[9]},
      {stage3_2[12]}
   );
   gpc1_1 gpc600 (
      {stage2_2[10]},
      {stage3_2[13]}
   );
   gpc1_1 gpc601 (
      {stage2_2[11]},
      {stage3_2[14]}
   );
   gpc1_1 gpc602 (
      {stage2_2[12]},
      {stage3_2[15]}
   );
   gpc1_1 gpc603 (
      {stage2_2[13]},
      {stage3_2[16]}
   );
   gpc1_1 gpc604 (
      {stage2_2[14]},
      {stage3_2[17]}
   );
   gpc1_1 gpc605 (
      {stage2_2[15]},
      {stage3_2[18]}
   );
   gpc1_1 gpc606 (
      {stage2_3[30]},
      {stage3_3[7]}
   );
   gpc1_1 gpc607 (
      {stage2_3[31]},
      {stage3_3[8]}
   );
   gpc1_1 gpc608 (
      {stage2_3[32]},
      {stage3_3[9]}
   );
   gpc1_1 gpc609 (
      {stage2_3[33]},
      {stage3_3[10]}
   );
   gpc1_1 gpc610 (
      {stage2_3[34]},
      {stage3_3[11]}
   );
   gpc1_1 gpc611 (
      {stage2_3[35]},
      {stage3_3[12]}
   );
   gpc1_1 gpc612 (
      {stage2_3[36]},
      {stage3_3[13]}
   );
   gpc1_1 gpc613 (
      {stage2_4[26]},
      {stage3_4[11]}
   );
   gpc1_1 gpc614 (
      {stage2_4[27]},
      {stage3_4[12]}
   );
   gpc1_1 gpc615 (
      {stage2_4[28]},
      {stage3_4[13]}
   );
   gpc1_1 gpc616 (
      {stage2_4[29]},
      {stage3_4[14]}
   );
   gpc1_1 gpc617 (
      {stage2_6[29]},
      {stage3_6[10]}
   );
   gpc1_1 gpc618 (
      {stage2_8[28]},
      {stage3_8[15]}
   );
   gpc1_1 gpc619 (
      {stage2_8[29]},
      {stage3_8[16]}
   );
   gpc1_1 gpc620 (
      {stage2_9[47]},
      {stage3_9[15]}
   );
   gpc1_1 gpc621 (
      {stage2_9[48]},
      {stage3_9[16]}
   );
   gpc1_1 gpc622 (
      {stage2_9[49]},
      {stage3_9[17]}
   );
   gpc1_1 gpc623 (
      {stage2_9[50]},
      {stage3_9[18]}
   );
   gpc1_1 gpc624 (
      {stage2_9[51]},
      {stage3_9[19]}
   );
   gpc1_1 gpc625 (
      {stage2_10[24]},
      {stage3_10[13]}
   );
   gpc1_1 gpc626 (
      {stage2_10[25]},
      {stage3_10[14]}
   );
   gpc1_1 gpc627 (
      {stage2_12[31]},
      {stage3_12[13]}
   );
   gpc1_1 gpc628 (
      {stage2_12[32]},
      {stage3_12[14]}
   );
   gpc1_1 gpc629 (
      {stage2_12[33]},
      {stage3_12[15]}
   );
   gpc1_1 gpc630 (
      {stage2_13[24]},
      {stage3_13[13]}
   );
   gpc1_1 gpc631 (
      {stage2_13[25]},
      {stage3_13[14]}
   );
   gpc1_1 gpc632 (
      {stage2_13[26]},
      {stage3_13[15]}
   );
   gpc1_1 gpc633 (
      {stage2_15[48]},
      {stage3_15[15]}
   );
   gpc1_1 gpc634 (
      {stage2_15[49]},
      {stage3_15[16]}
   );
   gpc1_1 gpc635 (
      {stage2_15[50]},
      {stage3_15[17]}
   );
   gpc1_1 gpc636 (
      {stage2_18[6]},
      {stage3_18[8]}
   );
   gpc1_1 gpc637 (
      {stage2_18[7]},
      {stage3_18[9]}
   );
   gpc1_1 gpc638 (
      {stage2_18[8]},
      {stage3_18[10]}
   );
   gpc1_1 gpc639 (
      {stage2_19[0]},
      {stage3_19[7]}
   );
   gpc615_5 gpc640 (
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4]},
      {stage3_3[0]},
      {stage3_4[0], stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0]}
   );
   gpc615_5 gpc641 (
      {stage3_2[5], stage3_2[6], stage3_2[7], stage3_2[8], stage3_2[9]},
      {stage3_3[1]},
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10], stage3_4[11]},
      {stage4_6[1],stage4_5[1],stage4_4[1],stage4_3[1],stage4_2[1]}
   );
   gpc615_5 gpc642 (
      {stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5], stage3_3[6]},
      {stage3_4[12]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[2],stage4_5[2],stage4_4[2],stage4_3[2]}
   );
   gpc615_5 gpc643 (
      {stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage3_4[13]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[3],stage4_5[3],stage4_4[3],stage4_3[3]}
   );
   gpc615_5 gpc644 (
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4]},
      {stage3_7[0]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[0],stage4_7[2],stage4_6[4]}
   );
   gpc615_5 gpc645 (
      {stage3_6[5], stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9]},
      {stage3_7[1]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[1],stage4_9[1],stage4_8[1],stage4_7[3],stage4_6[5]}
   );
   gpc615_5 gpc646 (
      {stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5], stage3_7[6]},
      {stage3_8[12]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[2],stage4_9[2],stage4_8[2],stage4_7[4]}
   );
   gpc615_5 gpc647 (
      {stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10], stage3_7[11]},
      {stage3_8[13]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[3],stage4_9[3],stage4_8[3],stage4_7[5]}
   );
   gpc606_5 gpc648 (
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[0],stage4_11[2],stage4_10[4],stage4_9[4]}
   );
   gpc606_5 gpc649 (
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5]},
      {stage4_14[0],stage4_13[1],stage4_12[1],stage4_11[3],stage4_10[5]}
   );
   gpc606_5 gpc650 (
      {stage3_10[6], stage3_10[7], stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11]},
      {stage4_14[1],stage4_13[2],stage4_12[2],stage4_11[4],stage4_10[6]}
   );
   gpc1406_5 gpc651 (
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3]},
      {stage3_16[0]},
      {stage4_17[0],stage4_16[0],stage4_15[0],stage4_14[2],stage4_13[3]}
   );
   gpc615_5 gpc652 (
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10]},
      {stage3_14[0]},
      {stage3_15[4], stage3_15[5], stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9]},
      {stage4_17[1],stage4_16[1],stage4_15[1],stage4_14[3],stage4_13[4]}
   );
   gpc615_5 gpc653 (
      {stage3_13[11], stage3_13[12], stage3_13[13], stage3_13[14], stage3_13[15]},
      {stage3_14[1]},
      {stage3_15[10], stage3_15[11], stage3_15[12], stage3_15[13], stage3_15[14], stage3_15[15]},
      {stage4_17[2],stage4_16[2],stage4_15[2],stage4_14[4],stage4_13[5]}
   );
   gpc606_5 gpc654 (
      {stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5], stage3_14[6], stage3_14[7]},
      {stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5], stage3_16[6]},
      {stage4_18[0],stage4_17[3],stage4_16[3],stage4_15[3],stage4_14[5]}
   );
   gpc615_5 gpc655 (
      {stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage3_17[0]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[0],stage4_18[1],stage4_17[4],stage4_16[4]}
   );
   gpc623_5 gpc656 (
      {stage3_16[12], stage3_16[13], stage3_16[14]},
      {stage3_17[1], stage3_17[2]},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], 1'b0},
      {stage4_20[1],stage4_19[1],stage4_18[2],stage4_17[5],stage4_16[5]}
   );
   gpc615_5 gpc657 (
      {stage3_17[3], stage3_17[4], stage3_17[5], stage3_17[6], stage3_17[7]},
      {1'b0},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[2],stage4_19[2],stage4_18[3],stage4_17[6]}
   );
   gpc1_1 gpc658 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc659 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc660 (
      {stage3_0[2]},
      {stage4_0[2]}
   );
   gpc1_1 gpc661 (
      {stage3_0[3]},
      {stage4_0[3]}
   );
   gpc1_1 gpc662 (
      {stage3_0[4]},
      {stage4_0[4]}
   );
   gpc1_1 gpc663 (
      {stage3_0[5]},
      {stage4_0[5]}
   );
   gpc1_1 gpc664 (
      {stage3_0[6]},
      {stage4_0[6]}
   );
   gpc1_1 gpc665 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc666 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc667 (
      {stage3_1[2]},
      {stage4_1[2]}
   );
   gpc1_1 gpc668 (
      {stage3_1[3]},
      {stage4_1[3]}
   );
   gpc1_1 gpc669 (
      {stage3_1[4]},
      {stage4_1[4]}
   );
   gpc1_1 gpc670 (
      {stage3_2[10]},
      {stage4_2[2]}
   );
   gpc1_1 gpc671 (
      {stage3_2[11]},
      {stage4_2[3]}
   );
   gpc1_1 gpc672 (
      {stage3_2[12]},
      {stage4_2[4]}
   );
   gpc1_1 gpc673 (
      {stage3_2[13]},
      {stage4_2[5]}
   );
   gpc1_1 gpc674 (
      {stage3_2[14]},
      {stage4_2[6]}
   );
   gpc1_1 gpc675 (
      {stage3_2[15]},
      {stage4_2[7]}
   );
   gpc1_1 gpc676 (
      {stage3_2[16]},
      {stage4_2[8]}
   );
   gpc1_1 gpc677 (
      {stage3_2[17]},
      {stage4_2[9]}
   );
   gpc1_1 gpc678 (
      {stage3_2[18]},
      {stage4_2[10]}
   );
   gpc1_1 gpc679 (
      {stage3_3[12]},
      {stage4_3[4]}
   );
   gpc1_1 gpc680 (
      {stage3_3[13]},
      {stage4_3[5]}
   );
   gpc1_1 gpc681 (
      {stage3_4[14]},
      {stage4_4[4]}
   );
   gpc1_1 gpc682 (
      {stage3_6[10]},
      {stage4_6[6]}
   );
   gpc1_1 gpc683 (
      {stage3_7[12]},
      {stage4_7[6]}
   );
   gpc1_1 gpc684 (
      {stage3_7[13]},
      {stage4_7[7]}
   );
   gpc1_1 gpc685 (
      {stage3_8[14]},
      {stage4_8[4]}
   );
   gpc1_1 gpc686 (
      {stage3_8[15]},
      {stage4_8[5]}
   );
   gpc1_1 gpc687 (
      {stage3_8[16]},
      {stage4_8[6]}
   );
   gpc1_1 gpc688 (
      {stage3_9[18]},
      {stage4_9[5]}
   );
   gpc1_1 gpc689 (
      {stage3_9[19]},
      {stage4_9[6]}
   );
   gpc1_1 gpc690 (
      {stage3_10[12]},
      {stage4_10[7]}
   );
   gpc1_1 gpc691 (
      {stage3_10[13]},
      {stage4_10[8]}
   );
   gpc1_1 gpc692 (
      {stage3_10[14]},
      {stage4_10[9]}
   );
   gpc1_1 gpc693 (
      {stage3_11[6]},
      {stage4_11[5]}
   );
   gpc1_1 gpc694 (
      {stage3_11[7]},
      {stage4_11[6]}
   );
   gpc1_1 gpc695 (
      {stage3_11[8]},
      {stage4_11[7]}
   );
   gpc1_1 gpc696 (
      {stage3_11[9]},
      {stage4_11[8]}
   );
   gpc1_1 gpc697 (
      {stage3_11[10]},
      {stage4_11[9]}
   );
   gpc1_1 gpc698 (
      {stage3_11[11]},
      {stage4_11[10]}
   );
   gpc1_1 gpc699 (
      {stage3_11[12]},
      {stage4_11[11]}
   );
   gpc1_1 gpc700 (
      {stage3_12[12]},
      {stage4_12[3]}
   );
   gpc1_1 gpc701 (
      {stage3_12[13]},
      {stage4_12[4]}
   );
   gpc1_1 gpc702 (
      {stage3_12[14]},
      {stage4_12[5]}
   );
   gpc1_1 gpc703 (
      {stage3_12[15]},
      {stage4_12[6]}
   );
   gpc1_1 gpc704 (
      {stage3_14[8]},
      {stage4_14[6]}
   );
   gpc1_1 gpc705 (
      {stage3_14[9]},
      {stage4_14[7]}
   );
   gpc1_1 gpc706 (
      {stage3_15[16]},
      {stage4_15[4]}
   );
   gpc1_1 gpc707 (
      {stage3_15[17]},
      {stage4_15[5]}
   );
   gpc1_1 gpc708 (
      {stage3_17[8]},
      {stage4_17[7]}
   );
   gpc1_1 gpc709 (
      {stage3_17[9]},
      {stage4_17[8]}
   );
   gpc1_1 gpc710 (
      {stage3_17[10]},
      {stage4_17[9]}
   );
   gpc1_1 gpc711 (
      {stage3_19[6]},
      {stage4_19[3]}
   );
   gpc1_1 gpc712 (
      {stage3_19[7]},
      {stage4_19[4]}
   );
   gpc1_1 gpc713 (
      {stage3_20[0]},
      {stage4_20[3]}
   );
   gpc606_5 gpc714 (
      {stage4_0[0], stage4_0[1], stage4_0[2], stage4_0[3], stage4_0[4], stage4_0[5]},
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], stage4_2[4], stage4_2[5]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0],stage5_0[0]}
   );
   gpc615_5 gpc715 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4]},
      {stage4_2[6]},
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5]},
      {stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1],stage5_1[1]}
   );
   gpc1343_5 gpc716 (
      {stage4_6[0], stage4_6[1], stage4_6[2]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3]},
      {stage4_8[0], stage4_8[1], stage4_8[2]},
      {stage4_9[0]},
      {stage5_10[0],stage5_9[0],stage5_8[0],stage5_7[0],stage5_6[0]}
   );
   gpc1343_5 gpc717 (
      {stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage4_7[4], stage4_7[5], stage4_7[6], stage4_7[7]},
      {stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage4_9[1]},
      {stage5_10[1],stage5_9[1],stage5_8[1],stage5_7[1],stage5_6[1]}
   );
   gpc1343_5 gpc718 (
      {stage4_9[2], stage4_9[3], stage4_9[4]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3]},
      {stage4_11[0], stage4_11[1], stage4_11[2]},
      {stage4_12[0]},
      {stage5_13[0],stage5_12[0],stage5_11[0],stage5_10[2],stage5_9[2]}
   );
   gpc7_3 gpc719 (
      {stage4_10[4], stage4_10[5], stage4_10[6], stage4_10[7], stage4_10[8], stage4_10[9], 1'b0},
      {stage5_12[1],stage5_11[1],stage5_10[3]}
   );
   gpc1343_5 gpc720 (
      {stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage4_12[1], stage4_12[2], stage4_12[3], stage4_12[4]},
      {stage4_13[0], stage4_13[1], stage4_13[2]},
      {stage4_14[0]},
      {stage5_15[0],stage5_14[0],stage5_13[1],stage5_12[2],stage5_11[2]}
   );
   gpc207_4 gpc721 (
      {stage4_11[6], stage4_11[7], stage4_11[8], stage4_11[9], stage4_11[10], stage4_11[11], 1'b0},
      {stage4_13[3], stage4_13[4]},
      {stage5_14[1],stage5_13[2],stage5_12[3],stage5_11[3]}
   );
   gpc615_5 gpc722 (
      {stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage4_15[0]},
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5]},
      {stage5_18[0],stage5_17[0],stage5_16[0],stage5_15[1],stage5_14[2]}
   );
   gpc615_5 gpc723 (
      {stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4], stage4_15[5]},
      {1'b0},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[1],stage5_17[1],stage5_16[1],stage5_15[2]}
   );
   gpc1_1 gpc724 (
      {stage4_0[6]},
      {stage5_0[1]}
   );
   gpc1_1 gpc725 (
      {stage4_2[7]},
      {stage5_2[2]}
   );
   gpc1_1 gpc726 (
      {stage4_2[8]},
      {stage5_2[3]}
   );
   gpc1_1 gpc727 (
      {stage4_2[9]},
      {stage5_2[4]}
   );
   gpc1_1 gpc728 (
      {stage4_2[10]},
      {stage5_2[5]}
   );
   gpc1_1 gpc729 (
      {stage4_4[0]},
      {stage5_4[2]}
   );
   gpc1_1 gpc730 (
      {stage4_4[1]},
      {stage5_4[3]}
   );
   gpc1_1 gpc731 (
      {stage4_4[2]},
      {stage5_4[4]}
   );
   gpc1_1 gpc732 (
      {stage4_4[3]},
      {stage5_4[5]}
   );
   gpc1_1 gpc733 (
      {stage4_4[4]},
      {stage5_4[6]}
   );
   gpc1_1 gpc734 (
      {stage4_5[0]},
      {stage5_5[1]}
   );
   gpc1_1 gpc735 (
      {stage4_5[1]},
      {stage5_5[2]}
   );
   gpc1_1 gpc736 (
      {stage4_5[2]},
      {stage5_5[3]}
   );
   gpc1_1 gpc737 (
      {stage4_5[3]},
      {stage5_5[4]}
   );
   gpc1_1 gpc738 (
      {stage4_6[6]},
      {stage5_6[2]}
   );
   gpc1_1 gpc739 (
      {stage4_8[6]},
      {stage5_8[2]}
   );
   gpc1_1 gpc740 (
      {stage4_9[5]},
      {stage5_9[3]}
   );
   gpc1_1 gpc741 (
      {stage4_9[6]},
      {stage5_9[4]}
   );
   gpc1_1 gpc742 (
      {stage4_12[5]},
      {stage5_12[4]}
   );
   gpc1_1 gpc743 (
      {stage4_12[6]},
      {stage5_12[5]}
   );
   gpc1_1 gpc744 (
      {stage4_13[5]},
      {stage5_13[3]}
   );
   gpc1_1 gpc745 (
      {stage4_14[6]},
      {stage5_14[3]}
   );
   gpc1_1 gpc746 (
      {stage4_14[7]},
      {stage5_14[4]}
   );
   gpc1_1 gpc747 (
      {stage4_17[6]},
      {stage5_17[2]}
   );
   gpc1_1 gpc748 (
      {stage4_17[7]},
      {stage5_17[3]}
   );
   gpc1_1 gpc749 (
      {stage4_17[8]},
      {stage5_17[4]}
   );
   gpc1_1 gpc750 (
      {stage4_17[9]},
      {stage5_17[5]}
   );
   gpc1_1 gpc751 (
      {stage4_18[0]},
      {stage5_18[2]}
   );
   gpc1_1 gpc752 (
      {stage4_18[1]},
      {stage5_18[3]}
   );
   gpc1_1 gpc753 (
      {stage4_18[2]},
      {stage5_18[4]}
   );
   gpc1_1 gpc754 (
      {stage4_18[3]},
      {stage5_18[5]}
   );
   gpc1_1 gpc755 (
      {stage4_19[0]},
      {stage5_19[1]}
   );
   gpc1_1 gpc756 (
      {stage4_19[1]},
      {stage5_19[2]}
   );
   gpc1_1 gpc757 (
      {stage4_19[2]},
      {stage5_19[3]}
   );
   gpc1_1 gpc758 (
      {stage4_19[3]},
      {stage5_19[4]}
   );
   gpc1_1 gpc759 (
      {stage4_19[4]},
      {stage5_19[5]}
   );
   gpc1_1 gpc760 (
      {stage4_20[0]},
      {stage5_20[0]}
   );
   gpc1_1 gpc761 (
      {stage4_20[1]},
      {stage5_20[1]}
   );
   gpc1_1 gpc762 (
      {stage4_20[2]},
      {stage5_20[2]}
   );
   gpc1_1 gpc763 (
      {stage4_20[3]},
      {stage5_20[3]}
   );
   gpc1_1 gpc764 (
      {stage4_21[0]},
      {stage5_21[0]}
   );
   gpc615_5 gpc765 (
      {stage5_2[0], stage5_2[1], stage5_2[2], stage5_2[3], stage5_2[4]},
      {stage5_3[0]},
      {stage5_4[0], stage5_4[1], stage5_4[2], stage5_4[3], stage5_4[4], stage5_4[5]},
      {stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0],stage6_2[0]}
   );
   gpc135_4 gpc766 (
      {stage5_5[0], stage5_5[1], stage5_5[2], stage5_5[3], stage5_5[4]},
      {stage5_6[0], stage5_6[1], stage5_6[2]},
      {stage5_7[0]},
      {stage6_8[0],stage6_7[0],stage6_6[1],stage6_5[1]}
   );
   gpc1343_5 gpc767 (
      {stage5_8[0], stage5_8[1], stage5_8[2]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3]},
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[0],stage6_10[0],stage6_9[0],stage6_8[1]}
   );
   gpc1163_5 gpc768 (
      {stage5_11[1], stage5_11[2], stage5_11[3]},
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5]},
      {stage5_13[0]},
      {stage5_14[0]},
      {stage6_15[0],stage6_14[0],stage6_13[0],stage6_12[1],stage6_11[1]}
   );
   gpc1343_5 gpc769 (
      {stage5_13[1], stage5_13[2], stage5_13[3]},
      {stage5_14[1], stage5_14[2], stage5_14[3], stage5_14[4]},
      {stage5_15[0], stage5_15[1], stage5_15[2]},
      {stage5_16[0]},
      {stage6_17[0],stage6_16[0],stage6_15[1],stage6_14[1],stage6_13[1]}
   );
   gpc606_5 gpc770 (
      {stage5_17[0], stage5_17[1], stage5_17[2], stage5_17[3], stage5_17[4], stage5_17[5]},
      {stage5_19[0], stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage6_21[0],stage6_20[0],stage6_19[0],stage6_18[0],stage6_17[1]}
   );
   gpc1406_5 gpc771 (
      {stage5_18[0], stage5_18[1], stage5_18[2], stage5_18[3], stage5_18[4], stage5_18[5]},
      {stage5_20[0], stage5_20[1], stage5_20[2], stage5_20[3]},
      {stage5_21[0]},
      {stage6_22[0],stage6_21[1],stage6_20[1],stage6_19[1],stage6_18[1]}
   );
   gpc1_1 gpc772 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc773 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc774 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc775 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc776 (
      {stage5_2[5]},
      {stage6_2[1]}
   );
   gpc1_1 gpc777 (
      {stage5_3[1]},
      {stage6_3[1]}
   );
   gpc1_1 gpc778 (
      {stage5_4[6]},
      {stage6_4[1]}
   );
   gpc1_1 gpc779 (
      {stage5_7[1]},
      {stage6_7[1]}
   );
   gpc1_1 gpc780 (
      {stage5_9[4]},
      {stage6_9[1]}
   );
   gpc1_1 gpc781 (
      {stage5_10[3]},
      {stage6_10[1]}
   );
   gpc1_1 gpc782 (
      {stage5_16[1]},
      {stage6_16[1]}
   );
endmodule

module testbench();
    reg [161:0] src0;
    reg [161:0] src1;
    reg [161:0] src2;
    reg [161:0] src3;
    reg [161:0] src4;
    reg [161:0] src5;
    reg [161:0] src6;
    reg [161:0] src7;
    reg [161:0] src8;
    reg [161:0] src9;
    reg [161:0] src10;
    reg [161:0] src11;
    reg [161:0] src12;
    reg [161:0] src13;
    reg [161:0] src14;
    reg [161:0] src15;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [23:0] srcsum;
    wire [23:0] dstsum;
    wire test;
    compressor_CLA162_16 compressor_CLA162_16(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127] + src0[128] + src0[129] + src0[130] + src0[131] + src0[132] + src0[133] + src0[134] + src0[135] + src0[136] + src0[137] + src0[138] + src0[139] + src0[140] + src0[141] + src0[142] + src0[143] + src0[144] + src0[145] + src0[146] + src0[147] + src0[148] + src0[149] + src0[150] + src0[151] + src0[152] + src0[153] + src0[154] + src0[155] + src0[156] + src0[157] + src0[158] + src0[159] + src0[160] + src0[161])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127] + src1[128] + src1[129] + src1[130] + src1[131] + src1[132] + src1[133] + src1[134] + src1[135] + src1[136] + src1[137] + src1[138] + src1[139] + src1[140] + src1[141] + src1[142] + src1[143] + src1[144] + src1[145] + src1[146] + src1[147] + src1[148] + src1[149] + src1[150] + src1[151] + src1[152] + src1[153] + src1[154] + src1[155] + src1[156] + src1[157] + src1[158] + src1[159] + src1[160] + src1[161])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127] + src2[128] + src2[129] + src2[130] + src2[131] + src2[132] + src2[133] + src2[134] + src2[135] + src2[136] + src2[137] + src2[138] + src2[139] + src2[140] + src2[141] + src2[142] + src2[143] + src2[144] + src2[145] + src2[146] + src2[147] + src2[148] + src2[149] + src2[150] + src2[151] + src2[152] + src2[153] + src2[154] + src2[155] + src2[156] + src2[157] + src2[158] + src2[159] + src2[160] + src2[161])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127] + src3[128] + src3[129] + src3[130] + src3[131] + src3[132] + src3[133] + src3[134] + src3[135] + src3[136] + src3[137] + src3[138] + src3[139] + src3[140] + src3[141] + src3[142] + src3[143] + src3[144] + src3[145] + src3[146] + src3[147] + src3[148] + src3[149] + src3[150] + src3[151] + src3[152] + src3[153] + src3[154] + src3[155] + src3[156] + src3[157] + src3[158] + src3[159] + src3[160] + src3[161])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127] + src4[128] + src4[129] + src4[130] + src4[131] + src4[132] + src4[133] + src4[134] + src4[135] + src4[136] + src4[137] + src4[138] + src4[139] + src4[140] + src4[141] + src4[142] + src4[143] + src4[144] + src4[145] + src4[146] + src4[147] + src4[148] + src4[149] + src4[150] + src4[151] + src4[152] + src4[153] + src4[154] + src4[155] + src4[156] + src4[157] + src4[158] + src4[159] + src4[160] + src4[161])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127] + src5[128] + src5[129] + src5[130] + src5[131] + src5[132] + src5[133] + src5[134] + src5[135] + src5[136] + src5[137] + src5[138] + src5[139] + src5[140] + src5[141] + src5[142] + src5[143] + src5[144] + src5[145] + src5[146] + src5[147] + src5[148] + src5[149] + src5[150] + src5[151] + src5[152] + src5[153] + src5[154] + src5[155] + src5[156] + src5[157] + src5[158] + src5[159] + src5[160] + src5[161])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127] + src6[128] + src6[129] + src6[130] + src6[131] + src6[132] + src6[133] + src6[134] + src6[135] + src6[136] + src6[137] + src6[138] + src6[139] + src6[140] + src6[141] + src6[142] + src6[143] + src6[144] + src6[145] + src6[146] + src6[147] + src6[148] + src6[149] + src6[150] + src6[151] + src6[152] + src6[153] + src6[154] + src6[155] + src6[156] + src6[157] + src6[158] + src6[159] + src6[160] + src6[161])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127] + src7[128] + src7[129] + src7[130] + src7[131] + src7[132] + src7[133] + src7[134] + src7[135] + src7[136] + src7[137] + src7[138] + src7[139] + src7[140] + src7[141] + src7[142] + src7[143] + src7[144] + src7[145] + src7[146] + src7[147] + src7[148] + src7[149] + src7[150] + src7[151] + src7[152] + src7[153] + src7[154] + src7[155] + src7[156] + src7[157] + src7[158] + src7[159] + src7[160] + src7[161])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127] + src8[128] + src8[129] + src8[130] + src8[131] + src8[132] + src8[133] + src8[134] + src8[135] + src8[136] + src8[137] + src8[138] + src8[139] + src8[140] + src8[141] + src8[142] + src8[143] + src8[144] + src8[145] + src8[146] + src8[147] + src8[148] + src8[149] + src8[150] + src8[151] + src8[152] + src8[153] + src8[154] + src8[155] + src8[156] + src8[157] + src8[158] + src8[159] + src8[160] + src8[161])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127] + src9[128] + src9[129] + src9[130] + src9[131] + src9[132] + src9[133] + src9[134] + src9[135] + src9[136] + src9[137] + src9[138] + src9[139] + src9[140] + src9[141] + src9[142] + src9[143] + src9[144] + src9[145] + src9[146] + src9[147] + src9[148] + src9[149] + src9[150] + src9[151] + src9[152] + src9[153] + src9[154] + src9[155] + src9[156] + src9[157] + src9[158] + src9[159] + src9[160] + src9[161])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127] + src10[128] + src10[129] + src10[130] + src10[131] + src10[132] + src10[133] + src10[134] + src10[135] + src10[136] + src10[137] + src10[138] + src10[139] + src10[140] + src10[141] + src10[142] + src10[143] + src10[144] + src10[145] + src10[146] + src10[147] + src10[148] + src10[149] + src10[150] + src10[151] + src10[152] + src10[153] + src10[154] + src10[155] + src10[156] + src10[157] + src10[158] + src10[159] + src10[160] + src10[161])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127] + src11[128] + src11[129] + src11[130] + src11[131] + src11[132] + src11[133] + src11[134] + src11[135] + src11[136] + src11[137] + src11[138] + src11[139] + src11[140] + src11[141] + src11[142] + src11[143] + src11[144] + src11[145] + src11[146] + src11[147] + src11[148] + src11[149] + src11[150] + src11[151] + src11[152] + src11[153] + src11[154] + src11[155] + src11[156] + src11[157] + src11[158] + src11[159] + src11[160] + src11[161])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127] + src12[128] + src12[129] + src12[130] + src12[131] + src12[132] + src12[133] + src12[134] + src12[135] + src12[136] + src12[137] + src12[138] + src12[139] + src12[140] + src12[141] + src12[142] + src12[143] + src12[144] + src12[145] + src12[146] + src12[147] + src12[148] + src12[149] + src12[150] + src12[151] + src12[152] + src12[153] + src12[154] + src12[155] + src12[156] + src12[157] + src12[158] + src12[159] + src12[160] + src12[161])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127] + src13[128] + src13[129] + src13[130] + src13[131] + src13[132] + src13[133] + src13[134] + src13[135] + src13[136] + src13[137] + src13[138] + src13[139] + src13[140] + src13[141] + src13[142] + src13[143] + src13[144] + src13[145] + src13[146] + src13[147] + src13[148] + src13[149] + src13[150] + src13[151] + src13[152] + src13[153] + src13[154] + src13[155] + src13[156] + src13[157] + src13[158] + src13[159] + src13[160] + src13[161])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127] + src14[128] + src14[129] + src14[130] + src14[131] + src14[132] + src14[133] + src14[134] + src14[135] + src14[136] + src14[137] + src14[138] + src14[139] + src14[140] + src14[141] + src14[142] + src14[143] + src14[144] + src14[145] + src14[146] + src14[147] + src14[148] + src14[149] + src14[150] + src14[151] + src14[152] + src14[153] + src14[154] + src14[155] + src14[156] + src14[157] + src14[158] + src14[159] + src14[160] + src14[161])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127] + src15[128] + src15[129] + src15[130] + src15[131] + src15[132] + src15[133] + src15[134] + src15[135] + src15[136] + src15[137] + src15[138] + src15[139] + src15[140] + src15[141] + src15[142] + src15[143] + src15[144] + src15[145] + src15[146] + src15[147] + src15[148] + src15[149] + src15[150] + src15[151] + src15[152] + src15[153] + src15[154] + src15[155] + src15[156] + src15[157] + src15[158] + src15[159] + src15[160] + src15[161])<<15);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h5935c9ca446c81922044bc4bc3dcf1e5eecdf403c30de3704bae1febfb28a1ce5ce50f2b77065d4fa4182b541573e2345d1419b7f5a2933ec583737f342a197b922abb2b2aa72cf42ef61872387516e43ce3203df5c8913892bf5c96288729914001b4f918fc9a970f9d564071890b1d7862bfc3c7834ca84a52625392660bdbb66e9595c50d8a9a10dfc933ec1f014104965554a0a57fc34937b38b734ce87afdd07c5a964bc304157305862d8c527d11878c448a3f3ddb1dceed3b7e26751f6bffcd035378f8993f74abacc1fba10d63feefad1ed5384d7303b09bf322d8d8af6f0609c66209734a70d8e18e9a1b125409c467f74aabb67035d893cc7cf3b34eb7afac815fb9f92dfac554bb1be5c3ffad5f039f37d809c7464e71b0b0831cb5d261af5583a15c4dacdadb4d2d371b00089bd0041be7caccba657d3840a76091b8e3f8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h97601c9971c4bbaef2b1d0b8cdf6f06625a1a506a05c8044c21483c239da51827699facb239279dff1056b68dbeb3627eef7f332a7b3fe104a0704f6c9ed02517c6a01698f71dc56f5aab0a588e507c2ece4d391e2a3c675469ed0c89d6a916c3f3b04901e8fa6c03382b04186ca5071be5d7972f3c1b5c48d464ff221cfa30252dbf3bd3fae863af1d5e7e607fce15af2d224063f95810251537a2a8b11c6d1baaebe39d2e2c5e55cf3fa5b35e84cba428d9e276ed1cf06f933c82d7162b490109f192f74cff142d20b86d1e5c827dbfa8287d18692f85151c8780cf4dd34601079df2351d17f80f2b80d9a30f0a2ce9c8f26f1efe709a9eb6f9f412d7dcde204adbbe97d1f3b28535119e1c92917af92f83515c111e2ad938384a9ad6471ed08408148ef541cf0f4d60a3197df5e15035f2b7271e0a4e14dfd522ec50e333f88ee2398;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h3047620ae7ff855e0f4a76fc8660c5d47244812b99ade35c36244126ca3f65200ffe533013d5a284d4c3c7155ab6efb272c70ca362148b47c61749ab740de5380b4b78aba622ded025cedd12cefa379ccd906a77c130c7babd4f9d584bae788afe038755e1245ffd5290d27c65b8c9154fcde539b4c06727046c226feed402bdc3963e9c1bd2a8efaf2ccba392c84aaf1bda733740bd0eb020274874b927d577d253d33abd592a86945f8662c2c87d3ae2524b8070b73457df5262d0de77f39b6a53d738f74ee299d79a868e96175fa88e5c614a5aa93be98f56b82e1b7560af4c7fd695c76e4c16f91adfbd7f746965827001d19c2c86d593bb458ccadd6929d8c35ea499e4a684b508c1a52a8c0c2b7a1be748bc6625aa51d143138acb2522f920d4090aef7535d2bea811deeed00db49344b27d637d15bbfcf7e3981300b805953069;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h5208103a8ba4a2a8819bccac45a16787ea2973914ef39bbe8d070e2e280f301c67d43db5f197fffe2e7813047a18da90237f4b9ff8f0cffe9fa69f563472ddd5a1d38a5641753d57052785cbb0d15f31dbf0e045e0693ebf773437716816b0bcbaa7de273bcb3ca65962d7e2ebb3e9e48f72a316e42172cd9ccaf6e2b4a9fcb9d923dea2f23b52f0c763774ddb89b26e22433ac27bdfcc02a7cb0d40780f60e583d1c4afbd8fb7a83f106830eb601e7858b993a8076a84633c1707ce6884b6e0c23492038ec902b911614cd853a82601f580837f6c6cac4f07689e526dd2ce633ed4a9e81a8328f70cadf7f1a8df324c6300f8836af52af822a73944400c1327575204b9eee934ef148e400d509141ed7a2215e4ddf963543cf6d93b3ab7e352dd16dc37fb94c6cda7fe448f79eb47094e71d7b6a3366b00a0dab0136692afb1356edd15;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hc11419a3350e2b58d21486f9bf22d5ef48191d8559dfbcfae5940aacb4b1ee96c25db01292e233e7495fd353d6ca479a9fb0bee19b915f9aaa25b3e2a298030db6880020554ce68a2de2dfe4351950de22aa4932de7f632821868b2bc522409df3564202fd9c63076373eea7e4b27056ed56a049a2f22fc9e23cc16b2c6bf1a703bb07d4b080157007ff370716caa8a5730f21745d3c59a66629161836caa467ff544dd0533f01899177faac5437cb253de00dfe69782007db46453fa72b820efe151d83cd553c23f61e57aa098c8c39d06033a392e83b984396d9c18bc330172429acfd796a63e350c10d893d01007f403827a142423af75362bed36ea011b1e5975273bae3c8edc8d9b6cf520f903951f2bbadf787febbe6dacfbd319942215b8e95c9a41c312e6f017b6e17664840137b09174a224e31a558c04f764c2dbfdd096dc2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'he2435f6d39a3cdc859a12d18ba53d755a3d345d0101ef2a802b201401f9208746c2a126621faf4105828d3fb11532654bae150eb616ca6074b854ccd217f9af1c657ff1125316f9ad803756d822217edc24175d305ccd2e0e39e78eb48756866fea8e34194924ac79241f44e945a2ffa8ccf9f454301b3f896180dbe9568953eb405684f6a8278ded0edbab9f48fd64432e55dd7e8b02efd078a98fbc7fa9f11c5afdd13bdf37b5f1b35d215dc83b47354ed2ed0a3c3fa62ee8a7ab9c7d52e3f9dcc8d6bd6a2c094b19300dcaa671a2b06e9e028c78cb54ed840c45c51a211810a2ec0370b2c01d7033df079222976d25556a9979b1688d17183e3a389013c2e1178920e7515a25e3276d8af71864d24891f1b3e096430941369abf30d79ba3c2c0c92d2051a0e8ff659269d6513270042e25751f05b53a567a7cd03794668125c95ae2b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h4c39038833fda9c9ae1190cc5baff5a2ef74814a651cf3b0e459ade622895531d4b7e3cfd595cd2e620e6a51bc7fb7919b4660490dd076ea6fa4bce48152c1bb9cf3f5e1067dff32e60b5524ade739cb5aaa36fb36b7896410b864ceca8d7bd8da8c29b4d64e86b0f1d8a2bc2fa9837b53a0bfba57fc5cd7731abe2f2b4f3c2cd93e00a075554e796977d06b900d894a2fe36eab353a2d9c3c225db460124a2427c3f01adb7849295db30f9207c30e89e5ce21ea050feaa40dd3458a53d997273218886efafbe0921239c94444f84c0968c1fec6b28d5792ee3f3993baff913c12db5dc3f1adaf71404781d463fdc003b932f61e6b8b03d1c35c6629dcf63c2ad394419780d77d51d016b355eb9d13a7e53dc24cd5ded4763eeca3adb6594f228aecdadb9b4fca4158bf58c176b6ed92f22ad13936f9773ce5e3e0dc27d8d8c765974e02;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h174220df82fa2a069495cce0baed57debcb2e495cdcb1811278f9daa2cb75eb1f0bd58cdbbf8f7c50dfa743f004b0ee82a37932067d0ac5e51fa455e4a9c5a5f6b2ec8341d3b1ea5e21a6b55add8a3cd100d009131bac0d684f4e4f10c1e57082325042174592cc96c681ddee18e331d6a76561d6c1fc8d62a35b4b55a02a94bda694245663259d0ef95e11677dccf7da8d0e7cf45c5e48d666c9bb80f2e945a286fc1093f3aa85c8cf7200ea850821546540c434a1ab9cc4a8ec3972be16cdcfec07880ad83a5d2108ccec432bd68b50502b556cf3761ef46f0df88c6d5d487f24a054f840a4a847d7c3e330747e9afbf3ea2ef5b88352a1128f8af5cc4a8996f78930af782547ef1433256619cada9353d5310def23f00eda2299c2d74f106f5eeaeb2d5c617b68d201229adb6ce5cb68ad02552dcc6ae1863e69c3f7b5078960849b2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h1628547755c2185946a652814e5bcb8881425fe062be2583af6e2bbf4f4e6032f029fc2177b72f4974ea03bd69cc7e279f78400c07a54c990a138262ea3bd3405b20c24bffaf15a492631785e920ca320bf17aa52100d9952a796de679eb690ce3a450f391b0889029140cbdb4e15527d64e36c1238a7d8c871cb2a8a0f026ea0db3e539cb4228ba68c4c311ef5c62fa71b990588e4494dbd8880e777bcdfceab6df8d4540b4af9b88df868b253db89f991b7b2f690a6a35888a714ceaf9e670420b0c1de127d0a7c169dbaeef5c1a4d3f7c036a840b4455b67f80d9be5b8b1c06cf70bc306bf95b25fa745fd0c9d388c2b9f9895afa4dd2efc3d44564741bc51ef5c9fd7d80e2e0d449fdcc2555670b9f7a26bbbc496c892d112f1eefc7865e15e74cad3a645924f29c773314b3f82a8a163932890111da99bc4865a3a9dc38f48927e2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hb279786f92f4317511c72c3d4a8c908b9f7760040725c1b5f309bdbf4f51a353694e8157c8cf8b83233ef0375b6ed39a05cfcac224643d3dd3706f58e022d2b274899e26b12fba0c0c138ea7fe214fd8357afaaa26f5a12cf2d20a6e74b85f3c01a4e60cac070b0d745f0ad382cf6a584e3db9d45f905efa7035956c38e54c312f308c3683f63dd08f7ffc992117217531db1b153a1664e10d42e68aac91c86171233f535020d39e9c197ccaced6f04b567eefd2e253ae4ff3abb2dd14917905556fc5f29b27e46988b1a85b3f23ca052f283f481172de7ce0a6a3fb8923b4f3919e63e0bfe57866a5496ee25200186d28f57667c84b2426c9359583531355da9d0fdf5bdb95845d9ff7cde73ecdeb7391e223b871e2f927fbca1d35182a8bbe4f9faeb2415e2adfbb49aa4a7f035503e33e80672348173061ff13b6babf0a55e4dcfeb2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h68ddbd3fbe5141e926312d26bbd20b159b8513f962709b52c05f4a49e5bf1e1b0690011dbaaadf1493301a7380b109542b18a05c5ef5b9eac1739abc7f69722a124fd7dba773f9f1f7936a466694ba15cc5fba7feea65a67cf576c405a523d17b1ae5efd392d9b7458bf7caf06305c1f62acc88b25e12e9d78ee47ab401ac03428f7bc5624245d6442ec0ec9f7998d1a62c54cd9d8e62b6f779a97211e943fa1cf07076cb5641dfc96f0b8fe7b0e16b550b27d77b12c12ee262f4f76b3465e09a21d266ea5ec50015bee62feffb9ce1eeaa26f8fc0c3058153bf59500bc64d736d808f963cd26d06e5b095cb0c91cc7baaca4226f2e426dee20dea855c67c0c33cee05b00fb778f20912b7e7594d94a0fc1cb171f8a55dd8860af11450e680d914e72df8f9c04ef940b6636a838227f7af88424338baeeb45b161e932688e1b76cbd4344;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h1b783add0264a3e80eb5ce3fc37edaf72f0e28a15a53f2f80c2c0baa19889f5a7908dee160c7ac0f7b9487d30114a8dbe3e98b401a98dd7c415d12509b2a8abfb7a694b385dfff9f407004bf72b57636629471c044b7346de46ad6406214a65c69a27a008e947f57855a2c923606b64f5b9b55babdc52af461ad0c0856c7f3def4347afca297ac48ba5afeed532401d9565140ab576de025693d4ed12e6d696a8f1a80ceb718e9b1a661dcb4a4ab922170fe10e5792d19d9b0a74a78c71dfdb6714282e774c46f59d64c85cb4257b3ba826c545a10ea3c6f6f4c62a879cf8c815b48819d188b54df17ba34c3e510a89a20507dd290e01fd6005633c0f5bd42905d01bd19d07bf7ba22e714dbaaed0f97e45a05e681a2c55e9ad48c8da5168de5c58970d922992dc80c2e6091c755806865308bbc735db9a0f94aac8a4071a811e6dafa70;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'had0ba5239ea42c6f6a9920c5b2ae6ed172b1bc66a96b1c25743e0a88cee900ec2fbe7c4fe7ed7399652c2297871126dd04599b38e7bb1be3474fd20c8342062359f4f11e9e9a334e21ea7200174b00124b55e03fbbac2ec9ff49ac22c2a29df0dc673abe54bbf148c350b777568b099a09fbac27adfbeb8e93d250e296c93f4343858e3d97993c47aec9d3e17b5367971aa61dce6ddb93cfc45612d1c7b007622083a6eda5fe970b27205de267f9699b1f212fbc5efbf318be4f7c23ddcd774246fc9411b1d39e2e279f31b77a7b554c5c07628e2c0d9c1cdffd44549a0cc9f899c3a88ee6583d25f7350a8e31598dfd90639980bf3730b770db91069b4961a9a4456703c8d3b7c6d8a9e14ca4cda889833e00312cc7290e460923bb45eb0be779f72624c418eba2ac7cbf9356900a9ae69c116b6949a31fb17020772ed95cbe1abcdeb4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h17e61fd79e16f9f3d837ee5ee2dbe7fbd8e4d5d376f07e732dc56cedcac1c3e297187f5902b85a0b611d06b8a2cbcb4c1f4738765aa7fa18c2ff230af55b5929c43cd4171ceb4a81789a82f7c798232ecb4b1c352bb6b1a360bfd585db68889dcb553b586f1d13fec768ffd874f5626501774d597239e38450476d1377ccbe2ed3c6fed785f3ca646b31136af30c774a08339abf1116fbf3a5506ac80730877b5934796f51a3b118d1d88d009f21028c8adf4f98bfdc1065cd74a6d819e4949b5c1206368b57c169009502a48d8e0d987b3cd1f4d52261c526c873bcc590065941eed4b4c4d6b5edcdfe77abf5afa4e5be5c3e68d4f4d17f3e2b5416d8f2b5e18f9c81aaadc2f6f9fb37e2cd850a8c73246c1b06259f4f32222823b8e6c7ed7c78dc9b401b2a6e1578dac42df44756a0f05916d1b5bd5a86fb77d6f75c0f11aa03175eb8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h7290df1571dbd8a2a93d5ea02c51e8418d820c29d8672e6d2bba8c35242593358744b8c4fcfabe24d2c93244ff8c828d70972dcd78f4ec8d41c80cc3f989ecd636b669ac8b89238683e1e5ab8a05f2b4c85dd8e3c50e1d882225177dbb5ad047f68d6882727dcf7aa3845bd025372fa1987b99212bcd06787c46356526bb1d78f8a147cd7effbef8bff742bc818622e6d6492eda6a466eaa23507750be802311be74b9dfaa98e7486471518224b1c29bce55c08d1cbe8f3210978770bd3a017116c45692ab20950f8e11a6a3190ad8658086c98f7039081b555e4508b1aafd66f451c2e6c0f23967f492d3b385e534bb307ac0ec5c722d81ffbb2642f84c548d1bd0c42db2822bd5e81ec97254dc48646b8f1f72caad4dcda58180b5e6f0788f81301eca3a0e06f1fb9ab35c60c432276f5cd318e593839210c7b97038b88b719a1ff158;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hd1cd21ba0dc72dc62f64ecc4cae3f3b58132b766787b9b96be8cc7cbabcdc383e6816e0ab1c6cf0f3e62154d902d2398d766dd6376d0af5d1d5f9eef377407f18905c89aa91fa3e3f64b71d905b1db94c3e8c59059d221e95c413eef260d0e7ca517c4183d935eb9b0b6fd21f05febd5f6b7b24316242d66f71b6c764d1f5b7ea9abe770688ee21e015549d2a5284e1b74e62d960ad5d7555797395263e0ef46bdc341eb186ba321cf798f4f2e6fd644f4c844c45fc86cadd7f753c8f288d1653c1b9b76d4ed915dd03e95ef89093fbccd48bc8e68785e4af4d7b41c5af8ad20cb8d533042117b2c0a1496cb4ab5df24b97ba74901884dba1e7534128bce2864d256c1f05a5afcab562e5c5f08d347fb87c98cc688f0e7e21275ad19f758a86bebbf16134ee57833feee82344578b34e7a71270142e0b3c8c2d29b3a4f1c5019ad54156f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h91ff390b55b0ba7987563d82e899904044d0860114eb4135e9f8575d4cec9dd04e1830a203bd7fcfdbc29d01ef3bd3766a46191670809181ef6fe6ce314a43e1f5ce61babbb4234496c39ec85f911d107ea16a5326067a459bca3da1e90e5516176a1a511d0e5dd8078719f75cc42c7597ee1e91babf30d2346059062b37392460da7b5089baa018fb0b85b922b954c0cca9ff75cb5de68ce70361867aa33ff19dc1b5ae8ee576b7307293d0236c3be3c26c0b571c7604cbe98e91572ed2bde33dc5cf615af4fbbb9117256a392fb78097da82057fbe71f28101d204e665462a7496e84ac1b873a6eaa40e52037528c99a32ac1e944c3899a64630df90a92f17347df27f426bee43fdfb611b4cd7d1a4742c3bdd018f95c62987a974340ac96859c8354cbd2867b8c140c80a402515701ad8ced6a87c798d86e21c95595d9cc61b7a87b6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h3c5ff6d33e3b076f7a1ee50c89954ad4b9aed4cbd1e758b6719e7040c3cfaeac7b17f16fe7f8b9c6f1cdec742bf9d281113d128f5c5c3cfe069a6e56a744788c80618afe91629e40d165a4cae88aa70ec7a9950884d99518335192134a5bc3327114f9242c42f6022e3905dc7088a701b0197f82ccefffbfa0dcd224f268a1402a0f5bf747de53753e2147e8ebfa5463f5cd0b9bb27c0b0a7119f23fdb6ff9061e369a72f870b87fc9a46db7b6ba605b10d142dad12ec1174bf9127f9e96c28095e47322bb35822a6150179b751b6b2b7fd57ec0ca3755d8d6cb333cd58d18ab7545c7f75bfaf9637edb6682e0fcb9758d256c7c25293646c91703c574be9380e09fcb4f3564b4784f1dbf88b18ef41d3c0f7f96daf3194ab34df50752ea0cfd28fb2890191f3938ed731ebcafe5750df3e4cdf5416267275467e020a0fd5df380e21b86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'he73b2a17dbab94ebb827d4f07901bb22c23b89195b3d14453be79021532e9868fbdd214dff9d22f17a5b0b381f7890014ae711b4551357bc8e94af4a16969b0115e83192495f210c4cfca80bb838c371477983b67be399f0eab173afd2c0debfd97cf785a8a3a906d855483382fc52738fc6b8204e1ff2ce18c63f6f495eb220518e660b7acb8e080f198b73a57a491b02b795ff314787de56beeb759b3e8b7e4cff0fe4b3836ac724aef92deb4501e102c3ee732a89f3d0d4f0c8fdc1f7799f16517c895a7a402af75cbbf60fb3432486f3f3f9ce1bf8c79f1d50ea33d42023e6e35d5550fa53b0b02660c81de0b442e2ac5a2b5cfba12c75f69722bba87609335f3cb97ac2315a9e7e27076154157c86745b831d96dac6ba1daf899de489c0b38926b6af94174438cab5bc0f2b9b5603baddad6b6b45923f09016b52ec9aa5080505fc;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h8d983117b1f55e15dada516345e5b66b18aef553273045de6db9970ff3f443c77a1570aed3a9012e561387bc64a7bcbffe78d6820e563a57b809989aeb0f7ad580867b69d55435a27ad46f7b55d4244f206de42dc393a0e33bf48af407cba9bc631ea82ea9e4dbde8a7155efb55f8ad0ff5ba342ed8b6c06d59c56cb30429de9ab92f890f4581f7302633b4843d0e9ccfc370f19845cafc3daf19ab7f15703adc9a058ced922ab8252a2c64c92cb53d7c70d59ddd7c0e9711e1f59ccb603778cc165f4d4bff270930155d481b4f16fe728af7abd0ee17936ba2f7a741f197e61b6352e336bdb8da3c407fbeb60b654ab9fb125b79aa68f40eb15d58579c7cf7fde3ca5615553440e28a3ada65350c964ba00daae70976979cd4c42849448e20339888ff1fb54dffe203535843256db6ff44dffa91eac6f2374c9eef5b4b96264bdaebeb9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h13a0a0fd1742dcd2dc1aa86b82fd93b115b15c07ec585ea1f1a4cb7013ed84e4117afc71968957cb044bde090a2dd5f9042c887a6fa73a9869e069d9277925662b1c162ea73b36d942d54342715395bf8ec846b50164070765db6cb37ec647b743b75cf37f0d8ca537f3f2876b0aad67bc6ac22f653e6a79d5db11c67394e664643818c64539a14f1d9647ae8470e87281809c2a31a044e6a8fe65982ab10305a7f444104d973bd5bce3bacb07bd38738d05465a29cf9187024562cd90e31d23f924bc0ed937ae1cfe96fb3ab317b3cb8e5e3c13840215fe38f73b7a8d401d35ae30c3bad5fcb7d07b21ff7875eb5b1526e03bfac40a206342763de992174bd9969ad80803f4db59a3b8661d274e13e49eaf6e8ea35a2d5cefd62a8694e83e2d1b0dc4ee2765518092a9ecbdb042d9a54df8b7191c562116f776a1d513b09492330a4b07;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'had6efaa10d7bac90a4cebd655acf244231e7748399e1986d2d3ea3d3c061b033278cd4805ddc05da7e657756d414676da9e0a11fb58a4a996becd621aa045f45cc6edb14c758fe20d0bccf6072106caf9bf7eb1b644511abf20b5bf8c8f4cc41b3e453f1142c9983bb7dd254798269cddbd2d62b876b4585e906cf77a73764a2ec2b706b4aec8798dd6e030c20383b6d33e05b7056bc60a9e791a46c274a8b3492962375f2160e7164cc2426aa27939c47ff908ce1083b02571d1bb7d7402086393aa9f65d0419fc16fb0083f6d7dffad07c8e04f43c3cdc4f4fea1bbc741795663c5e56f93095e09812a98691b0c0a4c1dac816b62bb30240846a486f5c7b2bbc787f03b16ecf6da7b43ae4c156962d66f1478242e6a3a0cf317f29ca06d2fc90d2f4b8e34a3cac97912304dc9671125d78878e5a6be529cdcc542b4562e2cd4d045977;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h653e935b2b2d41710c4e8bf684e6123d8bcdeb2d7a08e6add86700ecc6fe4ead30cc45bde2f29825efbfa861616eefa18ef30d828e17050c89ecc8c2229baab3e481eca2bab0860b18727c48b38b8a982e0288c68882c469278c01be39dab7cc5f269fc09ce51ca6fa5016f3fdfb78714c4084fb54db4f265cf675c6362b9c87899e004cb91273a8d7fc7c3e2ce0c93cf0f6de5fd9a32f1a3ff537c5e462deb2a3baded98a78136d4df1acdc553f0bb1389bb6b500978ff14b43b3c7e88549cfe9b945e80c738f8666812bb2538e10f1f61acf28e2035f2340eaca3f2be0b146702cd5e6eb841f117e35eb5c944db8e1d4a41d1846d55bd467cdec560e21005ba88933b86b86fef9624604d36ab1d58dd93c508dd9be3e5068818363eeaa012b4b588b90a6813f8763bd3d1bb5e8367b0e37f23f78c043f75128b4d7291f6c80e8f63d0c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hae04d03a911f5a52ef798488ff45981841da2de1329681043492f6209c71128dbe8288ff205bd8c111b588bd181aff1ac7ea8f425f8badeabcc3451034aebae1a2719fc00cc3eaf1d97638df191ae33c60f02f3cfc0db17082ad1059558e10d560db7e05d8fb7d85dc03d629b96b13001dcf4d64b19c2ae68e884f5f4c33a37b14b4de4e6eedc6a0a8d119969cbe0b4d54cadcc85481a7ab09d5f9967063294184d0dcbd3a6bfddb8c74e06db0a3b84037b29d355592050018c248f8a3b23b6ca64fd7cfb741708270051e4696b89b18a2393f70593f9bc2a1373b286e27c8b393983476237902eeccaf2aa99c682ee349fe6f65446ec8bcc643e5c319dc2c6d469567d58e44e3ae82d167eee6b8bb8df32b80aebdf64dae8bafa378f5d6ac4bd85be0d783abb9aba028d44a5382584418cc8d4fc9a6c430ff12bac395aebc7a7f36f29d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h66112d26bc929c1f7097aee2ecc07d0ad321bcae3c058628bbd0d16f9d9828f8191889a68eeb9ed763f7774717b507bde13f93e88be8365296115aac09092d28e4ea4e79db6b16c4bbd2972294190d8d32e27ace5e7af5008bdf89c4942da593aaff18667308440ec7ef957b546420ff0d8cc3aa93da059dc1dd2e4ec6b9e24247eddabbf496759f0ac88ca6643ffa7b3d30eaa56ee8b59b01450c79106b4dd9910127c69f4daf105b01fb47c57ae753e487b58792783401552b6bf4ba1f1db5b3c619f4acc58ab702697bdc6916191c6b71db053ed91534ec887a40cc35ef8464132df5b36e6225b4855ab8a03a880dc57c123e06f4708e5a7d7c7a5cca11f94dd034e9bcf82b847cb641ca6f8254c3a03899a31abcaf51cb3d331a129e981abfee5185a42b9cb991952783be0ea51ed365e8e73c6cf8ce52aaeceb290c53154ce5745c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hc3e7f1052b278e2a384a9c54b5d187e87017951f8e0da79d01a72b32a789bea5cb20bf1f4e86b9a043ddebb89633eddd3aa0e0b390f53c2e8b5bb18d7868f7caee29566c9454f67c1e1b46c07b610f326092c6a8a034717f89628a6f773122fc312e316aaa4a6a68fe69308c2c722fc0e6ab37f652f1752c6342cdebd3b9f048b120be9c7aee5890fc34353abbc28d865b5725144fc6a8f13c7540639a6000194feb537e4fcfc6c7fecb02348253f130c0a4407f6524b7559a3216ac659d3e2471cc32c8e8859117d22cb521574b08c427e40ae3804636fe807d4cfe3f4ad1b2c226bef79b92aa42ee1c2ccb7d890cdb4db0c9669c59b8b36f4bbcfa7eed212835a28ace2b9f2853daa565d2dda52eebce99c9f5f23a5a22bcc62f9a1b8f18c20f0412b7a83b73bea18ed42b1a24745c1845f98157d56ce59e96f9de295417bba1eb96a3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hf3842166e3908fff355685eb997f7c57f18ab038fcd45009b822fb8b5993f356f309b8b91eed0815a9a06b1d39780e417d044de0fd65b36c7ce80dabe884194111b6ef48c17aaa9fa9811739fddaf16b3bd0ce9dd18cc15a1733f479676773664a735fac7da476eed7143871a9d2db4cc308ac76d3675ca9669ce6b7e58cc1ef88545058370eb4b0ff841daf8d8c56b2a2dc60a2e4f9033f23c560faef5624e218f5907ae05d8d2086032564638d884376c8462f86d0a320bc85fa45186ac7a3b767d88668ae97e5c4b78c82bef00e71a139eea97c6554d6e2d51ec2972267e898afe1acd8ded8a58cafaa3314ef6656953e77d1949447296862977fc8e2d85347eb11a72c8b9e10b2d02f008cc89f725b256c550fd211ce74746047ba422fc53cdb0a3ea44a42bbbc58e218896fc5336a7723af4fa0dc4cd65ee99975fcf5bda24cb265;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h729ac149bce7b2ed8488b299f883b80a1739429fc464d28e8aead5961bee935e0023baec46d5fa95f8a532b09e1cd2d1de9898f75c1748ecb2d43638b06c18589e8bb96c0da5873e0cfa1434968e32f74427bc35277827f961b17ab96cd88f0fe383cb6479d30f9c76f032721968ca9d4d9dc645b64c83d201456aa37b4f9f10031c74152d1d710136a8ead1d05df13d4dc27ae1ce71a387c05671f45fd0904063c7e9b7a0ba764430447a4a07444cbb768544336a7be1a22f880a08f29629a55141c386551bb22363828e7cb5736b7ab44f5607a7fa9bf92b1767e07fa8daf7578f0c5addc0bb2e1883500033c5525eaec9db592d3f2dfd5e02d0ffdcfbfe6a795fb0a8a86bafe895a502582a1988d25349cd59f485cfa87002bbd020aa55eaf99c89a9ba56d345ad118413e2b51e05c579c617b4d8680d4355bc0a87928022106653a5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hee0d08fe369bc6f33a60f9b1875b25d10b92d27f94dcd907b16a7bce51654a88a610fd5c6f3940419e4c82ffa230fdd6b2592f2d2ab4230da1787ce837030627c0dddc2e80c555e9f5af53d45a42d4109d67d5d75847c191494f9e195eee658cd760283c016d1173a3afa81f58f48d10243b9b65635b1f0d4fa2abe8d36f2ef1b886e10ad06da5f72c4e51ddbaeac5d9426fd5ac95339c9f940c7c6bede8ca4fd060357373e4ef1ed07840c7ce05865e250534310c83319eb6350f2044ee8c2c0a01112adb319e367550ccf300364c0881161d89a2241122082637a6043879ced25a45e9418513f2ad7c9e4cb07c995f69f4261dfff1632c5f3f938b91f57c59cfd6af8283e873966fbaf548d5e18a23b381fefe2d7c9ee0429b9dc88367b3bf026926ee7f42d08fe0b55c03a720bbc545e4a34c61891fae9f2809c5caa9766c0647deec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h87eb656cc14aa771aed0dfe089e94c327f405c62e3a296b2b5a232a1bd896b3282f4b4e105725dae31e31e0286561e7a89af138e5c565e625bb93ffcc83ecab7528486a889a96203b19667966eb9a2dddc5daf786b8870240d64235b55b492e634b7aea28c9463c105056dc45ae961eb204e3a9cd647fcfd2307200930995e6764867053daa38b19de9aab4d60c9892a77bae9a9a0db4ccb76e814758697fa9f305b1e83a543f94562a3af5a998d814f84951efd63b2e0829dce2f0fbe70c3deb14e0eee37d967e9f89def84f4d1b856c75d9e66b050d6809ddea195e40939fcad07544bdac1fa8c41970895be0d149ff35af4acfa3caceb7cfb214a3a121f63077cb61d668a3321be8540441449c962a1cae62eae9a0fd95ec9cd70ab2cfb510944b58fda9e4f164e293a476f0ea1c8767eb9f27c79677af231f9458af0d6be80580e5e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hebb8fd0c2614f0b3d71e38918bf235198dfc53c338c55d724e0a229f49a5a3b9956dd20224aaad5feb8681a60c139e8fc105313f30a4469504502ec73e80d9b53f8ec8ea8a94824e5b644ae32bf6877d4398b914ef7c71fc76ddcff44a2d19af318100fdc36e2a821a6af97c44955ef60aef28b0685328405de371e05109a215bc0cae88efdb4b38e396acb54534a08ff63d00fb10d365e4ad4861234c7aef4035e546a6716d89c411b07eaa2fa8dd0b754e42eb818f23a754c3330cf5a364333dfeef752385b2f4e28fbc083884c12058c481d3cc7bac9f0ef689d45848e2e737855046f8fe76bbef33d8db78f115b83ae03333a0a98d4c9ef9d15dfb89a3124869844b423a2d8322205e64025908d8ab1c22e82c32705abf1efd0261a1d40851712e0e06bc33d651a69f30e354883acef1623138052b8083995318f24345258ff65ac3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hc7dcc8ed77125e5cf612104549bd126c42ae5d8719309b07e9a412769229bb37fc822bb3e08eb1b4cd1f951faed9044bf34fc9f9124073dfb090f15235ba6e155a82475dba4e5e08a9dce7294987035eb56c6a5ccf801f6cdd01695065d542e34f34a720f38b15c3bc9d8e4d046a2498d11d316904bd43cd7ef84218f86f8b47c5bb2e94bbf99b020d92ea4cff478a393da4fb5c31f8411ca1ccc910ea2de8cda72f10ca36d4a72490a1b86c6be6f536f6d0ca8d1f48eb59fce0fc5e6d438336d30763b53ea8a982e71fb12fb37ba51f0ac83b0a3c481af77bf30455e866155531a4f83a4717bb5d4ce631a763169a8558685bf489668c6b466239d6f57d97a4efdfd1bc92292fdd445d6efc299e8e3903c9ee96931fd741575b3d2204c2d58b8a3b8cb74482d80181bcbb529d785abd39dce8b442e2aab17d74a77d0ae61bc8bf58ea83;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h44a3d52b39b179ff63d1aa2136c40ac3d6f4a059050dcc4d469ba39c8df9d6ee7d80d36497f1e56ab83335a2eaeea062b49f9a2834590a59ee88182fc8223df372fd428211b690b7771e01185d48497823c075e7b735eefd6f9e5b2bf22a16e60cdac430132b4bbbbd2fdff48434d14bdfd440dce6de26a317d9a4516d95b4057e5e6bd08759ebd97aae0e5eb176df4effc6b110cb0658ef38638094ec7d4f08150200e1a597e4ea33a8f4d78ae4360db537a23aff84abc649e8288876ee244e2f37d55b793bf6c3e8cd3e8a1ed29f9a2ff76acf5f5df8ffcd1914956bc84bb41dfb320aaed12791fae9407dca15b163d156ca7496eba86f4ab269275155c4da0494321df962539c1c6bb351bf42b5fc8df4d3bfbd765fef6daab9e5d922db852bbf11db2b23a1f1e0e4b52ac4aaf9d54e91022da839d6b79f819ffac1c5976802ab39ec;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hf2ad1d6337697b9662b5aab519e2cbeaf83b19ad68bfcbccee154fb2bb1b4a3e7113ee76791c8f101cf9c9597330c4038403eea1207b635dde8fdc8b03b40bb9c8e35122a7a0eeb111cbf4f1c23a8f4357e97f25e55037bea60ada7159422294c7837b6d87f973e93d0dbe282e9cc023969c017c991873f986b4049d87fce2e775fd71d54016e027210e24a5b97f8db1b6ae2b91936e63ef629b2b77ab55fb8dec5af27d2bf3c2034fc1482d3c948794ecf7bd66336adaeb96e19856136dcb051ef5f3793bec977dfbf106a901a6c554e3ff90820ce1c403c1e4639a19287c809643981ad39cce5c53176a81e4e79561108ee22e3e1f13102e549fcb95a92fa061f8e87347f6a8335911ffdd37c0e39e164709f7c4efcc4c72a4474c1cc2307112806d02334be801b213773cec5d5b358985f6769f21a61e982cb6e133a17ec3d080b272;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h8c811a3461cb321033257060d4911637752ac1f2354489d276ffc413b816665cb3829e7ed015ac6c38372dbaa6f1d8463364755ca74f0719ab071b6a9ab12aec373cca80edc9ef9f11f93734af3997906ad3fd004098739c3aa12d691b5a94af607710e57886dff5560c059ea5a7bef9fbca195a6044f39e25f657e754fda06bf74b1f6ad2a159db36efa812ada12aa3881614e617690e22a5fc187a6e780ef454af6c521b6fc4f27f044d4bb0a70a89829f664fdc47e4365006267ab923f9b25d0cc8c1a5494185c8dfea3ed5b73ea4e58ec77d47c4e3e79d079ae60e3e94e2006f1e39a432ec6ff1b65b04c749a932336761cff6e266ca0a4cd0ded5b48afaa74449033f243cb16b631ac7bd5bea8c952ed3056c0b04565fb9bba8bf51a8a67b90f113389031f2e5930473a37d0ae34f20b59928727fafbd0338d657c81182373c7c3b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h8c757ed84308b43831469fdf9d9061415dcb05e240a248fadebc57315c8cb43a9a0cc8ef85a39ac5f920262974be736eac7553d7edf384699fa27aca8d3c3b17c25195df549216d947db8b2f835d6615a695977d52b26fab72e175cdb609cf07ffb76130fae4e5ffbb7e731e8b51889dbaa6d6f33e0ff322a41002b717d5969a2c5456919efe23b9be8b5c8dce4a29d12c6908f7510cfc1830be0040780bbb24642e2184dcd4e16d363e77d4d9f7353fb5da444c89004884accfac8b13a84b9fb106422d50c46aefc29e4756dde9380a3da0b9f4096c075dafecc08cffcf2c29bd790fc4fc117f4e2bc99353d2c638f46a2adc6124265d2ed95e77e8ecc92342851202a60d0d7aa444d0b65fdd78c72f9927e6e9154cd2c74502a15ae66f0a2d40c58bc2f95f4accc7105f165fb8f16250e94c08d931a6c81a58d92e26d3169cf8842275;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'he7b8094d18ec7d5ee2a08f43566c1b188ed59eade54ce3e5363df9e50de8849e552e0931b6e6a933f7af27acc8f15eae87493cda2004a14cdce7bd65af679b6557a5673d1d0244f47642fad86394387383ad3cf84c2c1d1638030dd4d40a0e141dd96a54367580c834f6c08a4ba9cd5f4309218ab09793961302a691381b49df309bd696979390b38bac9245ede0bd8b68ae54e4059834616a665215bbb8ae511d04d5e0dea69b7cc1facb43153a66d0d3c9b8b0cead120228c48065541dc0be4a6b5c6c1736ab993bff4f786aaddf851bed80037d082fbe915779fd95c1317f7bccf5e4fa30b5c5a91f0281f5450ae01ce153ca8cde4061775d4ada9ff4b67e295512356fd2047f6d3eafe36c68c13240acd963616564df75870000fe992ced4a56537f20a8a5315695d06098e900ad993ce5469e0f8019f14d13c25f660babad7b2595;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hfec9698be8b3e7e08e7e0c385fcd8e36e826ca4bde27551780c6a72dd71120234a3df5cd6f6ecaaad28e8d0bb509ed600d5b80c3fca326a3b767c530eb85654b81d83b08b9c687c435756ce47babc56b4eb3c43ea5449022639c41cdaf2d9fe0eefdcf8f15a923a337f59660a8b6eb480eaebd8c0502f01d7904a2e2d8918097ae8b3cf2084835dbfbaea5840b3f5f067d562a734d3a773e585962e2fd28d355ce5c9615ce1bbc9eec14d37540150a9ef6d664ca725513ede14d3267882921c54b81641f2c104b04bc204200c376ddf283dc18bd2fd815e160eb8ca87c98019c9d34e6bde673dde727981a513f2a9be98ca33f3bace6a4e42fb9c926776692a979ff74c6c2eb30c6bf34fff1162e173c4e3e368704e62e1aa900cef77855d7b730f1698353ad4e052ffe08237e0002f4303137f3a02ada7dc3b07928ebc9b1fd1b8d2ad5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hd76c12aae3536ec225e8857816e1c90e6be7e65dba0162926607a5a7e00ea60ce55124ed7ce78bc3438711d02880e5eb04297d7a741c8dc1a31156819e479ae83fb794371ef73add0074d2f671672f841eb8c7d4e03615cce508b32789074d15a01d69ef475e6ee4d2bdacd3eb171b1774163242fd82e17f5f0d7a00c7349b1ca4190491a2b7cc870eaad1b16fef63d8034d89664f6e303e5ede5bfe78d0993966c1b0af191ff6ebca1572da8f0b0be9f19d9ed35074f2028274935467c577c3fbc78cc5226473140bfb92322da00054232c21e4f6423825fe80ea7dd426c18f592b07465b430f11507138a059d84bf357c3e0697c498cb68d640dc50f54842e919971fd915c933fd437fcbb06e1389a03a090cdedc355c99863e7822c334a84d933af27bf327ba2358fda8dde412aec5f0f9da150e849b070e0084898e3ca9f252cc4a2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hf325c4ba21fd52db0e4f98c11374bd76ae5538c78376b9cb918910bbc0874dde112bc8460ab27beeafaa9955c6b7cd5c6ea3f0b47f899ea0354590a9cc5abce7de086e2c93f0717b23ee34977697db39371d115b33b9761c7e6aff007424b9d8022b7ed5a45c26931e88da6f2170c16875abeb94930ff67addfdca0d5c7efcca0237e8739f18a6215200124d05c5b2ecf8a9dc51a82d55a8dcd81c028314203958dbdb7287aa10f009ca2cf9919f51ff6f8b63b1697adb8e9ece69e2348a913d0e8d10d94b55dd73d4d0c35bcd72c7e7bc7158d70cfe3a48f9751a3da1a5bd6f1e73d47b922d07a52fd1b0dac7c4e64e321acc07382ff3b0a0012372206c26ff63e74e9118ea2f78c5ec8983a5dc9e5da204bba44e798ead10404fc1f2a82a7222a6960f2beb17e98cef7dd815f21d9d30ef1192e04a6cb3dc736efb6338428b8a9aebf8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hae4249971ffc89506ae854ca04ea7a30e79d8f05aa98b36b1ac82f6caae0957a558e86a85fad0b3fed411513f9dab6b78d47496efe8e05cc06f87fe92b38857158b34510dced66fbf54453ddacd7b755777574d38e880d4107eb4c08b71f059efe45c2d65eb589cbc74a584b4dc9cd10de7618915b5e6a366dac39110d6989afa0edcbe945e25b96a0d41f9ba955a89bf7d946c8680efb539e5855d2535fba6e9789aacd243f218fd6110b308cf81b7cfdcd1c973900bbaaf53d82008c02083d92994eb147d2768894119eb02de3a463c30613b36453c94861ad8edf0ba9f912421a566056cfc87d0bc8a50198f86ddd2308f8d914780ba006b73ee30d2fd6bea42e33dea3c3429830a715fcb73efedcc678563fa68151500fa0eb4f2954046ac04f74f9b473b4fdf5f730b5427650cc902439ab8053f8960241c2941c40a11fbe9d294e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h2726a0ba2c4ae8a1eb8bcd5d4862769a52255d4914255d06fdc4c90b06bc208e6b5fc8485adf3c4aeda4cd0a991d404a9e4bc711633ee26a112216bea9f90677585966e4b449a2a03e23afda6c2250411312b236947f0613c031fd289efaf98c1983a67aac890ba3750f9ee8c07bbdfee484d0fb8fb9168fca89b78922423d2ce46d5b41673bcac94664ad1947d13153039c50d4c308b0f00772e3a133296fc38f176719c3535c96ac67103f25b56302e0dbb5d5a0494b1ec121f19fe34f608a90af9b82999a16517393731a60b464b3538e89ef88cd2554a49d53b19c387bff63b60fa4ebf61c809a7ec2d804e011e89b0ef8a7edf97b2406a7477a927e3cd6aea58dcdb0b64464faeeee16ec5fc96d80491acf88ddbd84e827afb3583c8ffd4d18828a4e00795473c4fc185af9bbaa843988e01f5ec84662938045c0fa6309f32f8473;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h90deb566a5b8d436c5648a39a2d1e0e02fb4e5ba106b8c4363e5d672b85107365b7ac202b62893de9a39d19613e1cf4f01daea3dc2b24b3bf0704cb726bbd4edae1fd00893c91eb2c7aa45cbec741c9f8714702cd1b06e6b06ecfe45d160e4aa89247a33f7907477d46b6f2e2336dfc4ba3d3e0360966bc629bb013ab2f3db4f1b684c091e5a1639e0dbcc4bdd2d22f6fc4d704162ab743d581efda7f20257547b745ef9d76dbab583b0fe480485c5f754387904aed7355d500166c85cf5b653595c1d030ba199ffb29060e1021047aae7636ad130fc472c577304fb486e15576085ce9258e969c362a93003096f8903d8d72f950cc15be726d67b380aae122736032c0b20c9b13f47a9c0423cb7fdbe807806faf7b80fc0156237b89d74c702690ae8d8d625c73bf330c32bc7ca37b25998777d16848b41baaf33873aa5225f6fccaed4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hb6b1bcfd52b178ded61fd1af84aa485d0140abeebd4d5260caa2900a143d05dffe31519e383ec5bb223f8fff12dd7d4f3ff06c186ad6c371a43bde9147b610d3c9c6f87184f63fe9ecadec7fe8baf491b3f70ab2d527c23270123ec1a81a8dcf561a04efe5f6fb29a53cfa212eb4f3affc1841e57ca4ab3f622fa9b2be19fd7a985c68d41b84b6b35af99ae693de46517739339bd35b4897192028c158f4c9f8e89b56576655d42459747fc7433c1c2ae8ca44d0e7120637f6927a8cf5164a7c6d35731664d45736b7ed6442191c4ba2dd0b35ea6862452b419f8423debc2c30cbb518524fcc72bc7c88c77d26bca36426eaaf4ec23ffd9d099623afdeb8f99df077025fd4d58e026b30a291e97d232d5bd1c424673f4d3e46eb74cc3600061393d487d1d0ad92ae2077535c6a82db968015547902aaa0eac15eafe7a5a9f6eb94731604;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h2171dda551a49bb28cba9a68ee4d18aa94c2385951fcc5b85cae935fb342f37d133b1462e6d11253db786e0221ef8ac184acde1bda048c948c5549765642cbd8836edd08108b4d9623c4a646ad565f3ad8fa84d062de1bf8fc5dc3bef809aa9a8247e84618ea116c62e82b1d1f908305e2682da280456a82d8e7d9e81e4bf833895bf0dd27fe6ce737ee383dbf787c3158146b12927eea663a529a931713254150206837029a9724e64cadea55fc00d816261062341c7580ac161bf9b8712c1aa322f4ceaa4eb462ca30ee89041e5fd5aa9822472b79e201b015846701d4e8a6db4f6c10f9686c729ac1af5262e3511ae7b392af96ca7f3b89814e2870d786ad817d67bddcbafef49c020d3d7190ca3f01b65bc69b716078ce2eedc158ea047e6082c9ca884187ee17176c26ef22d8cfef2576deea4529900ab8be530bd9e65b2bdb1f83;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h147037cf013650cd2eeba8778c33c0f5b3376e969ad69c4dff58fe9d3938379dc4a8c0d27763856f315838042551512e743d47a39c6887428134cf43685176ec1d118b665590558c5ed043f155d1e273510bdadd4e98e7e2ccce02a1a2f5e7d9d85165622e6f1ab1d9cb7a4bade3d298fed99a7ac46869dd8cfd3ea84c831893f858c7b6cea04a7a4b9cc5ebd7670f3f38f15fd8d74f55522c460760f2a12adc8ef6a838166b73cc768c4a894ccb96371566e7c74eae0121d96244da96179a6099642f5e442160dc27cf1b2436d7be6d38cd8446dd129db37147aa269e793fa64eb2edecce2e17605c06c82eaa16d28488b578c2ac23ce1c28786e0f91b6afb423dce58c2d99602abfb8685f42e6c9337e2e06378205a625d845bb4749d47bf6cf98309f2ebef127db39b149692522a82ef95760cde3f7a1d6fdb6d466ee8ced69cbfe8b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'ha0cd9d62c318a3751f97a06929d087c01e7195d85e7fb737f810b20238fa74d04ef0bc5cb7ae2f286bf4e085852a0eea391c2f8d9ea89c590c7b42e686aaec7f2f03be92cc2a5f41b82b13b93785b2c20f7fe622e8633e49b78f6c27df5293990b0ef994657f55db02b640560a7ab0442e261540b33bb591de238bb5ff850eef9930a2379255607786359b42f1b39b3896f1ded0ec3ea347ff67a549923754b197d8061df5215b705dc67286707008443edf6e0d1afd7f7eba1b306633b3e00586ff509ff9a9585d1b77f71abcfb67403db832426b35c59f16cd64ade0f9cad55b4a494c65603336124466259598206e6cd64553c951ccc89aeae4cf1a816495557a869e6024c9f1a26268394b0d8c558299bb58ac3a0011e0b7de14c8a3ae14639313dc31e69d9a16d54493aebb2bdc44fd95d2842440bca13ab3d8a1acdd66bc83f88b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h9975931cd30d64a2ac5b0ef17e3a6c8e7b8cca3f0e46f7c49413f18bbbb437937173bb84204013f132b161dcd882a32f9f60801d13ffbacda37867ed8bfea875a74a4708afd0c54852bf57a7ec3c4c68b619ec9ee52cde1fc59ca614925b8bf5c8fc5fe50bdbb8f5a3ea8bf943cdad50b2068586c45efe2b3a4e9af05176b0d3238cce59fd117d460557630fc1af7a7d48db8073d9bc7909cea430785ae7af3bfcee8012fe713c3a6b6859696085bcfc295d2e68f873cc05b782036cca69b2b52e6db67cdb693e4012f59f0ece3bf695e94243ab5ae9760b650ba962d68b50f5d12370183bb8f1cc719aec4dbfef44e1df0e050cd627db3eb12df20fc404c0f9d22fbaa835fcd36fa7de41d3dfd618f0af4667da6557cd2414f39e899b1b22a3ad37afd27698071df561896eddd9d2c25ad48b90941d442a9f73ba5b59406fbd0d98531d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hba1799f21e4930b19e53c2848b0ba0c38437a57849a4b8f4a4b8800f39830d9c12e7e4e54d2f8c761cfa5ad74f31e2bd735890d9811a22a8b1fb101e299c5a12be3f2388b521221f1de9e9e8ad6b9e35973be8ebe99bd0abe75d87f2e4b2877b2ffcf842a92af177fd899acdbce4881cbd6ac447cb52cdea0a550f023445e72947428cd2fcb0a634fb062e1d2568e9e76ba7db1e45e36c6fc7ef3aeddfbbc276790687704a4882e3672c7c1d7b713e6b7d89e35bbf8beb4feffd1840ad58d6d1a9a2ec02ad568cb064fae50d3851910d96dcfb16d0f0b93542cedcc51b6a81ff13772227c38d8b010d576635032c7c35acc51cb085bbe77f8f3f0a341ac6ac0077cd786207aade93f58d99e317085e64e8762d90fb2e1efe767b30a9cd92e1799c606e70b13549d1138e8dea165c391cb5bca4c3023a36f55ca8eeae9e8760060846af76;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hf06b9f51b13d978aa78453d5be90803e38a29a00f692f79b04c0899a268a9d71fcb040076d84dacce16b436910f3e81152d4b3ef63786a80dea84aa59738fb3b1d10f2d88ce33d7994a1366224d2ae43137974225d7a2c6469fe977303303fdc3c948ed91d19ac2c6fc2250e68f69832a15f13cfc6ccde42e045f2df0adf6f4c9dab5ecd752c4264d8ad0c9e6974d1e89ad6d11128cb6244c2fbaf6c24f7eef1cd01dcc2edc1fbc67c2813d26e213e181ebc184cf3ffe525861bcc1f3a617e745ac98c744d7e029aa4b6c3365fe6911a0facdffe37bb95239adfe6deb2096694c319f260f4f46cbe36adafd016ba05666c69a5630a4952cee84108675d1430fbb42477da7f676bdfff5c84132b4a9e9912267fff9005acf6db18d0016fdecb4b6eeb46f8ceca6487503ec8a74c07b492e375649565e75e7080714ec41e00ef4e032e8a88;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h69f2198a552bad4b677615cd9a300cc87839eb5a1497fcec20e59b1b3057f4958bca44978971ea9c6aa91f51decaf60101d381587b4edbbd093987ef74eace32259bbd700b55173f52a67fb2a8721604ec8e7cb5caa6a96d32766196450b5cdfe201adb7bbdf8bca6e60d6e6c46c6c83382c1a818f5fbb1db0b99d9bf69c9c197ca40e73a85d573789873be1fe08da9bd7c27ec5101d2168568485e1443b48d7336df83c8855a39bfa0c8cb966309d1b10b2a397304ec814c3838c96fd9299427d866a892ebf52068a873b159ff0d853b9bf5923101b1ecfe8c5db9303e163da235f0749d541b6bb6251243463e36ee4d069ebc1a127f15dfdc5bb2e71edfddbc71fb15734a00157344419d9d4d6b7b539f6ad32ac4abb092c04def241d4c9d0b9286ea749ca39248dfe8de52af29f3e420e45c710ac092a3795f44b9fd0815207af2f03;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hc5125d68b4d10b8d2fcdc64a7514245e9c39dd25cb8269d00dbebf647ec56670cf2defc07ae45fa1230e1d72aa86c0baca3f9a1b24ad09198a3d2c95065456adfe8116dbfa3849944da12bce52a8f2f05ffe22bfe481de9d4e3f7a502ac866f60027974eea427d1d178ff5035bb2c1390b1fb3189369d6acc077bab27fd44773b8b55804a3c4e31bf3fe45a6cda9ebf130a71e1d63954122a66d293575109f88cb7cf4e0296f4c71e17df494963e6d3a1f53428006da2b5b39d4b4743c999b98f108fc506cfd40f53024c1428762267e69916c48296027a6ee371de16687e18130b1c587f11b6986c44865bfa8fc4ccfb2b7c8421f6002c679468c4a25813f8b9885bfab05c9844c29455fc686302d4807bdb8cf9175d8aec3c7c540143d55cc5e46078734ee4ab431931d417c8660aa6167b854e6b692fc0ffbf1673710e2f79364cce4;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h66b08d886c2b1a835cce4848f61b49739909cd93c1d3432b0955806c5e01745b9de51c84a492ec557fe3c5a37290ba99f3a986babc3c5120ee3de73bda7020e30718cc68dcd324cee2fe5c35d89d46e0c83a5fb38e72d932411bd1e7bcfc7c98a32736229e8aadda32630791db7ebb6f2514c4778919d676cc60ba83f7cb5b1c1207b58179facd9942f0cb5090ddb6240783e1323b2710e847754efe948dc715e97bd0da9303537503072e708e50c354663ecd35bbaba5382c7b5d611ccee05752991db41320402f7a08759c42c76e46069ce9d91310448647d16c29902fd70416db0ea675938add7e74aa5ac4a6e216eb2097934a06d4349943baaf7f12f379a6742940f96078756c2bf117f40fbe2b970ab2adcbf57c505ac4193f8a16c291a43504decec46fa4118df169a2985072ab5fb03113267aefeff6d795eade33be6b9d71c6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h34337efc24f62ac99eb990db98af5481b111e19565888fedae1f9ca03851f9074547d4383af8347d29b417c4f2abf63793332fa87a2ee536c53abc68a3201986c05e288788d95ec5267bf9a00f89aa83e94ec7f71b0cc48a72484e7ba760a4c62c46102e7dfcba847c5853f63c98bac134e8c663d4142d1930d046ce4198e484e8c95ffab6bb02ef78f3880d29c8a01e0cd06f5e1bf2e7c0aefc58cd615eb44602a41f1b2d5bc1b13809162f30d0a6f2cef0688f3f4e154655759b5cf449b78877e535bfcd655448c7e41f50676be9045395feff63bfa5e3b9abedd9a2e781bc56554ac2390b0926e6bb48ff1860c3be83f137634ffc9486a7a087e1d265e1d3942492c92a962c47934a2375436615d5a0280461f65bdc4071ea48af25c92b96ed2d488a139707da5aa89ddb5e08a04cf30678042caa8855d27e9fcf9313cd59d56a0599;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h2ae596e883dd7e055c19f1f2e5e54c4e99a44c26388396c61cb357813165584238f831dc9c8d2c55638db88c54685889fe4a62cac3bf742b8570b03e7a75e73a97a51b3d8880faff1451880071ad0c5ec39dc7b407d0b59cbc92345ae52b2fb00003583511ff33180d4998d29a91b4be428bf111a5ff6bcb51fbbf01ca4801cdaae4c8c16e54b413ef04deef5c1ab96961793fad97cf6b4ad9d7c3f5b75c7cba5191c77d3442fcd63fdcfe8e97e04da7b1a9f7a32323b14f3c9d6f296a63519afe450b92d5a41b31c60ca5067b2aa94ad8b646bd38c65a0f5c14b4791089c7ebcc8947e8d2018a74b0b7cec5eefe4a2cf24871f58b8ac9d4810ef29c817337edecb749e3f8306672f82f04aa0938e37b601ef4b7a20efea6776e6d2ed5ac1d1e29d601b2dde46a7c293f8d383ebf969dfed9e0ddd89651bedef20f950c24a70461f9e1c8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h4b3f16a8ea33b6ba23be003b6c5813a6b59a5f7849b0414435ecb8d910f16bd0abcf87f8e8f4ea526d91684414acb90c9418d74d33ef96d8983c89c915742ef37ff485d8da573b20b413b8cd3568cbd80a2c2d8d7564c88f3fcd38076fb6281d2260d8cdc182c113259e697d3be775b42c83f22745355ac1bde0a002d85648902a37a1467cfdc5021b60a1987fbb4ce3e6cbcfcc6ac7d687431ae83187c2b47fef8dfbc69bb8a51bc857e86946f8cadfa36727320624f4607a825d9780a8d9dfb88cd6afd2e782fcaa850b76f372e46be334938b041e0dbbe48b4b0777e7b74162595d488969000a0e46b7f392009f163686f5618df0cec76e5dbe4eeaac910678bc8da0b25483161f078023c013e2d9946ef412709c098fd2b77f0e58421931709d037930445ff4fb27ce5055f9cde4e36702848111758a4199dee5baaa99d6cf3d35b1;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hf0925ae1f4394c44b937c8d5061c41f2308a19a6f3c6f2ef331c6b1fda978992ad36ebdeb53520a1b1f3085bb5d128da404ccf09a4e0e179d68d81116760cb51e2b9878b5e3eeaa7999986c5ca50408e6a9d22a52bf1a3ee5ae91f40377494eadb08793474fd3282422833a01143e82d1d5409f7cbcd592d3e1b5e8981be3a7888af3399d0ea11805b9972ce6e7c61f55ca6a170f27122002b1bb9002e9778c5831ab0e7efde8f66cc8b43b244e54b45f8e85339d189266ac96231ed3a5d8029c4d88131f2ecd44250431c64725196894579dbf45c026a70c8cc04f3c502dc13f58344a6c9b1f4019755e20b7ff87dcc988a537173f6f30b8a63cc76cbdf9608c1e4b6fd5f3d7a8cd021729d6eadd076460e1dc4eea7c7e7e8873f718c5567c4af3ba37cc1dc76de5852058f0435698f10f6b6eb3c11040d8b903ac74802b9224eb28e8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h5b27b5489dc4a29b931ce11776d628414a437e7be1f46342a5fa1d8f56222777f6f83d36bb1fc7c6b3167058a4a5320753935e380f30545c42b1c6d77a817c6671bcf14550752821c3e8ef8d7d8ec2eb5931aa0738f98b1ba283e5369ddd95fa6a9a350e9e7c43a9da4bc8c514facb9a896008c6c17bb87436865b6b0048d15d9297f728d974db449d5222b3729020787e0c16375a70342266eb70625818b50d7feea29afdfe2e73060616524e3b9586f6d9f381c09ef77871586032b21747a6c0ad8e5289db5682a392e9ceb8799d2b62e3ad32863157a087d2b3792b17ae3aef6243a6b035ab9f940ecbb08ad6ca935fcd79b04d2d1dbe6302593351f05a2fd8a767b82a8b3681905799874c3ccbcc6d1bf69bb2f525abe9eab3c478d436854af26b672c6c9e9df0fa5eb039eb2f2d7754e4aa8522dcbd31303e1c2af151293fa2be4d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hd846af8af07772988efbd272987cbf49aed7b9b993126400e1a251f59410a398c8d0c036b5b44d17561d8b52eaf84376642907a168b6941638f79ca476add15212dda19aac7105e3ca57e1389f4f2f4a90ab3255134c80d986bc59da30ae4cd33cb542da755bded39d639f855ee940916c649af1428e2749e6dc612af4c60528551f65752e19b7dfd3c3fd5ce31d2101ca53567cea94c84e5989c92cb23f2a53dacbdd0e087b6a3fd30db6e12430a9570dad6a8764478f424041380062ccaf03cad9cef4742e934c598626bd6715da1b303923f6758425f4c78a4fdad1d7e38018bfa29c7057e5d5bd9dd4248f05ae4e4b431a0874a34d71bcfe84805ff08521f3140312ce3da3342f1e02563ba960550434264b9e960e82da2c997a2930a0fe90fbef729d2de52c5b6cc29458ea63f7bbbb6ae81039cfe7d7f42eb75678143402769599;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h270111cff176407e91f48127c1a0ba3a6fd0cd4d14e28175863f0483faa4c3aa9e6a9966c6277cd277ddc3da15c40a242c6ed0b4e1d380c3dc922cd02e363110289c9e562df0e45da959778bb77dc0bebb11ede7fbd65989a3bc25079285939e000e8a6e3a643e21d2d2c80d8523ee5b698e42ffa3ded2b83f6f769aced0071ee04ee9664c7e31e37f73cd82f4afb5c1dfd2044792fcb2745ff313b52858207fc339fde5851422ce606411b32e3d10f7d923b287f55b36200f401674a06144f88ca2da9fe933ae66fecf2cb9c7637cd2906997667f587b7ae80e2fcfc7404b3f2fbed1ea172a8774e5b764d65fef029ea24479c71a68ae9647caac2ec5255e69a59df27121dab1f0d528b65f5d301bcfd04eed8a8b7fdffa485ddd70d001edefc615460578986324b0ab517bc58dfe15aebab6be0f85f8dc65d74966ffe8bd64bf5dccbd;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h8a8727057d660b42785d78849dd256cf1cc2771b7443f086dab4c76a42f4125a8e38db58364a58c629331ae6db10adba04222c333275b590cc819e0201b7564b5600f816e0bdf1b8ca92318f3fb15cbb7da53b776ed13743ad96d682db77e41d872a86b9db1a0eea5a5eb409dae25130213ae924e14ccbf7644492ff1046f385040d055526f1861c4124321c899e8262eab467d312a00415caa8902e4a9576834d7d588f08d8e60eb275927726bcf670fb7e34dc2fd65dd78ee61661fc97ce70c88617b2440300b47ffdac714b7a8501e336a05cf54bbf0dc24f324b64d6b42916ff9627f33f9568108085b815e7b8273f22fe80fa9a378da0872342973cc931bf3a43cf61aab8c81a28190cd2d19f2df98463ffecb58318f799be034c604eb3527561ca017b15decf303d4ea68fcdde912de141b43b0ff9a5091b0b0c10c323650d3c0d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hfcbc80639dd1b81999d2929fa155d3f4fc6e586fd403f9e8a535a7856c2a08f5e08ebe2bc848c46d73a41b8eab8bf36cf48293249d2526be97520a21a2ecc91bfef8c260f77b8815aeaf754f2b8cb5a2711b2929932a5504665489175b42370ce9d14a6188a47a1cb5a2c281124f54b77953b93ff0a0cb59e93788d68e3e3882c2ef97cce30065c3bea7a0e6a33faea74c73d06f7302b9191f81f194cadf23aebe981e852e328ac54081c8d9f2e23360a19f398eb55e6abd40d8e715894e1b94bd7a6624a48c240aed4838e03872ec12443fc20d2755754418bafbcae35c2533e94ce9be69c1959656fffa3f6c6c9d101fb8e71a7ac9fedfa4b69d51afcfc1a82f3130fc7041dd6f2bdb3b5af604edebb9e9fd3bb54d72ce4b8dc22d7a2f1bb892df155364735f33bf75611104fbcdfc5fed989ac4d679e8e62dd8d86d69a3b997057407;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h330602219c409ed693de251df60bfa8b0f62fb743e86977deaa97078cbc19fd1b5205738dd02fd33d13356b973c3e9ea85efde64aa5146fcd3a19791b8166a018a033e58cde7b12b9c51ed1f1fef5e07552a684e0b06b5facd40813ead15971ff38d9a2204e83a36653bfa4eb94819b749fd677c2051fe55375e6a8f5bbde0319076c82f71ebea4d858fd86fac9ea0610b068f1eef6c4e84080eb8a8808648be65282d9acda35aeb401b807789f5595dbfd705a375ba767fec3cc893094a96edd5895cb4922988cab145c42bb22ca203ed021c321bc971b4d3d11cb612900d212dc66013c34a0ee60d17ead6f0c88ae488d555bb608b0a773f3caa60b9784b798e0ef5e13109682c6d46232fbba7dd72190d654bc5e8a7bdff315b77905a151762eb19ca3de654145979f7cbc3c69c95ca6676d8b9fe4a6dc35052950532d655b5e9f5a9;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h95a38a972d6b3ac5d62d20d1f4ca8722a931353f8e30295854708038dcfc70a48265caf34e116de8e17a95a735b0604c7037d3af7cbc48aa220ea4f23dbb4378979d2c646dfd6a06b954d5ef3f7b062db91912130029b0bbb63a906a9ac2c80088688a20f7166c4b6f7fbd75914a2eb013b6d8a3fe8ad2230d4a59b7ff373b4ea0a013ab2e8b80323b63bd3d10011ccb33035c406554a9724e5a6f0b624ca188d6a252b8d23f6a8d7917126ed29180a560d200292ba3e1d9d3aec001c095cb6073fbc32d3d15afec1a0ecff2b5f1ecc414367a2c26cd6772bceab737f32246da5d11a19b4c48572047fa97b3584ea560aa95e9422ea96b5d634e9073a52619f02425ea8d7130a9be821b368e350799aeb608c1bfb73483af043e1ab4dcb3401a7ca7355613aecc1ee8067934c2005370e29720248d3ee60f8bc4ddc5defadd304c16b15e;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hb0d02e973824723c5d74fe159999d2f56577595df9b6eb77af8a3522dd5bd02e37807b2b964f5a3e8b279f6c42f5a9adb9f3942580ef3f341ef9ec40bdbeb828c60640eb479e1065b1f8d3c10d9f7fb68bae14fab564391b5f683616947e8e1cb806e364280eb9653fdc29341c82277b345e05e3ba1fc0faa2209ea20522f578aee7e0942bc800d1b981ad3bd6849173a774d3a16b2f911ce63e0d92366317babe1697b4e27c1524bd2e7f4f2ed09b986140c97640287ef9fc016d1b57f7db61b105f9233ba8fce40e5a626c6d8a82b9211e9b10dc450668955ba78726d6479eda20265dc291e91a074286b332bc81e78f836b150795fefdddeaa8a70df5ebdd0fa77d8b2e20ec85d59cdb4a36effd0272112c3b4b9795ef085414c1574575501689aed65b345d23dcf186ba11fa2b73d3f37d8c2d57c83ab559f086db2826c88f283d6;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h1b3451b9fd5a9cd81ddb1bc50b675760bb784e1acf9c2541dd32d6429caa75317202e502c56cac38bfaefff77338d4e872605680fefb5794a378144aaf4d5f8ea46755d2c6369aa7fabd328fa57f1f4004fada2f413509b9d09eb52747e7ef783fc08ff36876cc163fdc4bc46f369b1e73c553b3dd97cbbc444eb882ee43f8182864e401ae6bb97013dc662cc8505957627fc8b27afdf5d0040a4ef3b71a38b0d0a54962b269d89511ed4028b39ef1414e66876145b8cd990ddc611a60038f166b8055f2cd057aef91a954ab58a691b6f389be504bf43697e206abf13b8cac1917676c9e15a483c47bd567b133501f0b42ee1d7ddc7213025d3eb39c473ce0ec9e05d27a98ed457a0e6082442aeb244accf4379f2a9c65a0e984f6c7d1e4ee5398d6f36718ed9a97c2ede1fcfbeeba9802debbe3d208424730ea49910d5aae5d9fd81fa2;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h55447b92e2bf8fcaf127b41f184bc837886c248bcefe54c996d9e74df4a06f6e6771a235735971e66f8ef179d5b4f4c631e7339b35611f8f216f3f780e41599d89083abc6b1cfae43e9bdb3ee24b2831175ad8fb3d98866dc393e76cdc77c79de7b4f1fe9f2cbe54cb67b5551ed1de42366b0d7871d6d4ec092e4a686ebb7b5514152c7bcda1ed3e67ba9c377099f663a6266801e7524fe0eda172b70f2fb65c86c57ba20917bf591351ae897cebe2067d4baa5f207b818509e9079e2d522a12b6350bfe77af21ecdc5e4340c876d4a5fd3769ee9c019e9cf936e2e76cde72f78687ca2ca469b20502f6459c5106be9b5293ac0a1e11d6de26adae04c1cb8947a82974d1b05ac9456b6ab5c204e011930573fe8b4d4149d4c5c0d859fc0261ffe50b98b9c23344815d0c6645847e3d4dae8f6f8af828114c27f9499f295018b8b5d59e44;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h5e6f5b641e1bb403d280354504f1d6309d5d9cd6f2da80d8bf615bf4749872e16033d61d466057e3f0707d68c0ceac12aaa2842236d01c1757644daf958ec0961a1be33947c3f564cd7fdfc825a663c07bf46f21eea2c816bbb1501cc304362e603540ebeddac9f010ce3d93aa58e565b76185d2ea57d1941665c60aa5a4011e115d1f1ea2745a7d6bd224a805ddd9e65b77763eb220bc5525b4c8a9072e033997ae57a66f6405e5aab530230047d2434f936512404c660750a453a78161721a7c872b594ab6b2f188cf11c3cb4b63dc21329ec7531a54920b04a4811ab43b2ea5c05c42b767dbe4e6036b1ec52218eff8e460858fc80d3aea7cd418ee4a046ba7e0a52c9ecf02041329c1b51b64634d4d8b432cdcf1bddd3c755f7f79f4654dc15daf5423082bb312c7f734d1ac72778b9e4f6f2eca9c972f070e9846d50cbcc3090fc3;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h6ba3e846af0c0f37045122ac4626ec6696419ff85724503fa9fc182a6d925b2c2527386fdeac450ae95a9041a3dc79589ec7a36bf0c5171048a340150251a3f069abc683af2c212421a58fa7f046780309b2e34a83a6e76c31c3a7c05364f9293f045aa89ece7c2b14a72d9e94b1966f9a64618bb8947be3537c3678290c3c8bff07ca02a4a1969ee6edcbdec9d3658929ea5fbda2bf997ef208f4c976a2323a7c0f70f3002c9135411424f182966892ab12979a28949672abcd28b4d553ff29d78c54c0d7d4ce94b4b1afdbfec352bace4b902be44db93a81a1af8f237a1b584875b171450e4377ef876b24db954b89b5e2a826dba07b32616a05d54a9aee9a008aead866efcbcf65cb8dac3eee0a926a1224e5c8037b0d33274c26b0a6e36a5fdf0f73a629c168071195a9f74139945ec883e59525e728055b2872e16bf0242489bd05;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h51c21ae5b2bd512c7109b05501ed8d3561b68460a067fc730640e6d8c14550fb23b4009577b4d499cdc5da1858ee084cbd8ea65b58beaaafc8d9d440a9a9e142dbcc3efa8a2b7eb14428b0768b757113f2779c7962b17f47e80a511b098a3790e75b279efdfcb24ed528124010e1890d1c6d02ed99024ba25ab53dbe6dbec801f7690af0a5eb07b6c0fae58c111063620a53d5d5c6e2dc4d6b8e87d0289c4afccda41853ad7249eda157cd82ed570ebd7baa54b6ebe8225699ff5519d77d73d67bf47a9217ac68dd53caf4d9969665b56a16d6aa7096fef8df781eb5d09854450f416c0dae2c8a8e75fd54488b0c5e5707334b59ff0dd26cd58dd854c132563242e5e769cba0066ad98495d61b82c27cf54b0d263f51fd7269c11240f21604ff64520e7b94144d20cee1d5fc6472fac7cc63c2764bac360950369b587e0b49485f2cb708;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h6484cb604a5782756989b4af9b25264e475f1be97df78e30df2ff97f743991b973d9ec522cb386ea09b8ec44abc4ed86322c8f4c7ccb14f849078a70accec5029fa60c59e6382052af2e8e05a4b35cb787805d7b9811489a19dd5b0d01d67852f057b3824fbdace3751e45751ce3ee61d16121312be498b1bee3354bdff16c664daa4f63d24d9742442e7a8830d44780cc764b10c29efe1be311ed1d8d7d643d3b06cb54417ccedb37784ab80d8d5b6a9a3d4b7d6d4b7c8ae74ce6ae04b6cc1d59ccb5934521674de053eb39c597184e873f8fc16bf582110dae6a65d3825a1ed83d5bb68421796982057c10e8d10a5f9461f1df9ea11e3f9ccb49e876e8a841be181fa50e41963f29ce4fda11e40749c0390e263feec99583e81583324285e0b50ac1127cd0a929279ecf24e56f45c245888336eb46636fdbefc6727012ba5c6659f3c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hb06a3886f603b56928535812c9f749b61701d43de55ac86159ac73a44879e48669f843efedabdf7fdc9055a827eb3441f82a65ee8b4739e38d793a56d9439bbc5bc832fe4f76aef48c7137d8a6ac8d15b9a90ae28354455f4f8c795ba4ff390f2460937d919fba2c9db45d6e5ee440dc92747e8356316495c57f1f5ed8580af642eaecff80856fa760d1e8b8bf586a8aec56c8faf64327ae5722f649bcd2d0f2e04fb40d56e28201c94836f309d1702ad198fcfedab8e5fd3a6c920269226c51880b57bcc4a52e0a6a5eef1f7087ce288d4e4ecc92c4ea4a42b8a34033b1b8b82f27ca43f6791699c973ab048fb7eedd13f88558bfab854b04172d1f47cc44c5c28e2b75182cfd3e696ca4a068d785a1146947f3dd08353319652d96a4413ec78c430df80ec52aaccc4c40c1d425556804534f041d63b4411425440ef1cdad1c4a3bb91a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hfa86e7e225465a823a457cc31ef9092c95e7a60507fa3c7c6dfd90a9ad5ac3a68c3dee68047f0f6149698985f50f39c19d13ca5b5586960f1ce967f54431c2cdcbacf2925ee40ed53ea9ef5f4855ce7e7de51d245fa54ce7400f3c1f226e5962efde2af6beb54d3e60cd2f2cf905c1c71e53f520c9151a4e3819dd7618ccacffa1ea87396514b0568a5ff7e1d0d58a37c14e1ef9d8dae096f92dfe30bfd9ea8761c285936baa69b357d37937368060cd2a6d73c769e2944eb417dda5f46edb36d45be139fb9982361eea6a07d754e6eae6e3627d9325156094c59b8c4d40b1bc87de50c3a3ec99dbfd3a5d046a77e98a8fe0db693cd86acaca1d6f8474ca736a345b7fb3d3fd9ab959e0761867b8d98b29e5bbc1d97fec13c648c1ad08763d1e9c7aaad61cb898f1d1d95a2bc8af12cc49ae727e9c0e893dd4c63c608be2f34e264d4152;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h4ca9319d2460fb63281d0583d34d073739d30eb25e3183f4a26ddc67737ef4e1b959eccad6974e020f278f261108ba0c4f359a5c2adefba898594a4e3cf5d5cbd1d6cfb8dc257315f2faa63700f933d2a281658fbb39c57fed4e57f906caa844770c20056d8a58921147b4a2d8e11042468ef98fe7be86f15da1d36c5a806bde301ac392ceab7bb0fef1c75a9bd4349e21a417a1bfe37805520bf2914bf0aba374582b2bd00dbfa679930fd92aefa2496eae37e0c64e41e5277165fbb976768bbfc1d660f26aa7dc790a3b26e615a4aeaf001f1d49325b31c721a7ba441282596bb6ca55cda77488d522898e0b1810d8f7001571f8c14f865127ebfb7510acd1c5efbf0bd3c74511877ba9624e10165b5226c5393e0c04fb92a45b5165c1a7739c95487058f6e1136ef5fff4d7e32f8c693e382e68314d0275e7c8c59bbb448050f79b9f;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h3fd4cfff10562e65cb22b8863f0020775966b212089c0aa31fe4000d33d71e648ec6f839fe54ae4fd311b051eb6821c4e4e57380590fed0d2d428bd184b8a7974add2c89f3ca6828757099c451b421e43b851d1bfcb8873253111e58cbcc79dbdeedbf84144f0abf7d243426ec8ac5eb8ce1932eca29272d5475c522d3233bf22ce81040aa4f69516e9388b261996189510e0b03354b23d445346ffca23ca0db5034cf3d940ce9802e58882d4d1553629897035b0e3f77a7c5bff4388a54618c2a8dd21f60835ca79bd6c0f787736771fb28b328989d866c855b6d8de692ebb30cdb19937d6300ce90818b98b1ab62f2e0983c6d12561fcf98b08932f6390bb1cfe6166fa1d7e1235b7e42839d55f30ca2de0f10fd15250e205f227a5318c3c6737c53b1e71ab2c0d062080a78bac896ca014acf9160c60ecaafb3df8010093d7c2b02ba;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hca9dc440e53577484058bec1b36d6d53748ea7c6a242924fbd72e6bf7f2daeff96d0cb8edbade643d1c41fb7fe6d0cd502a8390f2d60e6cfa72f6ef7f7d83baa461b7b53aba3646e73353f236523619978baf452b1f27e5ccb92b734fd0abc900c697060a83bce792377d3b8a7de428f218a893556b33f40f27efda157060fd4511ba7653a660d533b6bfc6222818d1b02f9a7efd29a42be6d89c304b0a207b2bfc7d3acb52509afd01a309e8906213f9493752ff763e835bd126460d923672cb682fd0fd3aac97384a31e91184978e1d2129972eee79efb2da9497ce9aa5bc00c1248f1c7bd73c0a10104e796aaa796b44db6bcdad57823adbc3946b72f87de7117bcaf8a11b50a4b5ed9160bf17579fd901abf46c1e7149acc80642b9a069cde33460376ff93a14f93164de6e220bb71cb4153bbb3adcc384f6073eff8e93d688f0075;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h6b69759eac6b8fdf1e00ed7165efff7690de8dfc21d23b8928963352487ebf96c9226ade1708986a683c5737147f66f126f702b246ad05bb9ac313cf389f7544aa68f7abe49e9c225bc53f86d24f98e4ca59f0d726fb47d7bbd20a21e76ae7ac8a760e9e0aae4836f45272bccb714a5c09592e40d6d5a52a2dffa1167c6fe568e1d2f653b2db0afac69613ca87b70dfe6151b98fd311525f4e9f4361dbbca6923aff57f0777636e8890c04cdfb28d618271d6bfd8a295c0547490430063691cdb1fc376bc4302ba27ef9943f77416b3a001024692316d68d8a064c6a82af16ea7349c64b7073b0ab6d844757175a7edff7736aea1acfde0a02112d6085c9016275a0fcb2928f09e7485d398b98a8243ca61e1a15d12f72ca0f806505a78a22a93227648f26bf18facb443c5baa75c18d7914ef96b181dd9d29173cf27aa8941d6caca1b0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h9fa51bd431f30b8f185ed3bbe47b3f24f150294bf5335021d2de3fd5f9ed8a39d1e2308166ee2f654ff630255112a980865a31166c97388b172e2b25d5d8293f002a3b004b2f0c0cb33e712b35c8931fb178a9a83e692e5a14228607da54c9464f594c26c0b158be76e6c45be77dbb938f4060e6133e12a7b6469de839ef13f3dce35148bf6ea2bd6df491f4a0e065b1db59f9b585a6c8ae2480b300a378aed0fc08793e9fc4566001abc737b0fa2d43d7e99107d7c87f1d1d4d22ffd2725922f5a3fd8c167bba6850b4c4bd5b5bdf1f803be85db2f9b33ac39551128991b573f0a5e2cb9f9d7d4be057334071f7c267e0378b96d771a0597c025e397630faa436b2145f17811e0de2f437b8f80db79370549c8f3172d133c935102f19c6468527c8eedc233d9e773bafa3580c6fb9d22d282df3a54453fd8db925a8b2426b56a51a70fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hb2eed7b0aab678ec05f1bcc42459093de41be96859a84149c05104dc40f5a34a54adae6fda8abe6f21fc9248279e6905ca6a5d086b75af3d63c97fd4f5e0e086aa01adb6dea7520396f9539bdb69880fe6f4118d7474b41076ead13fa89341051fc7d3525bccede0f80003b3c6b29503544962bda44ae3f48873e94592c155a7e7b427add96a1f446957c956888187f15403c685d304544186df26c8ae6f8cf8194fd50bc5a78acf3a924a6d4485a50dd9460b44043cdde8cf5353632ac352489edd0e882c9228786a16b540fc931c39a10c0db322719e9d61a90d37364eea0f4005d76f08e03a3e4f9a361230c4ab3125b7bc1b1ca0f5fc92f078ab4725c64bfbc3f150ded9d07c1acaa6bb63b961883238c9a1e93b5b530dac36d1dc751ac456d65505d32d4c113a61a07cc95a4e6ed930d50d1badb373f2440d03da6f64b4ac51a9fb;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h63e2240d4f020a1b48412323ed9763e122cca0550f7fcf87f86d33aa52dd1c95e89d194fad4fc113105ad4e981f82289c8d565a9f892e6d708f4e9be719d480db94d9de5d039423ce2f803675db4a40a442bab1ca37d844cb9cf03c925bd62479fc29bd7e32129237aab38fda2a1a1b612b48391c10c8e21790cdb5bcdf9c1263b720438af1799b0808479952617d44d01b8fe5ba32ec4cc15f44d2c34434f98c8296a55998b6123e77be757ad967e6b32c1ffcc5ded9b5858ff893c077ae0c46d9408bfed36a79205e8bbfca51c0233182b6b9a8eff6661e8fd1b670a8b065ddf8b2217eb75ef9e858e2fdc8df074b09c670c7c05c86e70165dcbace9087dbdf240c009e4c71e571b661ea32107d81f83c9aef1fb5491a18180ca5e8b4de80059e975d8e4a46e80ab03e40cbbc9358e76ab7ab614da2886699a348ec65bc89769b2434b;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h369a625438e6e65034a63de66b5632e66de5e0803af23582a069de718b255d3c6f21d72cba63cb622e50952049976000eb50683df19514a8cbdcd30edbbbd17b267e8c750a47f6eda83fcb3b36ff928e7917a39334787a1259ed9bfb45ce184909163224f608f5fc9a0388d6600770abf3bd9830c9d773f6bff17057333834b4d9d184f7d416523cca2cbf7b39dda6579ab4fc05b46f66ff40abed4debea0fab4328871e9c30757e548e22f79630afa8661ad718e7841af294cbb942a6142d8f63fb9115ac5d3431926a39a38097e0b62b385361a0bda39bf7b8ba2941700a8fdfc98425417094ad1c813ebe3edd3663b968545e2023fea646fbbbcb152febbd29918f4fff6bf3177c1f825f35f331b97875085e80c6e23d0104b298d8167c236f97946eaf65092e68b0eec390e8e4a1c4280652cb570641879dac7286af24fc9ea36f86;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h97d525afc518c60e2de717f606e637b0bb494aa5c9d8f3e67cca6e484650ba78f1c4f16302e10177aa683e4255e43e4ac11d86079c123da8e32df89020dd62d30104205175330e7a654935079a9b7bdcb163ce8b568e88baf2aee53139712cf4ac90738eb9630e55eece94f869e12012212742224e27a249bd87148dee422c2a3f85583945d638802fff20437007fe7e49334ee5c5c321f352fc1d96de0f2031a37ffba82d07df2a4c9f9a72770098335ab0036afc47174730a5c673949faea237ff8a4a0a9cd317081c356158ac36fa7aadb3b825589cbe404358bfb252913e1ba490dd6007d2bed6fdccee7ed10f30e0a031cdfb4c2e5967411a4e321a86bdc6a9cff2578c43fab26e799eb4b02d865a118f0adafa83059aa22332528ab37242723059ef3cd4ed5b70b85c4f38923d2f1b5c2132229b958c07b82fb8a33cfed17b87c5;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h4b699677b352fab0a6f4ad5aa7409c48cd687fdff519e4a9181bc3fc2514dfdb07f46ac674c9a969dc23ef42d353fda642bce3e41f979399378daeaed0c40d91a883bc80b6779af36bf5775b8e44e23eb8a079fb906c3407a2de5f2bcf7acd49e89cd9a41feeb094186161ec1caeb7b7232a88bb6cc61bf5425d4deb48f8aa010a5e544b559c734a6b56c1c635239b1ab6033068c756350f73764564ee8ba96f6cc8d029f98ab36c4ccfb9a9f8f24769c89bf37dbf86b08364198324d1f7610c70b58a2c80314f59ba8dc6fac4cd7f6ad99e56655ec71ca95a8b2c7fe5f1440eae74e30d9c1f5fb48c3b964f93b679af1749200233a75404fbfa39f98bf7e0137ca9bbf51d1966cac9e1a762efb500f36d72be78c04eb707536c39c080a1c5a6b1a9e5ad8db0e02e90fe1b3d61c6d1ac7e46934b8e9f893994b0ed54dfba06ed080a5b8;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h8aefe43d8f85527f4489c7fe2e4962c897fe8de7b33a26e4bb70ab9f3e812090b70fb7b2fa65a91ce853668b1e10c251e476ddcc399d03c4368888d7a497243b2ecc07584d63df61fe056427b327c03b0b9477d3e09a67dc272e14bebf9280534e18b069dc2d1f5a1595b4b8e665b87c3f729e036b1ffa46d5c47a9db0782c4f6ff06acff025a4cf326ddf106383ef5f466cae248b258087289eb750b50313ee77eb72450db1601096a21af53edd170689a633c9359bec9b972c3661668394ffb79e15c4c0273c6b216d7d2bd4dc5adf059c3f81b4e4e24c1ee3666a1286ea27dfb31ed220e6f78f3abfa67a3edbb177b2ae39ee47f36d4751f96aceca0b148894ee551c5d1aa658de45e5ca1869f61827633d90476ea99b26fd1fd314508013a39db38d0ed1e037e6003443b90fb3321fa57bc8763f21be42e9435921ce9d50be06be72;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hf8d2a00930f62de59646430061e69976c8b2c147b74a19a3e1d2e9ac8608a6315e2982a39d255a9a5b1d12507ca0f8daf553625789b9479070b9007cd06c63802cd54f037bbec0923a21ee293cfe74d453ba4452b10ff95cb3bc659c637daa8cceff789c37f8db758d7b23c37c0fa4709212724bdc8b16c2dce7b9b0174a45ca31e192fb500cee40227ab78e033671a08747a5f4ebcbccaa448a8ea1585d352f3062d1dc2a60b0223bfb376f857d0043ca965a8aea0b097222d18df06567682f1de0f26a3687f87c8dc52004fda3067203ca15fa3f4994282ca83e3bfe5bcceed1d68519ada2e8b0e6d57d66342c7b0877bed346fb861e0f3ac45be46b3784a152507a6aa533e03eb7e0985359b6f2e2f7a65aa9f47b8ea19d1aeae97e375cbe6460672d1429fbd79d4ebcc71369a728a2bf4a6a06c18ba5f3e78caf3428f0e5ad377e04;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hbb3420c79cf3e199cc46f5bb0ca9be886429011ab8d666a32c55599f397b4a9bb8b0ce96e4fd65fa8644e2aaa143911a0f7b62086092fa762a34ec795976967958cf8b72227ae13003fb55afe9ea7de5f9340a0cf3f85639aa087c107483b1fbe4df1dbfdd00e6fb43f15cf4f8a22042d0dce34748bb4d2ecf81dd5c9ff7107413d383c6bd3afb98c4ac1b512323041988db0c53753f6b25b5226d17cd6e1bde43ce3fdc2be14a450021994b42970218e2b8dc71381e6e2d6bcbec91f574a27b784d767abcad1500d8e96973f0f5334a00fb4f06ae1f462aee0a5129b134c9319540e0588b38e8ed104319b42bdb7fc607108192d5f0651b4031bddb30b53c2bcb5a72fea7ea3f5e50fd681d803659888c7d8d457f8aa2f744fe84d3a2747fa92852ef8f4b64123aa1b34e8cd8afc486b6d400b3b09e759df32ce18e6b745c870706317;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h85719203d82bf0a05edd94b6f0eed2a693c91725fdf9e0d64aeafd1ef6350045c3b97a93adf2cd6280b9e39b0911c6e46182bd172ea82d10ff212833f5bfd3931a7a9750d01f6b1d8bfccd08ef97a9ddbf6e9329a5e51701832f365fee57102418b530a9436bf968fa8dac3a7ecd56cc0e4c4806783a2d302eb462fedb8705cdd8fa2a438b6f0ff4c34e241fb4dddf99631985adacf4180a2a5e9f4589de8bef478c5f4badbc1c446dab8196d4589cb9d0b1acada42cf82429cb13982c102f165268eda633d9355e7cdee80e2a90a313a4433b7be851229526405268657fd93a07acf574218343d68ab63a08d77873af21704eef4c725191415b5af06534b56ad9e67c07f9ba30e449b30161be7b522fa3bab220a3c9f26b86a7655fee180808b527c42d67b10c6713ea95e0977aeea386f6e362647861ddda24b49727c5dbdc81cea39d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hedd695e49ff2edcd930cb981f027618225bf6803fa1d69f558944ae8fab08de8b16458fca5427ea889eff737dbffa06a705cfbf83bb8b07160fa987854c7d28065eabf1a08c636f8e13fe996a7891a984ed0f138d674e00806a87204d3bd13ef4631cfa57fef6c2a5fd08c7e67557ecf1b168091866a74538693aff488b5356a10e79a36d062e966a810b3b60e20b4d27a87cbe8eb56a5bfe3dce46e7b4c148e8fd09e551313af2506d63033add21fc8e20977aa5fc457b0e30d83ddc63c770efe91618b174644c1a4bf6d823995f7b453cf4420c363b2957ac23450010f3307be35221cf9be6dcc52ad49e2f5098b12c21c50cd9388b95e48c935f50cfc3757589a5542016331fec43724bb7ece0f1eee79ae81a233eb55e1956a72b35882ce61530c33dca7d3d87a5d881fde03f9b2fbb733cff6ba2ce7766dad12b1d617752e411d71;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h35150c06c86984b43a1615fb0da621d2799106c6442e3776d6b285c65c181a6fd2dfd6cb3dc2c7d98855f7e4e1b6fb2daaab218dc03ac48416773de86bef2dd0dcaa1ec44c429230c83d72c9d770c420e8e7bc28e0e4e204ce764d5525842871bfb21cd6a869f5bf8a81231ce2bcda5a52c3f110a87cdb2bfce88bfe509be7f0499be37857d41c5f4c141587af063806afe07adde7cc8a4ef37cbaea8e6738fa6dc1dd588461eb2fdf22202ad1fc52dd3410e15edd780a4e5e7d60afdb9dc2a99f8a2b66170218ec2bd9fd8a005e07f53cd3338efd42c51c2e01aa1ab2bf781aa132fbdbc839c2c27f4c35b5dd5161436dc3681ccba1ade435a71ed3234ef2d03e4bdcd2e3e1df5999ea8d4accf7838ad0761cff27efe170f3a6545eb33d4158983cb9d43637a63c17d544d9894142d543d487dcdfde83f4db0506a3b964ec42ba5da109;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'he95c9192bc87d252e5479df2a2f8bef849a5896e98098c03f1205acd8026f518cbde9a826fe6eade2e4da5e5c08de95209bae60e6e9314c2a56d0cf37f40ac77564ae02f501e438f10113b280ce49fd4f54b573ca27c59f41221a7da8b61fec0b3c8a3ba83112ff471365ff223fbb6bebe7590b1b89e530fccdb146d00ec512ec4f1e32f4d7a9e478c4ce5ef6c589d29f31a8140aef6d16c6a90120088980884339e1d4072e1b54b552c2b20305706e53f2d5e7c4c72d5da0ba9c8f66678d8359b792ad70f08f8f994c253bf0f6cb3f2d0c7e943fcb42f901c370623c4ccdf17034ff52fbc3bbb8814b543758e5ce12ae290f73fdd2dc18ede5a27b2bab5381915b1c2e4c88c73ca9c211e385da09beffd62bba41fd29288dde2a98f946f94597ac27a20dfc9d3ec35d17f614b153a19923090443202f6d7e76ebcbba57d3cfd86e502b7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hb3fe16e47f862e120a0e83d02fb4a72d555eb3443fc39d8ebda14708a50a51ddecb6a86bf45d01e88882fbb1f5fcd5112925adcfc8782b19c55eaf9d7baa3f40f7b1ebc2ee183379d3733267aca8754aee38da09231b24349e8bd824b3cf666388b35f6b9ca267245c69d01c0570972979d8efff01833491c89f94fa8b90399d119bea1e43e0c678caf69cbe1e8dcea7610f9644097357803c78c8d90f6a81e4e7071bb8b2417bf51d35b9fd74f8d407b26888f6c767ea5e625675f8d184abc2a72ac5b8c277c62ea231260035e324d3af16398e3cec4aa01d312c5dbf612de6ef26ec181e4a109a2f9b4b0f9f3c651c878479a3412de196b97df633462961a9c86c296d64243841e909b418ca70ea4de8a5007033e0376bdf51135271346920fbb964b4f26a5179f4c8d062fce7f8d009da84dffe2a710059491f2b259f08500d0452e0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h9089e5c01e82b7c0a26f74326185ffdb3270242b68e1d85856e6e6884cfa2079ae133ff8afe5af474ecab179079ecc120134e47ab548bc91d4c3acc74d9d62ac49d7e211267d6a2c4a9988ec291d0ecd8202685fba5fd3b6a772ec96e1d51081f7ce79ca8c1eaec68446cad0ee5088b9c7b46d6727ecaac062ec9c4ae8259810ba400dca52a09d6fe802973b8a1476f8b5fe08f98107060f7e85d1d1172aa43fae54b41a2dfa3052ecfa44e0558136b2fb062ee85b9daf6ad14c6087fe8157b145cea62568370431a5a246393358f4fe7c155700edba4a22a9a42f6a5fafd16eb17b0f178364477668747dafd8d4ea9edc5792d02635576c258f578c9a393750c930241c05d42d5ee48bd297b26f1bf4cb2f19278f34e337e64bfde02e3ce894ab5adfee7edb11ccc2dd788f6d051ec33a5c870691787b4f90b4328ee218d6210561e114;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h9157c20b173a7e135134a5e51b16bc31274725252dd267774e8651bbd626ee880d6328c81bb7f582a8b5fba1346356372d954b4808925135fcb95ab3d33ea4368a50ddeae77a3bc61c27c7b8d196fa74bd8b65850708b887021832383d5677a397a37bf73da8893f53825c223d5694d75b9203e39e9e514a41262f5e6d0b56abf8d05034f93bf38c8f629e636cca06744f66206af13dd342acf2826577d6161d7c6a3b4a619f01badac22bdc9e6a34320c4f585cea8102d8787c07ace9db4f15e0e3761850552cb177c4d9e5cb906030b5683ee7f497c3607a352d4ab3a527f04ba594b54b421243bdb695b2d022ee7d1128716b1b1bee5c30ea6aee8410830956fbe113034956311742a94cc474fd36e003c19e9b4567f0bdaa11f4c9e64a3ee2c2980c37d330753ff5553a47b4bf7fc3161093d41a4f3279de4cc427f21cf86103ca9d;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h518d24b158bd91752e962637fd4af45ab86e8e16f6c0a52a83a7c6d2cde621ec926440f1892f8e44193eb505d21a5bbe7ad8ebeb95ae352973c0ee4cf4d4036f968d5e7ed258ffd3c5576f3c84d7196f52a7504ce9d48a0e6ef3da443fb7e93eb1e3a2c9c182ff8e6ef44cb1ffc1085859f2e803e6001bfa1d408f6803da93c7f32b2f96fb81eebe2c80f3759ed5d99ba1acd0ae76db070214c70a3f700fa9a570712b10e5fa041e4696e277d95a8822adcbaaede8c9640985c8b252c41998874f309909dab556bea41ed9f742728b36e8cadba377db4b2435b997a316330c760e34112b5b6253711cc40ceabdcc11fb17027181640d6b758b3472cdeac401a19d44d96c6d763eddee19b5a8dbc1ff2981946312ba06087a6ea8f29e5aab1d277d45384fb4df5137a6e4aa281de39d0c2e76cb9846e9445b97cc75c89c91308cc04816a7;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h337fbdaa9a8972d3437f8a91b17c777d73ee9403316ea2c207b0408a7f03f21d82c725f58f6c97cfacb065ea39ac4d07e9cd785b81dfa16679bb715f40787862e1838d484c28e8ebf1c85d0e667b80be99e19f52b002cf135e5ef00b84821b9c35dc43b2d86be84ae093424ba9f4bec0d3598f5298353878c5a58817ec317e6fdfc98f4371f45cc8fc5b5d38860b5b8a794d01d6319568058f8316c6933a2e9cc11ef7f617550e1cb52539ab920a196cf0cb8bc7a70c8d52ae1c3f897ca97e1e11b981d61b885482431d80f7a93800e4e186f05dacad71d8650891134560f8c6ccfb88bb9ce7db7d50f9b944b288306553d461120d2b84f6d9fec50432223ca55e9676ff6344bc6ddbd4fa8ae90e82ebbc374f8a403d95c92aec99b81be37b1f35e9d307717a11c48a653412625b38f2fadc25f5cb573fee45909199ad9d7c97e6ac3a96;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h3d1f228ffd31e6137161eeab0a8c25be2fa801ec3327574aff4e3c10b0aad7fe8795fd17584d77a84ef48204965b9bad0d0d933fa2ff9e1ff3d1b5ad5c4bd801a8dcd94ceb035d9bf280b7b4a0f2af8801b4a4271d31fa7ada2295638f9959ed1c3f361f21e510b7b92514130df0dad3cf15d13dfc71485be3256f005132428d24ded4719305c05e39482a478b6df496542a15453052075dcb6160faf97daa94f71350fbb203b704e033c1048c81a9f948c216c0a54755588706c0ef60bcca1d8094441eed5dbb561504fa293a0a1a97458d706ade7d4a9891ec852ea29419cf0ac3d8f575290ed8efd1df65ea38a10e5f4c23d238a962ec00673beef4db998cc78c2a37f13332c15cf84233b57b483c8d376d5e17c84cc043218b658e7a15db05fb58e01d4d95e6ce45bac2eb3ef3101e60c741cbf0d82d63bd3b11f8b8d843a7dc9184;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h217f461f4024bbc08ca72d178c0fd4a2542806963276c3cf04559597f6ca4e8fa88280e353d446c3d2327f09216b4246286e1a42883ff63375210e9fb224bf48af681f94b1cbbe0e15a0d9f2a9b03ba52ebfe003370997033568b82d604b08a1dbdcf842751a44409828a28beb84f63bee36190b532a5ff24223f304d665c8b05e77959b789bf387a43685c7cd51837c245b9c44e78891b6d829903bf06e49b9800d3dfa58ee36e4824bd1db8671a2f565aebf9a4b835a53dceaca7386bd70497c9c68fc3e47ff36836448ad53abbb0f74d03c54643d19ea065c360c2103195ec46bc3a2d6db1c48a591598cad5f4897ad7d8515bbce4f79c8a660bae39217ef7d64d2ae4030501958ed3b00e9b9d802469108cf7d132ac977b035afa6925cd7006f559e13ace7594d275dddd659c670f3d7e86dc3a9e95026761aa2c3bcb88c8bdb173a;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'hef9bea62da0310103f2aa0c585692b90fc2345a1694f3d77f05e23033f219d8266cf4db1ad79e90d0225075ce61cb33a259e4eb233b7f41f9f7216ef8c0fb448a254816e93b8dcfb162423a68b81f4ee9e95d4f1cf30ff18df5fc6c223d9eac5dbad967ab8b175d6b294ee79d1e6215eb248626ebd9dd887241e527dd696d26e7c2f624cf0799b5b06e8b42228bd03a6e13676542a06db42fea91deab33aaebb7a1d32046833bebaeea90519dcb32ab48dc444feae0ce580adac286f971602e1ac83b30d18f11476d0e41ce5214c7623d36244891afd377691ad9242c039655511e25c1053950851eac62e3d8dac3cf7fe3fa1f7062f79fffa6714bcf013bb6472e1ad0228f71c8d306a00c81d319a2613e6b874f519c64c798ff32e2f039bd5c3251b73950cf72645d7a6a564034ca508932758953eddbfaa8c4395c0ea6fd3bd3cdbb0;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h55a4295de5b638a43c328c9c0fafa538c0f5621f8ab911503fad9a15a95b924a880eaa592a76b550151af26fdfd02ffac498245e92c6247af923b3211ac7907f2074f57b93b20d66e06dc437982445158c8bc5a1e51d7506bd2d873fe143823f098f15b04dbc75cb2800654632703113af1ee8145a5d8df8c6b812c71c2250bac8506c41107fb19ce94e1ca71ac524157ec5861fd52743bd394264bed9c3130df674b2f909cd0d4f433e75262769d657d72ad7649d5e3fa0e5037683fca7d612baa49c9b6cfcb1587cf0212323c266d65fb399dc29e3e0274e1d2f8fe466f9bffc9f5bf75a0c670ccd3cd4c1a2e6dff4d122bdef1959c62003a7f642fa08becbdb7281aa3808ad143263d33b0d4ce3f44a88328e5f43ad4c03fc90f9acd93d4f83ea43d5fc703e2b4f7dfe6fbf970173bc621f8a8eaa6d84addc27fb86a093cc937198c;
        #1
        {src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2592'h4e3673c9fc98caac42874893a177002ac936da4dbd6398b054fe56a3b462dd336cba96496f55a2a69fc11e238641e90ba4c6e03b1912e976d953446b532cbce9eacf4edac24250976aa476c3c51e2f27b9da3af92fa0d91fdf51f04f97f2d17d7c2384524642eed6859b19dcedd570d8abe3a494c7631e8f0ddeebc6137379b6669543f7c317ddf274e35bc41340916161ac914c5ff0c1e4c1ffd36919a33c6ab30ffba6a99043f4b7463ddaaa0d978bd25df4e7386622468348d2becf23d4c8405082dc5544a87f112a2510149283751ad93ae27c1119e9879e8b4e24197ee43dabce944194b759ed8385196cfe87abc48aac5596cd3de2aaf9e13c549c934d3efec21aaa575ed65774cc6f054987b2485e9608a41382e51c286b9f8112256383b45c7e5aec0420f792e64a78f4c38829543fd50479302ebdad6cb523dbca4d05f7bc91;
        #1
        $finish();
    end
endmodule
