module testbench();
    reg [17:0] src0;
    reg [17:0] src1;
    reg [17:0] src2;
    reg [17:0] src3;
    reg [17:0] src4;
    reg [17:0] src5;
    reg [17:0] src6;
    reg [17:0] src7;
    reg [17:0] src8;
    reg [17:0] src9;
    reg [17:0] src10;
    reg [17:0] src11;
    reg [17:0] src12;
    reg [17:0] src13;
    reg [17:0] src14;
    reg [17:0] src15;
    reg [17:0] src16;
    reg [17:0] src17;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [22:0] srcsum;
    wire [22:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2cc44c612061db151b65e52da7fcb7ac4b9a640c5d3aa44a96c4c1cd2e800a525d574eaf391fe6e92;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b7c533a1a87436d31443b0a44cbbbf3b4dc1460992aa7cd26ce9a3fbc329024e6f10cf1c6d88dfbf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8643493b843dabb507649b63b499579e0456291fbe33b9caf2ed4b0c8bc983e6bc0439f73a02f54dc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9494ff06508122044e442ec8ba9f27ddb640217cb36f7671101f7c476054392d203cfbdcdd5e1a2d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5487bf1a667314e5062d248adc5bc338014f606a80c644d3607b305d7aa240136f91095c6226abce6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdcee6a61d50e04a51af3c16cd29365b5dd638298ffc540db4332776709da2d134a32cbea3afb7678a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcd5f12037a36f55dd697221f9ec1937054fe29a560a04beb399c4c4b2f10470a028edfcfcdb3d1d29;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd79e0e44ad07ed95a4373854d2c2d4fe62ffb4fa63676a2c16baa4d2bb890902c9d068b9656e7279;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1e093a23630afb78786fa56fe6bff2a13b528a4516b8670f3258a2a4f355ac46e107df2eef60f1b1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39551e83d3f400b03517b4e7ce65290b2b94692c088bbcd589deddc7e113331df9b0e68783a4a08c3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1107ed2047f27dfb2e36ad5c021e8ed479e9e6e87cce24a29d953e3ff1fdcc14f28eb661737b8d9e9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h95af17f45e367c0480d6b463ca6c2a2261e5117aa721e0f385c039c34f3a3ce169dfeecfd77402b4c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0838fbae990ab71475993a7444e1763dc44aab639e9b5e872e6fe5a90f5a714cd5da17abec8edba3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63536acc59c616ceba35ac07efb250b9d83aa849b31e4dd7bd52f947cb3dacd8388c5cd6f3e22fed7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h62703aad770194245892740f9bcdf9a8e0be4e2e5e629d1f6c5e7f3e01fc8e542887f980beb247943;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc13fb88e335aa03edef014aae0e9a34c539eeebf6f98764703c1140f6901368fd37fc6ced7d019e41;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6ffd82bfab14eb52797c9bc6287729c61652147c34d3867ba1ece75468cc42f53f47b30805ffc67;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha9e9a357d421e8a9c6abbcf237ff05f9b8887b9823dbf6e26c8fe9896d8083e3a88a8fcbd566ca0fa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h634c76c727258cea31372a56ef72f4cebadbbca4568f74ef906432c8461382988fba574bb82c3a7a4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3edbce6bd72c04e854ad88f30916686f5012f5ddabe20f187b1b550d741df45bde6c5332364bfaeb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd3686b3a50a13b3abe4a95d5de3d2df2463c298663c2687744b214984b58130b303300e5e689ff7fe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9cc414231db38ae9f26b8ae073a1318436887234426957f8886c53a190b602fd80341aadd172ac000;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb6102e57eaa9c326aadb569fa70cde785687c37066bcfbc56721a2a76cbc88b6560ae4ddcdc2085f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7cfa3a83a5e9335bd0b038cee315131f5aa9b3673a060e68823dfc99ff547f0b5b25099efd89bc79f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5349ade6ee9f1aab340a5544113ae4caae200a430711640c714dd92206234b40308f250a43f608e5b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d7a00fe0d3a207044ed7aad7e2592674577efd7c98b86eeae0c7441e57e071482d8871aecaeb085c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86ecdbd8d1f7eb6a9ed79f5c88362c6fd863683575589578bcdf4fa9923312c51fec45cc77a9908f2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha81f86feff2cf156c993ebc01043f062ecef3d7cd86b36f78ef938b094184c7ee3185a33dec04307e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d7818df388e74542dba2fbc1cce1cf605efe763205843a9aa31138efc561e92cc934e9565e3298ee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbba67f2259c5f3a70a2324be71e804896ee73f2b121944a1bfd131e37f39639a82372b99dc3d3357;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2f75cb7dfb66605884c471d0f84905c169d9ca432a4b356d6abf9955a181b2c0c1d6110c7467d95;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80ffcbacf04bfcd1a9d10f396a6b7a4815c8930ff1659528da5e8770d3fb3b9ec78f263fd78faf35c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59c0b34bbf992a84fc9478a8a9bb6f9bc2a5dcc6a9e297b396a2f1eaf1cd95e7631b710e62594bec6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h90703f0c6e81cb749d3f2c0a78c2000ca27f3f885bca1b45a62a096a42c1ca92eb5d4263b3a0409df;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf736e9e9cea5d9ec9b965f617e77d74af0beef95c78d22fd3f5036c800a0b37662ef435d6e64190d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha5a9db142054164dc224ecc0d24b84ea8011a984dba45c49c07930f700b624e378f29ac5e6704ee41;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9164977157c14b349bad1985f5c779fbbce07055b9495ae8425a6d8b5d8b54677f8e56338cd121eeb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b99636745ccb2447b4b159a950d5c989e86d03a589c023a06324b513a990356afba5174c1a9cf258;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76cb4e293df4b02692a2fb8131451aef02b5dfa7bf9576b1b31251c9a1d9ea5e4932525be17b42873;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f68edf680ac12f3012bfa6fb0fdddc2d3bc43abec4fea11d39f0c6a1c3f4fb02d509a2fa651c4e27;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h689e6aab8ae231462da84e52e1ec34de3cf65c4934a07ffdd66c580e2b1f5945c342ed08ff2cd3fd3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79920e3f118eb0c4659621c339b79fe503520777fa0380658d4ca8f607464f7280b8a4e14826f175b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc400d42a359d36f270d65ce8a599dd383fc9793e6ea8f40f349220868c6981f3c5ffad2423543e27b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ed117afa78d1c4bfb3b763e8ca2d3b2b4d4a9cedc0fa2355c83975ff22e1d08be9a466f14859e15a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8edc4779a7f62c57fddbee0e408c65fddabfcf3443904857371c0ecbf71b48263de1658d5ecd28ce9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5af27c058cf01fbdae9f344db338fa282a364166ce1b99a7475c6c397e5cbb27d66f9377148fb2b1a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdf9fcc10eab44f9951161970a61ccf8008b681a4499878975520c11b07d84c992c9b80204e3e3f7ea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a06af69310e826b8097e2f2abecf75861a78fe97bac7bd0dabaf8624c857380c82d7fa7785e0b0d8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h219daf565397ae9b3494ef7aa67bae8a7ea5485669f5613819446990a86460387d81bd7a39557b6fb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4bf99af94bb16b9664251809c043dae8dcbbd06322dfedfe0921b586f4b32dd403f2ef290d93f4d6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf47c1e0e3e9dd6317f313065daaa543c1712fffe7b745891552df59e6bbc6f802499c18b546a5398;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h963ec0652ce3e56189eef59e6d6508a4c9574a3eaea49f8d7c7fe1b2c7e16a66fc3ebefac1cebbf4e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h66d5dfe061964696629294a6f435c128d7729476d613dfadbff5aad02b9e58cc7e4b4ce5683525c86;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc321ad0f3ac0232e92b5c6333e3ea22ca8133cd1f840345a7f80cd23755724261bfd01f370f7a6158;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19f43a71df556cb01441b12a739d0fd09b6cc2b9fc52ff1e368367241201085506c0d1cff58893a9b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3147461a92cf0e776d8dfb8277d7bd45259d987320992a6b84230356edc2ff7d9ddb4dadcd0940da;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdf2992ebebce3882291b72b448602d6b0b1207eb01543ad4f500e717ac60d497213197410d810021f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf024a258563f4b08eb097742556ae418c855ac736ea899048019470ec301e59f3fe251df1657a4f6f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h985df407bd40d644ecdf757d52c95e4e768b70c9e0b03cd49de2070befc74fb4f6b9095f205902c1f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc0b91167cfa46032abc65067b7edb750c9bb2b876bacb59ece3192c5129f057fb097ea0174fe0e48;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf2c770cdce45d0a4208fdec05178cabf6663b204050a42013e806774db5276a1c8299a2764e869779;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb87f3f4b87331ae2c2f36b6c8fa1d436e8479589b0336c2fbda0759d5bed4ac1c2519a714497d8466;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82955d2456b591167a75a1ee590d2a65366643c9a568b9542cf7980aac0a60f1686de32c51c3ef0d3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h89d4f6015e192ea787a05e4132259bffcb1568ef37fd4d3256e4acbe8f6bd6cbb2e6c823a716bd40b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb22f98222277839ccf166e1d8be101af16ade821dc362440490556cf348a87210315f326afbd597e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f2129f47d47bb95df4abdc4baaa4d3c8968f87e91c47d37c48d4f60f2e630738c8064c28a7ed4bc5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfdd2b67b3712fe6ede1e3dafe445889b83e942f4f171b82176f0db79f409beb4afeb767de517c936b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h78b39f2d0baed010293051b07f1c3fc07c3edcc8109fb0405bb346e9e18a2fd48844625019c827717;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4f2475f0e2551533abae36c6b104bf1e7e1d79cbc4e57f1c2a7b902e2b6f5ddd8461715a0dd9cc2d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had0fde5fd9a6ca3c13a1a5e1241f2f9b8dff346f2544ca040087be837a9f630e11144f1d937cfdb78;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfd4d5f8bd886c4fc47fd8e5c97a2c69d66b9f521871ce4a310c317eba302d4ee08be3ac3c1209bafc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hffc3621150a3cdcbcbe1cc70e44b76fe02d0feefae2cd7abe64e22517d0620c504a52cdba6ba9430c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a3095ea3d70bf353a2f198c2425debd5b196e339011f5e8c49fad57ae8737144c786c637c932a266;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb7feda53802786f36f9dad0e0aa9e44127d987019aedccc0f7a2b4f42fa4223c0cf5a6b88f7fc23b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4a6dfd74ac64a9b72364c5a1813ae28f3c7548b95313d8f6e23810b56db621e22bbf0de74b8c048d8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1954df19d7f7ad1e10df433c2c310c7b8f1a538cdfbbb7b4c6169191d2a1a6fdf819e9883d0e7b7b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18f84852c3bf9414f968797a011f718df564c5d257596ac2d88eb80f9225f097f88f7b646cf95b94f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7367d80b92fbac474311322b81219076f130ea47ed7a3e564f86f85db58315833d6f09c5177b36dc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha0b2e6aa36939430809732813584755c042a96f6002f3d733665b6f373fae7cc083d20dc38e37e50c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h205502abf04864921cd469eb3de5ae11883437d660ddace547a00f12389d015d2bf9d6b09172f4dbc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9cc0534bebaeff89f5cf56da345195017eaaa9d116f4bba8ce67559809ed1547851b01c5c2e6328f9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8389949e78583caa260fa54cfda8015318b350da2587a9cea90f499eb6be2d3c419d9dc74af715c5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf708d59efcfcaf2b649fabc419b5992a01d32ac6d22dad7d276742d367a2168a1bb301c5f6678c066;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h659819ead498fdb469e18c5a5ecd0cc17ac62e2ff8dedf5c7e97509f281e953d91e679039694e510c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf348c6429b859df3d316f1ac295a98eb45d49ec3f080986d78db87cc4bfe0e3225cbd1846ebde40ba;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h596974b2279dd4a263f569eafcf90e80d6395addd4b7bd4dc35f43d347c33b1457de1ca13d418c5b0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h64c286640bfb5fc565df572c6175a44fbb0a00d0dd24c0fa0d747d091b493d9dc7aecb6c098d80c77;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3aefd615c5f4c554ef4c825db11880c69270080bf28137bb7075ff1b97a109b233b8f504eec2fb4b8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1ec5b2b7c32f177e3ab9717722c22488c49a1d0efba4680a30eb1d9f5835a449cd604d21227ec0b7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1a470bf640f6c2ef5ca5c6aa6366f47a2658a3d89eafaf2662552a81b645d6b15ff16f77627cd932a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbbb3e7fa42502b299f0c44acd673229f5c07887021798ba7777967036239aa2279652058c83633d0b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d286af302b34827e12eb817094d2d45cc1a7a7f6b31f3ff4556ece18d0aef089c0822edc5b450589;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h40f35d41737ed7579127b85cb72f2377ce898dbb208ade20e35bc959864962307939b7dc6d02fd69c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b45ceeacecfdd5bfc77a2225732795d341e4e55dc9c3d16afecb2f24b4ea8e460c2a23d4ce22afa6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1691969a517246dc7189440122bf65f8b9ec2f41b17bdf381689aab87c2283aeb33ffd5b4ca5d262;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84a7d5a2fa3a4b706c3d0268d2d6ed93af478e7b5f80bbce8c3b68e1fb712ec57c27d6a41f5f85bd0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hadff43217c159696505088215b71505e80c54aa18fb1e9f63793b520f5391948a7c9ae9ba4969db3c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9303bc7b909ebe9e25431982337c1f2b8dd5fefc14fd8cc68fe03480cc28e742f0a5c63748b289947;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h746bf2e3a6c5b9bf1b06acaef55f97f33818fe5967e2d518a0340dd7747e3c066252d415621522e64;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4dd2991afd78833eddddcffd7d63d7087fe0c8a2f874da1b2dc3d35efa039da8f76f96e910902c33c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc53d90b38d0b81282791beaa4106c4ca43a3481a3747ae51e9e4ff0223c4d4445bc6b269a64ff26e8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he491997a6007861348649a9fce007628f2647f4a6ff39c9a7c9e751af65c9c27993f843122c4f21b5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef4432c9abe604dd3ddcd7ea09ea1ba15912b588521d75dd33322349292555d1aefb18db5648c472c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f203b0051ef5f9e7b6e2dfc3acd751f22a5ea294c2244dc9d7a86da30a13e3c044264596b83b1775;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hafb4ca74cbec8ef78c85454f4a568b9d6779d43f042bbdc546b5382de9604282f8600ffe35b51aba;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1f88bd78af1c9d517f4b225d84c427e101383522c87a38a416e592de5343b4f9e06bc55eb16c234f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29c7bf631211266241b72030934a1d34329b48f3cb4eb6c60d1412e01f8279aa2149ee9c86d180f8c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd446b455a207604d8290422fa11494022d496bbabc0bb2fe73d9ce7a409c3c1adcd3dd079aed4e6be;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8a753bc2051552f1ddf7f2fb1ecd7741a081fd822ff14982e49a4838dacb868245577d9264aeea970;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6264bd5c2bac49b62089b4ec65b81c5125e2b109cfd1f51e0e22a502068176d8ac06245625ef1181f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h483f0d53acb86d92c86ad82bd42a3a559aad1230746bc544eb32fb1b10e844ce3844f351c75121459;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc289ee82e34360ca748fe6dcaa8e151f48e32dc23c3f023add995d0b8bf15be0e86dc2dd6cde9368;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3b63da43a8889c3a5c13252f046d8954a6d0a0131c8331f3d3a2fb8c7598320645479fe30ed824a7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9ee87b1514bc9d3726bcfa2627f6da532eb6f67e7cef332d9697d05954b74822ff959ce3408b3e9e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hafb522bf854d41381f1c9495da7ce167d862d855df389b777c667258c724d98f48fdc13bf3856b3e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h722297b43588b549bcffb7a791660ddd9269787bf89abb368ad6dc7d835f2fdcd09d485aea007275d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c917569a0287560b43d04caf29f4e81c24b855064ae85ff1f8c34c6a44c8acff588ee2bdfede7761;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9058b440dffce3c9a9e9ea2a1c445dbed0e5ec4e3f40abde8e661028f9b622149b7b74794fff9276;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1e8c6d50d0f7903b8ed86014d085860c65fc8e09c5d912d37b08c8334194c7945947f2f38165eaf3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c82a9d1f48f74cdb723c08a86a800f2f34db754927f4e50cc2dc3a6b1b067b20d7a81f283d03bcae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5460c67bbb4523efa2b9494ccf8b664bfcd65117ee1bb6ac3480365b88376ce6caa87ccab7bb659d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4bca0453780401ce1b8b46edac0e3e13de472f1e0b52f2995ecb095051ccd72a19e0cb1057bba9a0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc35b7cdf91ab7a418d355c8c821fc78052c894861c85c34f76894046d2bb87923de1513240a084c90;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7090b298a447bb699cd77608dbdf9d5359c312f56d3cb1f3abeb6afe3552b68f832ce0b1bde4f3150;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2f75f41ac52305487d4a60b788530eefbb0a70fa908f9f55f646875e748995f187bedf4c99d606f6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc8bcdac73d8f88e6189369c7e81b91a216e13448c2dd744490449c1d7419a9f41e4fb5d6bd461b296;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14e8dddd1eb311055cab853757c65271beb345f3aa6d535cbdbb6ca255bd15904b5945e4dfaf1b624;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h978741dbf5f9394627b3d3e4ffc5cb24c0b6a1bbbc53407c0dc1f78176171761cba818fcb59f68a7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf174be53f841fdc551d37acabbe48e23d5ff28b77146c51b8f716e1ea891e956293ec9e087f6a32d5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c27f9b719969b1e0ba0354a1e21e5e05fed24c928cbad30eab32c7f03624705adda9f9805b5ccdba;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hebe5da5206bb37a2da8e6e539f418a2ffda03c297caa3ffa92a0fba31bc76256ce5a1a1dbc4141e6b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd29c0bdd4641ac58c9648ef809731bc8eae7a208e7b92ce37059628cfea0a69e3c86e014ab39acb4c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha48fdc4fd0a0f046bf7f5c3fe8b97b193ba53cbf94c7ded5efa3066677dff3c5fc1cf4244b56d6357;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3395f5d9dffb5129a6429ec0b368105668379af5a588ffc53ee445da3866f8745e46ac356f60c63cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1af92e1fce0992da786aec8c41820960dcd85b772f53cf078d8fad858a0748e93861f362101c2a63;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h696d53df660dad70c10de560e38b03b9c5ee4467f5fd85b2cb7e4c9a8db051073b102996d8059bbec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfefb2c9f8e8145807777a77f20f01abbbf8b2623869c8011d2033144fd569b2a7da018ac94b172953;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7adbfc0bcd3a2fee54a9a7a1b33632ad77d659d78037620d74095632146da3fc5b6e274dcde0a1a89;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha41394646e4a3ae81e27bd2b532cf1d60a79618dc042fdcd78e0343bce952575f031dedf6a9e5fa7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3992f82bee39ea378527afa70651ce86c8e7d9294a610c434511052848c2d5f6d3e19c7408820eb92;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f68e0cb7ddf9ae631d26b6a50cafb834a7ced93536c6e04beb6103bdcd2ad66acbf62fd62cf074f1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h56e598b4f3961598e60a2231a1b7892a463633459f1a6aa4b53f0f7c1f713267d6a1b6e4bad2fa78b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbbbd0e811a0dce9eface7544894eb9066c557d55d48085750f72d35524db6cb1c5a66a7420b99969f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4e584d63aee2b1dd3e1d2f522f06e20dd14479e683baef4a00603253a14cc34777a220d46c8ed8fc7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60b9530d6c9b3a4fd085371546eefb945487bf00938c2b0282d606f73e13c61c06a2142b484de0128;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd37c96f67e7014656e9ba099f9e15b36a8b1bbe27d47b6c5584a51c088b4c92db768e711cf8206d95;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h58ad3c3b78a017af0aeb0b878b7510c1b485e57e7bbbb7ee3878c2fec77acb1594ee967ce95415028;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h106eb52f680a2f5681b17d83857f76e43ce054f2604d3f8fb5ef760170db5129e966a75f6345acee1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha2b2da069223d2f9ee5667bf00e0095dc41239598a4b937bc45275ded46b46ed662f46eee28332dc1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7998cbd9ef3a1b59777d1766070e118f437040e3c792d6464a1dbaa99074cdeade168a34bb8f10c55;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h536a1bc30bfde74ef191e724a440efe25f02c17c151c80bedd902bc223574400f51d36eea2e9acacf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2442c811be9418689c551f03bdd887f7ad69d48457dd2698137658a1f07b9a6d43c7ab532b6f6d5ff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdec0b5911210e2b45e9c305bd9a104d69e585679cc990cafbd405abff15595036458a1fe8b55297cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1244d9d3d6566d6ae3e133b3ed92a30475ec6aead1a447dd4370b2efbab9e4928d5f903e81f804b74;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6289c2984098b6eb252165f17055f0a262f7a613bc29ddae956d3e35cf2c083f55ecd4ab83fd6f22b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hede6ce06b816e4a88f0b4a836e98125e48206f10d0fd77a3d9f632c6c51e91fe4d477aba53e9e847a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5653c201cf0606207bf7ca49be83413ebdb5b95de532d5965a7c1135bf1b6b9c379086e14f0b2597;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha289046fc19486af68bbba679082cc677968a61a850281403134655adf210f7cc1dc48aaaca46a88e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48353a1933d240d2f329a18d2c13f8beee3646451b85e1474353aad766cdd782ab898adc476c25efb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heac785e195e2717f34aa028d940fdf6187e127e1ab665b61cd54d8a27099a30b0ecb6060231ce8915;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb4f162133b29325d3a27e9f8ea2d293745ec81600b19217bc0de254d8043ffb1b6f4bba6d327c49e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfd5690d3801e36f3cffa6bdef87a859fde91ea8749894831bb884a129723439016ab0d04a5519e604;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hddf6ad577a6b1c5c3ef69d13ae79b81d30cab0f4489c592560cb27c87b820ff4f6e07f71d0fd216c8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c60f2064a8df7c36549c56212136b042e1a42748a736dc1ddc7a465867001f3b3ff29ebf8a9e1100;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0aa93bd668239d3fd229bfa2c9ff11fdfa857e25976fbbda0e086e9aac6a44c4ec60c3f6fea82722;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb2fd7d826d1b15d927a6821e2f30384cde33bdf44db9e4de3a4632314c128bb22c5f24527676439;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0d11bf4e8e6b6370d2e3271e32267f0f728879a0812638e34f8f9a4003eb41075bb50010a7855c46;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha786db54f953e1125f750f14ac18c19a54260a043a155a694f77549cdcf93806e88b41c4b54c3c425;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h859bbfb2057dcb3e73280be0aba49c8476fa461bfeaa19527e4feda09dcb4152f7173181ebacedb98;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd22919990d09f746dc0b1508860b30c8e5e9f8fc73a008266f909c1b0226b0686a025e6a2c13baafb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha50d7e14c6b114a4ae173fd1200e26ad4818ba4f22e406de5de14b243f2a517e73750b362eedfec09;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h789d116b082e74d7bc5f6abae74e7a9bdff3d6377a11562b612050043547f1963c13e4ca2450c6289;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc50cc88908cd50cf6fcb28aa300e003628959f646fd78d020eacc7c36147f0e76c20b731d44eb703d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h35ff69c305f08bde5f8c30ecb33252272000f58c75c98c709c0dab77cc1d77f63d17ea06842bef39d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb8cd1afd7bb1257cd539ab5bb566f8b1b83dc298c0d602dd2eac317d17ae41a4668d85d8e6b7804c1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81c6927a41d2032e3f5e240c5b9f49ba685bc2ad380c7bad71a21da8ec264590ca37907effd2a5c5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7f8574e2c899e873850c4474214635665176e235582c5e960c8d653e6d8a5b89a7247abc998650ca2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8da4111ace4a4f76e5fbbd14e37289ebcffac677b8f94b2d5a992457e98743ac60a8b67ab9b530d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ac2abf4005ff14638ee570f4e0561bfa419a6f16ff610554bb43b4967e8a53d17cf888451155725e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba1abad8ca4849d4e09a43eae421a3abd6d5f94fc516b2a6748548fd67b4c9dad21b5fe3f18eea839;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h921b74cec82c53952a2e6fbc32729fd0bb325b392c574133586bb83d5a774e47624107ac6b79d8013;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb1d6a550c3cfe7ebcc9f8891b43d4e61613c87f2f21400cc9f52f74f68f50409fa16a671ee5616315;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e42100ba5bb0e340fe1537ccd8dcfdbf7de292032a7c3478b2dc3ef2720d3a525554b49b13e3be3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd434e77985f2d20b3a9810271181a9dedfdf9fe3dc72d3fdc046df89e5b6da436cc99c2386744558e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b464c59f9e78dc640457fa85983bbfc9f613c5109c4956b93f42a2f6f8ed33b2745519b7d3d09053;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5206e70fb53e32a4f213f2464c7aca5f15865940f3588afa4bb157f5ed8cef2c618cf1a685936b7ec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfebcb7866b613286bbc409a7b62d481589a2bf7cd8ac31edce3b9b0df28550a3900deaa9eb3ccdfbd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca7b3711643ec608129cd262ccec4083e883a61d656a1b984846245a6791e7a452374a0d57cb20091;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4da913d8a63f9a7e4e5783ce5d11bf8745c688c4efa79ae8e5319d48cd83c6111350fecca36e997f0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f343a1fb500333e8ca73e7464db05296525e2d67cab3dddb7d68896beb9df6f65a56e0c798e4c229;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4507c603ee303ba44113d2db78048daedb58a6b677d883e1499f82d8bba113ffa79d203161502ad21;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67a9660c8977cd1822386b73eb5f9b85a743ca71bf90b3accb348ec9715574381683ffe87770f4c33;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ff3965433cf4ec411cf3868cd18857ff3faf954da39db916363828c4fca66783d2cb5ac782404f9d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h52d5abe1858904c53beef6e4f863181aebe7b7fe8e8be58ded147bff6a82e2f8b71d1d724e4ee215a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3885d2a698394b75d7d3cb034c3875a85f38e2fb5ab9c9f50d23aa474482b357532dafaf8c34c5a7e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf609fd3bd78933ccd43952c851f4bef55d4618291b6152b035b5b9cdd388999df831e4250535d0862;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h737cddd3ad5ad9ae58878f596cc2984d325423c2238f4b500478a50203f1a6b54d3766763706971c2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9f8e9a7b617fbb39ed00f665346355bd98d429db921650746dd2ecf458e652dd45eae6e17160dc67;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h674a4811a1afbf22f5a3ce63bc787cdca67f6f20748cba4e89efe837f7bbd3a0bf8d0590c607d7834;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9288222fbf321005f4d7713003ce13ff5376586af33b200cf9f075b6b64ee8278e8d36f9c5435737e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc1a047302b992c1848b352f2514bbbebc1edd43063ff82ee0ec1875fbe64d89570662cc7a0606df0c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5950760b7544920f2a4b0427108342aa287020b54cbb1c0d7574a9d11b96226b45528ab70652df629;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8426beadad44c8c52f6dd1727de16093c749f4936a9165ca704423e45d906d53e36ebbf153424847b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4ba198a82061e705ad731f115b1ba5568377dd702b783d6dd0f844c6ef96179ab63f7617415950cf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce81f01cf6cf49626722946fd9b5caf1690ba1cd2317c3f23e6169d5d305a1956483b935ba5c007c1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2fcb616f10715b28106addbeb3250b6d8c5f81b31ff411a3086f1de46d7be248ce8cd6eb3a894eae6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7309aa242103e186d6915881b771e7826c98862c4c00c94bb1be7fd63a969e33ecf4244dfc9195d5a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h207b25750ad7935c963f090ae2a63eb5a4d692663e4938a42b4fdedab7cc000f1b07b6a117110c667;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdfcd65c1d5ae2a7a5ceacf2f85ed9e6ab4ba871b798f92cd70bb3c800f101bcfedafe50118c380d78;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd473647aed6c1228d371093814eb6b2efcf7e1d1155ceef50bb5c3ad349d976df8e474303f2ce14d8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h609766f474d193e7c077d08693fe3a15d17085d827d44722133c5c6158d9af7ff4073ff60673bb351;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e17a38619102181ae3b2d0fbf9a2eac70da22c0cdbdef15d2e6a026b714f925f9c3832af9e95287e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d3330a5a59c67eb81a825c9e2c0b32f242742ab66e6cc6019cd939a31c559cb219b28f2aa13d402a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1820c9f0545db591e1c2e447b2b8161b9ba84854c09c26dca33892a614f73943c43bbd725243728d9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h88db340645b6c79c51e50586cb7c39065ebb44f153cb29e92ea97b9915e7b932bedf885b783c53339;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79ed39ca441eb2b5e7f8fc7b0ebf06514ba3c11009a84d952c71348b54c8d24da6fb188c38fe9ef93;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h85a8e215b661ecc528f23fc7a5d5daca417f9246d23540b60f20e0ab76078d7dc2aba1eb23823d6a9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9a169980d98ecbab91f0073e864c2a2262652fe8292c1014c9b975328907e47790fd093a313da817;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3f9cbe718f6c15787ff55be6112e70328b1a32f2bbcca15352514baaebf242d5f8aee8c7cc47b383;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfcdad04adaa2dfcb7e60a6d2ebacfda0ae0007c33c94610670cb875979acde74ebda5d6accd478449;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h46a27c2f11daf8169609fe9c8d98f889c8bbd5d69b04eacfd37a4cb1e4d1be18110f0c5c2bb74e5c5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf10a2673817a55b3d714157f6178db8143cd6bb10b8c4f9413318829691900cd5c65ac0169e19ae00;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ac6115461aa72c447efec75f40a3372254ada65ffe160244e7afeda7f2934a907e7f272dcaaf72e3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he256a6a81a7d04007197263b895d89608a170e4286c5b5c9d56bac4cacb6c9a36275c365ed1f26132;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd31ab544dc6ecfca293b85b2ea703a5ed109cf6a85b4ba0fc0c2e371a1d7cb0ff10d73255538229cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b8a9b2b8a00d058cddea5b713f862ec5aa5a396d0c43dd9eebb66b17fd1b891a988e8f7833be34e2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe59448ade7bc84ce72b3274fd239d787765598dfbe1a3a945d8d5bc12403c74b63021813c37d795d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15ef55e7f445a28ecb39f785b30dde58bd27d0d30b8c1d877f76d08cc2564bb1f6f917db628170abb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d519ed0180964ee64cc6c3eba98dc8ac4b5c7d48ae7573effe02851df6c4401c9a08a9495353d98c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h35225e44ebb0f24ce2a0a40dda5f4844750be1c6802ffdaee6f642ad5b15d04870848aad0a632ed95;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd9e665af80173f254348e105c0eb5edab06e83cd683d3fe8f826d73f4e15df037e9c9af74fa13095;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f7b9b18dbf0b55220dc6a663f60ef2536df9aa814be463ddbeddc0cafca023d0f3329b6e388303d0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d32149e6e2cf99ee20b2d82cc5b34d32d8065bfa67349b3bed13a3719581beb8f738e69cf3ca6a5b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdca6c29875df1c157d84491a9388cbc1b523fa5446cbcd58350dab8c5f9f3ed071cc4019f9e53fb6a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f083e0204e1c86ad69166a51e6e7348338de06947023174eac9cb451dbd1a3423070b37b81abd38d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcec0c3fb7325b786eec4f36cfcfc17cf912dac7ea3aae004a6f57b8ba7d3cf9d20cae253e1fce1ac8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87c37232618cf538cb5382f36e5f77594e941f887e40d2d5696914824a5807848b786617c8df85c48;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h729f8d72045e5f31c6f2e946cb7bf542ef67ab10fa1915a300c44c6f6743bfdbefb9e65043f8de886;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16ab0413b706883fffaef13aae208487b18a536da9a4630b5bc9889546ed2cdaa7645ab924a6ff671;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7b620612a6e7467d3b34534d7524a9b4bd5af556fa48027c0daa0c248d9e37b199446b7bca253c4c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2872b24798348c5e6fd05252ee58fe99d6c48b059e55bf16c48e746c101e195d12ccc6508a783d5a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ad05b3cfce1c968713e54be15f4e361e9977a41eeaf3a40e9bcf9e09595e0ad705e363c4183cebcd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f44b15bfe12106a5e6c31209689c3972124c6bb67f1d03b4ec8e8a93714f66988cd541d0d551a1b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb539a438ec361f61c5ac6473dfcc161a296fba6c1228928d8af6e8c70bbd3cf8ca611290ec1706dc9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h879b0f2982539132c0c5700f63830514c0161161063604c5e8c4d85d0cb204767d109893adbaa7a6e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haaee2528b15307ea60df32425cc292f87c24c751b516255e04c37bbf051aa9bed66349a60a5a8d45c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf05da23eeed466fbc5c91c118a2fd5f52bf31359077bbe197be42be00d3b156a0f382981631b8e1fc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hed3b095ba2515f6cc5774740afe83929bfb88213231d0e08914cddb8470f7d69c58f590efe1c160ca;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d3f2e8bb1a85437d2f8ff0ee90d563f4eb7fbeeee1d0fd5eee2c18191142f44dbe0b7ba343e052fd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef06cf5506c694690e3c581d09dd19e4cb67e7dc66a757616126ecbf00cd4150f13c4bf5f19366457;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h97f0aebe1f0de43f4e6b0f5e269e7851b8e3efefbf95a15a06c7cbb48d3bb86c9eef3b609dbac8a11;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9b583aa10fd27cca21799296a42bad623937b3b6c7235749417bfe711cd9310d34c25130be05c8c4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1cdbce98bd03a832484ea6a1a746fcfbcfec4f352b0e42decf6197eb4c063e2c13df0aa1dc574bac0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5e7dc537456547aac0221a4bad1573176dde57f7061990b2f5cea96792d151756af90b4a9b795c4c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb621f8469fd714e66461f3d698ca3854f5884c49a7fa60ea8323012e0adfb9aba52e4ef41ee521c30;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h485cb8338be648648b6e17034112331f715e6b2cb47504e061e04708041065c11785c3fb4cadddb36;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6555ce9d50ece28ac710d9c01caf84f6697c554a87cd53387fe732c0754930ee9b8b47f09dea92d25;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h777eaeeea49a7ac99597766e4f7ecdef460344b2fe002474d97178f083c50191cf020113b93fe2e81;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0c298875a1aaa3130ccb41e74b69237dd1385b49e9751c12a378567a068da946a8a5d30574ae38a8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47ec9c62de92527ee0c73a9bbd5f0cff02de468fdf9ed70bfd41b37d7d12623c20c7dcfb6b2768212;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb601b23f2f2674c6474b23199c1e9bbd2a7ccba99c8a79372bd18748a620eefa6735fc89ad096b1bc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87fd3dbe93e630bcd2128f199fbe6d330736b989649f71e15e1b28baa74c521c9ce5445669297d26e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39b2ec35dbdb1604845850a0fdfa383397beac50fe7f929021fc3a927a2aba2b5c859e274858624bf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f60b0a5ca8616891bbb2555e4ae35fae9b9193294b337dc0c3e28485a9622e830b39090eb44b82f3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haa8ba0e686a124f323cc997d039b08154c2ecb097809b7723c2e133d71b9d1b1fad005853e4af3732;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e5653292948644f48b6e687cc6d3287bc6c2060a304ed4e9645563744e50b9449f5027fb9c09ef52;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2853bf79a38541420bca0a4a106e55cd85456c368750cc76e2459ad58617ef9db3d5c6d5769029804;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d8f51677e355b3de88d1756ac9800e058001122dd97ccda9a0d4137a55782109bc049ec92f6d2e5e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2496b1f80996fc23992dd5db1a588ca6bf1099f0b5f632d7e52dad8f1009461d3c0b2ca0ccb25351;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3656128c1d8a8a29c38e65263f805d9a629552f248cb0b7b609d8559e3b9fb02c7a76152ff597947;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h692c19e4b26644f2acc173e9d4e5d06704961da67ac7c5d9da4b482ce721ec6619e87368b60d7cb52;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11d25ab046c272c61438974986830b2332e75d4eb395f852bf9454c2b912eb8302916481e1ee7f1d5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h62be87659eaea6ce2a5db013dc0c94169edc7e9292f28689c4f0271b5ed76f7cb38d3f05e8d6f70be;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae247ff609500cfed78cbee9827ff010bc6057af61015655c5b6631dd9380f8bdb7b44029b135be4f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13a1fce7723cc550b5a41a8ae6a957c572f769dbd82b9f1cdc9906b4370f0e6eaca4176919bacb19d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8785b057bd53b57bebae35ab0c14f3d373a92a67d97295f604a6586d8f865a7eaa8dd9d3b8e2a9ff2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had6111f2f90e6b9096598e5384527e5ffa52a427a001ccbf4df8d6cc5d01da28ba12e540b3ea5ff9c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82cd1cfa760f0a3b3901d36f50915d4c5e904a09c1065c049c63400c91dbe6c4f09902738f5124ddb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39f7044165024fe004ac34668bd097d2cec8593d4d0c2617ffd80d7e70732c890f3601b4e91a13bb0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfac7abac64fc1ba83ec9e6880c6e4d123f39516d5f155e66110ef614912decf8e2cf5d831311b73fa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h35f47d92abfd374595573780ffb98ebf4f9b57e04999da3eb2d7759192be6953c433abd4ab5d0f11f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h33cade41668977535e19807e7ba929968a80b59cb40b08d9f876345f0cd5ca219745c8cb10f19300;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hffda1139caf44383fc6f9362b63db16ced6caa130643957e3f9aeedc5bdec7c530a4eea428b71735c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h37da2b972f1947e93a66fd9635919cf4cd4db93187c68bbc0c2c0a5b0983280b626b8961eba475718;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7af0831b884dd413d02aa03f65c1973b3659da0a462d5a6b179bba4175d12355c32b90422bd5eadf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7e6080fb08651fcbfb0d97385113a96af20b6f2e770dfb5656df2dff0896e31be3321e2ad203629b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31c3362e92a2f29c5d16489a4f6eec8fcbc35e2f984803bc59f73504a8ee621f4b4d15d7d940e1996;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e98f96d8789ee01dabd55ce624efb411cc975984338112c32145f6767af931be12d3fb8751d6e528;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6fed5adc37d0f9ff0d48f1723ab9ed75d3f36f6bba15887a65aed252beee5b92f80c697827a867aba;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb31c241ad65313780abcf2a34b4b1d1a71d0c55d613e4fa67ae37aac7eed7b71d6f2ac6055e9fda1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hafffc9ab1db9f82e771ee233db5cdadaf5a15bc7bf05ee1299aa12456844a2283495cb3c156c8ec49;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb157c69d21464801aa1b12f9a1bab63905edc992621a446e462f73c8d86ce20b78ad747dbd416424;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5da3a34205624d1400632883bc7cc0f22b16fab0458c608cc89bb9ef05e7a0790b90edc609665d570;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc6eed1fe31b38b891e275741cbd32b0500f2b0afc7e399fc1bfc49ebfdd97856476fd343a5a7d598;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h792a48f4db5a868a8d8c8f858d8526e8f4722a22596c1941a14164a0fbb5c5b8b5671c91f6a12c33;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he66a8baf83b0a1f599bcf62f1028e9678931d809f92fefd2180d17f05843ed232a67df8fd0bd603d1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4584a870021fe16a7c7de74d77ba5835ea1c445abfaf63c4224e2ffc8ce7dade06d40d7d8a20abb7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12872a8117d8080dc0168331569e9386af53eeaa1f22ef1619a30f108b9c7bb5d29a306645228bb59;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8aa69584092f6e4bcad060b360f7fcd5412604954dd8398b668bf6cba5794c1570878d456c10479fa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4195252cee2cd633fa0679535218d5f5a6b70bb47cd57737fb61b0020bbae5cbc0970115f9dc34c7d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6301d39f708168ea8c7322274757136715943f5a9b311eb215d5cfdb76b03de27756953ca27b9103e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ca0f269d756007d76a5c1bbf8d6261b902f875f9e91a9f2e7e4d6f0345cf41769c9077994a8f29c8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd45a95b17cadf1b9894d9b5d1dec9754df039785846a03966e8683b8a531c3df6f15430c00a3fed8c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59cfa083f439c19ad288dfad98eb29a9a86e434e667620278249118705de79fa7bc4adb2753b2986f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h183c7a1aae03c1284511cf34927c77a69d5c77f0368f1dc6dd8160154d4050942a6fb0230c809c08f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc8a3f7f11d7adcbbbd05e25563c9285bfb4704ad55ed341b12155401bf5e98d8bc10aaff7171ee803;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdbee047ee76d933f8a680c03e77cf137e7d877c46bed9dd3db82447f7800f896896ddb45b8e9b1cc8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93222cf043d601a8e362096d09e2f4c15e221bcf198106c034cf0d3fd5883d52f54b0a096c3436fb3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9154fd285165e6509cc711c082cebdd29ccb6495974417ec8a5da3c70a2e67e1d0253ade02e894342;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c45dfd268a0c6cebd2bedd4cca9f64895bf2887633c5f02bfafc3ec4921a84b7b6fea48773a9b070;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44e7158b475ce34eb2f3ac911d82268bd5d027a20d98cbe0777f58b1f7021a8719bff47ad4a3062ad;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb2159bd9761b513e211e8d27d03d0bdd49d926a0ab956293386ee034f8acc42e01c18cd9ecd9cc659;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha545e604caadfceec8f4d9524fbf555d7b9adb72d10d11a89644b31357059b0fa820652a299d671bf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbfcfea094adc528099ccb65454de47332879521f4443a2da4ce3a60d442f66658563ff1a07a78f68f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h60c974958d2e78d868a113717739e12d46d352f9ff011486647f9f1e2f39cc21343aa9716190505bf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22a4fe9717d5a6a5284ffc07208101844cdb025c80dfec73f52b738f8c4847c6b901c6b7cc1275970;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0c8f2faa8816e9e31e6d1c1f5df72b10a9520fb3531900dc1f176f3a4c24b950efc27f5c6ba9200f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h90d26a98665d15374ab353494a08966d8e1e3a0382b0de8f7e3116968f4a58842ac6c6f27d9b824c0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha253d64302682c64b4857306d377a4a0be89cde3f0941cd2f665ecca6d8c9a57835018099eadb9276;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had1caec48d63a4cc611ed0694e24f2eec70bacd7cd620fd84807ada22e64a15146c73f7901357e3ee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h971af5e12430d7600c3bb1707bafdb484226fbb384dd8d446fca52805ad989c0f4bdb4209fc91d750;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5fed678fd34fff91a9c46f563bd7376b61a72f2ffad6364b46a007fe47823f59d3abe6bfeacd5d664;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab671b374c5cd7d07d973adb7b98afb57ab09a76603d25c689c602a5a57f6bb13dc28780774a49970;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf575d22b82e4e8a150f282e4fec6f7c3d24838473685ccecd699abea8c4d8b7a06dd00c3e899f0bbf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa61c24fadcea969501740234d41a007b84cd0c78946dfb9dffa907b76e52e40551f4463dfb74431e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5a9c6f5d82738e734596f6283efb84f6fbadc511b4d123524c9712180510d98616cf169653999bb72;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h239a42a6f7a0d844417ea9e3db618246cf7db6aaa0aedfe3baf918540754aad4dc29ecdfd64d86ccd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d129d845a146c94c78cf7df88fc318a513b9a223ae4057acddd0ee70091fabe9cac638a1c9296ffa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22bee11256e794fee2b940913239f99efb6028ae30853a8dae48393fe9bc530978f33dcba4e2ea0f6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hae141907b2d67deeabfc8fa6cc13f00916793ef3b8da2dd7af4ccc68bd2b3cdbdbe80a34a8443fd27;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he068eefcc92c45f22b845449b3c32a3b541172a7e9a30bd6d7bfc630ba1f1660e03f4f31120cc6224;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb66bc3f54dbffdcae66d3b64e22f07e118c11942658398ee00bf92aca970a7be5517bcc3aa623d064;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ac4c61fb03e9e4627226b5c6fdff53bdcf7614ff6d0a110246fcf75430eca544aa6f3074f6137ddb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7273745be2b48f26cff9b31a98d8568ea3858fb2a5abeaf72a7fb64f06b7a760b31b5817a40778b5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdfba63ee6df3159cf99b95a31873c521875a6f8a800e4757072dbdf70ef5aa66ee55db25b41ffef0a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63301aeab8efad07e2a4b38d7722be196494d1e8a91f2f53809f9d9211c4a4f8902361298c9f6141b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf99ec7dcd0017f1169a53c90a3d15b31df45b4074a8caab2cb1e771386e2c0b036054c65fd9660a2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b5258c27e90b10cb49d4606cb093340613c6142aeb71b1f9029a3cb354606f77b62fa4e34b73b690;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3737cfb7f6c5ec42dde93ea76758d18a5f5cf89efd729bfa8655c2b2c400ac2ea24cc922230d7e01;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9bbfeb2223775158c2825cfa9b0bd644f65de6d2adbda6f317f04708e16d0b45406b8e716637129b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77904c1fb9f2a822f826a519de29b52576879e8634fdf92522618d987b6ef26b1f6c4633baa58ef9a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he02ed6af5ccadbfd8f0ec506e3fee8dc67bf5fd95d191b2d0dd7bcf736be9df8875bf852eb816b471;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h15b80376c39fbf3c8e0d3cd5cda7a1e7f06324f15348bc2fc881240d7ae6673d647c3685f6efddd93;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h37036b7209ee9b6ef287dd630f89d37d124b3fa58a932bf766b7279c3c00096e24aaa8ebdc17aac73;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h93614f988d3e6d9db8062c28f4b0ec4925926c2ca902bd55d6b196103ad6688520125d2182406c6ad;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b962f6f883fd576206f503e78ab5cf489e38bb4da02cbcc197d46bac009dd96f347cb046836aa2d7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd0f21722b0299cb18ad42ab015ddc23554176ee4a7907aecd38ce7ffe398839e471670de29d5250c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6101d2983f6c3f37eaa4ae3cd26fc28df528181d284569ed3a9675f1fa4618b1880603667f5d2b726;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc0080e92121eb2789413ac0d90fed57579b7e50d6799a9faa35a48fd039e5f9da1b581983c4b1f74d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b459da324c2c564f2048ddda62b9faafab2208ed5c98e156dd2c3cd1db5e2267ad6942ede76135c2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h574cf253fff82048c4dd6a71c81518a22a9abbab0d7181683a2cc0ce99a92a06687f9518778d3df93;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb506526dfaf60db5dcb85e2704b615785604ef4fd4e66f6639508d2c7a3b033ac12176b98a21c0332;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h89c4a5e331f9457cb654fc75d177dfa5fe42bc7a4007843fa6905a043c56b427aa10cda94366b835e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc0496260602b8d37be5775f8b0e82e9317d84efd9a6e59a3f937b67692cd248693223c9a4aa21167;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c472b8022fa6d44d7076b74006fe2a80d4c37b64e8d83ad39aeeecd038b1ff20832a0e9705647ce6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5532c526baee634d97e1f95da2e7ea97c6334b9fccba15467fad40a95a6790840d38fa18703c9c970;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc9ce6e36c0de7916ac6a26c10bf87d5e8b01c15277cc792756ddaf7d825d5a7741bccaf3dde60fca;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hee60d6c3543a2a24f35eefea4b457fb77f688bd66cfc90a1dfaa142f191cd52aab52a88c6782b1d64;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ed8c87e8623036748bb9ff42b38af3f76ad8a68ef11872c514172c263d91eda1dd46a78aee64301f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc75271d8f5f09301f67249595580d67ac900e5a4e162ba1457dbdbdc5d271d84513e1dacaf2a1a3dd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b752e1ffc625c2b58f798b9e2c3a4e7acdeafc894235ff00ac6a608e0f851ddb2b362dd66e34faa6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd88e1bf22b485d0344e324da157c41e80e845848252f34edc9af467e51efecc2f129cd18e2698fa85;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h386e047377e318ff59f93bf253bd26e9355be0af7ae585b0737c537f4fabdaed9b5793e1bb71905b3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc5caffb19e254146fd81d4ee79b29f729f0dca53fad5175544ceedf8af2c380a7ba28ea2677860b8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ef570f0f6bf59f580b567da621bd90092b5500cd64c3c002246562f8dd8e79d5e11e25b1e356991a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec9e68b76e7fd47c592aad32ce42690c98d5f232da2b05d5f3674be526127e80a34d2845fe154dcf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h19224accb3b4c655e2597e5739518e31f39ec1ff2890833cdedbab95b41c64c033c748a9a62819c1c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e18c8effded79cffa70d6d3cddec68ddb72b5d7fe010fbc105cfefe137647d7901bc88a28f9dad81;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h986b2a5c6dd84876c30ef8adcbdb38644dc9e2ed66d6b591b9c528e1a5ed83795eb9a98ab2b85bfc2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2292f07715df6ad971b3f3bd6e70fb647f3604f53cbb68211c24a7e34085d8a9dd6ad283afbf08efd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hded76e0239de6a0fa97573dc6d475131031e14d5b775e143fe89eb41d947c5d88f62ffd87eb48fa5e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14298bc014ac3a85a96151b8268b598a2489c7b7164da3e90129153b5c94cbfda7aa4c2670ba42878;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heff3e33f272a1a918d82a1a442431ecc22e80f783b627bc1f0a119d27444a24cbed7acf4a04830479;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7a745d176a6b349f55972805af46c3a3c9518097e8caa463ad82edfe5566455666a21bc1fd2d4ba9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb876aac37669027902c15bef08d9d702236b2f9e429dbba6a39b709de78ee03bf8b457e3cb451c33f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ee597a5e395354ec7996207fac17e35e635b40b7837ec184de4474daa2c4089b871ce7e275dfd6b0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h854ebfe4c9a04085943f4a0a64d22a2973e13e03c6a81ca94f77db8521cc6368eee26edf5164c0c99;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2db402c57fffa8d0848337e286998bede6c2ae5e7ce08311559000b90bc913c3ef3e5cf1180daa28a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb53ba6fd3789ca98abdc7df7e56918fd5919ba6a7d2d9406f481214a46619c0c3297a89ed914bc6b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc70d2db75528e9bc122ef3b22559997b74932aa314e18b2fa6a20f98edd1df63de4cf9f5583a93e7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1e7c2ec2b2c55aa7a1fdca5af441fc4b80be210eb857acc0608433112f57b6ec8c813b4f4569a440c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb40922616f00f4a59b3692ec443dfefd2bdb646d315faf4cb9094ff61a63ba62ac49a94f793313acf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87e3f565d110ecc6e5ac0d8ea06cec1347e8f2e4f2cbf0c2ff2fd1338213e7eb0d38ce3d2fcc389d1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9a63170f0d97c6b9510cf1017e366c140f7a1a1e95e4ed200b28eb9bac7ff4a957f47698f5079efb1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b0c51da1f617ff6ea58c7d93dc826ee0afbb060f0f9b6d9139f3c07037bce90838ba5781c00a7e20;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3d034b84feed36f8526999dfd816079b9431e478d5978f36237df5d1c7a997582086eab9c15097fbc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e953ca09946284d6248cdc9d20b82bb00224f87841d2f10974733d9c6f4db3322b1f4cbb24537d78;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb38ab9b47bdc9a15125e76a818cdc711adc31b146f3b9f7a5fe3d953db6e0f846b8b0b05af16a4b85;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he27539d71bc1fc7d8f58d2724a0eef08f2c212e06d5aea71488c37bcd4720956329c16486be2c91ea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31b901fa2bb540d2d9818eaee168d32659a4770f6c8129830799ec29bc1710702e0b9e8a12bc9fc0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab4c6bcb7315c82301aa7b652c17db5b44a83bb28de2f40025bb42dc548a1b93236310988c765ca22;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4eb84e3fdb4edadb21fffe89639f7c89f1cd845b862b749790994fef67000f847bfe80da0c8c825c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3149dfffbfee14b350584d52bb093bdbd3db298d2270f2b8a73d2b51276e34e0916da1f6163347e0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18bb43bcde46cf50672885cc6b2c8620d69a47bdbc2c125776d7e4b5016b4065f05824565780da2ca;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f8d1a77235c998b5c21679d0e158337bb9a9ff1c31d124c544f43759d29f685dbf88288f5f865cbb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he885806e6e05d1be48ca2e1ec9a466283bc4332707d59a9156ed87f8211900c82a2598ee46921790;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc6cb1f512874c203dbad914b2196b058522282f463d9e79dc936fe620e6b642d62c0dd0022d12343;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc880c1eea610d7a16a2d60ee8e78c724a6d8fb6a877a904be2b54b42e662490d99428e5cc9d0af293;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ae2357e8aeeeba5a73e8ac8e5f810b9270729f1493c784a9278a17966f3fe1fde41bbaf376921547;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86db21f35e157111e9f1e4d9832a899d594d6c03b60f1787131ed72f0dd38c5bbe480cea65394d03;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7a5420aea004ff5066e01eae676fa301336a989e263a0962f693dc5c7df6fbd3194b42bebf10b8cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4103f31a1a273ceef394141518f394a594f6aa307d0e551da20fb1b3c663c14bb6f6f4a06aa425aa6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcac99a3e76f91e85b60b89e15e9b54b659fba2ee9bab11ffa68037e0ecc646bf545887329ea787431;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7d675f6d33f0d732a88c3c30ec8cfca576ae08ec13a4bfc4c5915c4096a4a67d2f590f52df8c45ff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3dae31170dc19b6e2ef44c2ee891eb620bd356039bcecbd19229b68ba5d2ff4ef65d9e6f02cf05a3d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb72f297b3cc36b9b349e0e0db465e957837e621acef86f0ac3f63cc76683db0c899a3602cbfad7d4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7b2eb852b39856cca623367bf0f9dae32c72873a0b4073dbf133e1e506b1a61f4dea2a944d32f1b4a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e8e10f7ae1b2e0c2e10bba30ac9d87b3f7b40f931db7a8e126c99b383f0e1752638e2f80d6905861;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2e4e8db8110385a9565726580d3bcbd298c216ed7582644bc5dc16a5f5cb94277a4a8d04056150f1d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7434aa2d7b6bc08fe2c4707b986b3110dfe3c7a6f964f65472479c0e1ba5cda58727137cae243b952;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h868d29f343eeab45394217da379b94c5c64872559cbcac4a925d8f0b7e5cdfddbb8a31898862cd72c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h406f2281fd4b1f034fce0c46edd8b433f6dbc3622ff1e24d061a5f4152b7cebeaebbad391d40f7f0f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5588c6d94444f6b5abb34c725398dcf9c109f369f5b24a56323f565b072280d453d732867515b1031;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb9cf123e785580cce88bb22c5dfe547443f3790286c378fef720cc00eb7b5f13d5528fd60540d055;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53fa9429c7718e4e82232f64c7f54f55b0dcda823d3a346518dd1a5026a567a0c238b306c71a785e8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2b6e9c9a96fe7dd0c4f84e0b251ea6454f4660d48f2ca12fb1922aeb13cc5d8cdca0924a9341b7ff7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h26f3f85c81f4be2d845488ac44c9e326ee49762a81541782ddc0e64344e42f5a8abe89f90b378acde;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4bc21681a94f5c4ab50049886707985b257b843816c6ec36034229b847b084b5ffca93d8d06bd7e4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h554b2c92ff699ee01e00c98d1decae0089cfc43e032ce1b40ca326ed1cd951a2d965e81f64a10bf0b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab8243d7608350a4daf2edf98fbd511774a31c63683bd3f268e10e2d046dc21401d4c911611f9d1cf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3541f91891015efabe9079f344d6a1b62667858d760356c75973c5ae9e6782a7a0dde8f17c704836f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h456f26a53448118b957ec2cc8ea013ed6996e074cff1873d91a02a11bfc49c2d8468ba3e11c626cc2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1cf00e5fd9f234b0e30a4e5fc0955f1b7322ddf100563464abb7c88f42d3d7b645f83a73f553a8368;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6e361c9561ae9848ae1c4e7c4aa279fc1cd6cfe3ea68ea722e0265d590218e8ff1a37fe50c493775;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7dbc82d8080cdfe8f8e656ad894ba12360e6c496fe96508c4767d62bb047ec00aae408f9a635555e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haaee35f7da3a2323d19fa221af86305fdb2a1a62fb09711b4be62b14d9bd18c2e488ace526433512e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf4aca10a8d7329f753a1f6b33f3e8a2e7f8f3d6aacf228d0e0fee70252642472366712ad8690f6776;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47bc8c7541dfead3f3f0c7e597a6416438fc28c0f954898189b089acb01e5ea8b0083c8e5cb6bc0f2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h61b2f204b9a169553cea0dbd956a12da1700f87cffb8a329691eb86621c95360f8d0996dc040dc8a5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe8d287e59a3c72c09f22e3fcca9f7a54c79563378569cefdb27ff0296ede59038fa77826f651f9c5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50ae1e68474c88d67128b22652eaa9930d630b5f4181f40ece193109af9697dd2420d16fe498beddb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5cebf43615dcb8b3f9821715e222530d3534927bf6a340fb044c5b3bc5198dd7f19f170ec0b05b4f2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd602fc287a5fc66784eab3121c5794c3fa3fdc4598fe0b67db97dfdb450bf4b01e9d23487512fceb9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfeb6243884d44201117f17b73bad134c166b9e4b3a4eab9b2546c266a832a0355fc8e5c5fcc42e622;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h162ed166c8669146161e32ed6368618b4949b1f7ad4c1413f8586292e98a3f2f7f7f8ae659df456ef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c376f8ef2b7c59b3dac5b2e104a5d4da4513939b781e863b4687a48cc31240ff1979de4e0ddeda98;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6015e266f0e412d0d1d7e525b4ddfdbe866db67be5f4c6678b0da5306d06355b15f4913b56de9ce72;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde7c1f67faa1c1bf3ac61a2350273aa38385b46cad9e30c495ca981d35cf42efc00958cb801fb3e74;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd63507464023a507e539823ba5d21e0cc0eedffc75256a0d545f1bd40d63a8b452ea66d83a64b48e2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he782bcf7cf5aa18c660fd14ee506e6528eae112b84848d40412fcbac8f58f80717d6f1b9c87dddc32;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e40920d5e92d77683a336ae448af5c02c1e713357e7722c25dd946608deabb9da3434c439664173a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hced03c4b64615cf9dab84951021d06b8a30474d7f6dfad306ec1311379c3908abf85cde7a334aae25;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfc1d5d2e27d9f91deb90e0bbe3126aa08de2fe92058d492ae9536e2b47a91d0f2aced8db4f9dd3ee9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70208979056d09fe712c5d362b7a7e45704b49e01ded002107cc714b846c181f5aebe096f03c9440b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hccca94da02bf34e1bacf7cfe624f4ccefe5e9e35a50546e22b2827510cd2be89ac18d9c937e3c9e48;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab78ffbf14515beb347f13dfd92a7767e5581f574dca3659f5e87dc0d0cc6a3897bf41d6e42f17204;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65067c12ddf7d63dd27bf0503a49b81331268e3210c60551e87ad021dc1465481b19324c7c0ac3c9e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1620c8b9ed486a72d4b4141d1fb96d5ea11bb87d4d3e3fca916da205cfa303ee1700ace00b1c88ea2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c460d82b130af23d03844d3ada76d44dd0628ff81221000e6c837a766cf4b78d758583dae6074a27;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h87a8410ab53b42d56cc47e028fff8f1be7f1aaa08ed1aa47992478ecb0082de39c22472687376431f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbe8c84ebb617ec49a350a3b91ec341b9539c653e036570a94e8d2d742bac86c97f2d3ecdefbee4715;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf690d8bccf7deffb117bce2e5e95b105bcbef437b73e515a3bdd4fe6b44cc3603256d7afd822e9650;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc4db850a62d2292276b69444adb89902a2143d2dd78bb1d42440d5e76e1d852cf969204edb88a963d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfcb42eb83b52074002b8c36e05589db1933fe0c1e1d128ec08a14182579661f391765ce33ca2e477d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h603994faf0a3d17c708a4dd46e3c17fabdbdd5d2abd14a07b3ea1ac5bfbb439dbc2929822443dce08;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha101b18db874fd3ba65529fd9c15f3cad5e53dd1f85c493b4e3ec5640c33980a31cab44ab0d20b37e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hafdb3d6e4825e1857ef6f8cfd66c25e48d234778a08d3d5180434db08f74d3378369d8422692ddc3f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hca762702bfda2c7fd4a05ab74667dc3f114717f876d0beec4f20167a88aad792127b7d05b8034703;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12199e521fb2b6792d32fbaf02a69c6168f3fba357e16fc42689b02ee0817413aadaa0a7614c1bba4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h258b6b1cdf153e5528b0ed7750bdaa3850b10c088d9969cd4f0fa7e82c0d1edcd0830bd58b2746d69;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b47cb13cb737f2d3d5b5d630698dfe1edc182fe728095a23ccc350eec2ca47e4ce86a1e7041e0079;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h178b2dba880eb75e729e902d225ba1bb124714e055231ab8770eb03c792e1a0e55b6261dcc03901c2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h77463325e71f5d2cbdf8d9f8c28e04b9b941426212b19dbf4eebc6e7269128aca3dba238916c4972c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd1a581a03c3ad121b51eab6fd109507156e03d98825430988a24eef86d1049756dbe549af1a954035;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h159cd71362409f592859db241ec3c4b35f02ab98a6df90ea3b9cd6993517e49ef72cd2a5c4f431c83;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6fe7b64860357ea9055e817d6bc87188f54f3bcdababc7259dd0a23e740ac4888b22972015f0216c7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h70b06b1c616edf7737ca2aa55ff58bb658a47c77b4682e73161e6056b131fcc6b38d158dcf8a0d722;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he62dc80a2ef681f4ea6f8126a6db8e92b86c1051081e2c3cebe402982ee7902fb6870059014162104;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h114b761f00f022512e85a214d53f10596574971baa48cecbecbdfce6c053fdc32827bd005caf3b4c5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5fd881bf9f64876ef563b3f0f99173e2220b1c4a96cf55c303d0dcec6c9dd48d2996d8d7d2eaf7ba8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5699aeaeab8f2ecf060cccf989876cbbb3bd6a61cbbd2535241a78fbff1c6145dd2fe252c1ecfded0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbc4d630ea87b254a965d354b225299d45d8faa0b0fc1c35073a3f0bc5b964b293e9c03fdad074deb3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce7e5d52b5db3abcbae982467408d987d2f764c87b6dde8af0b80db963a9f0ce263c256ec4cf8cbc4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde6039cffea591c18967bbd5d5b892456b858eed927206d051ff0cc9aa846d71924e9ff1447b56444;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29de096f79e3078e253b37ed7296955dc32833ad193c957608f5fc390a4ec093ae44418b0d04b8cfd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb4fae51d778004acc9a98dcad20fe9282b469b3d848e3a6ae023d5a696c147f78f1b4c1f9b5313db0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h766429975db1a9ff752263d4b57f4e172f4bc6828914ae550c9436d31fb685f2554d658a8f927468b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5decee1ecf709bad5768a0eaa44dc95d80225860f2718d1b8cc21d4eed065decb1cc2e48f5bd1ab38;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h67fe068ef6e4b31cafc912c3fa48cde64832cf516a1e6d5ffb041a627417876a9070b86d9f16d24ae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9c638970d897c5337257586b7aa62ba0c44b0bad4aaaa7e35305c21bb4394ae65e45195fd8915c66;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbae8d08e5ff64464eaeca72e1aadbf95c227e5b5f8783ad4e79f1e08ee9638901b35d821e2ee7df60;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf107e96bafc6369b44344b44fec78eac74a826578df144b0f6aac9ac4fd62dfadde1c5ace2a8fd9bb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ae28dbfe30ba775bb97c11f11ccb7750e41abdf7c968e918ed1c75138218ff43217e4d02cc756882;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h493be8139798eae64c2c6a3d087d8ab193f1af2fa18bf83ddaca29116d766e4ec0a47b2fec899d1ec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68b712aad32bc783ada95a57fe2a2383bd90295910ad4c5d1f2cf853878ea02a5d58fd6e966f8bf57;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb963680ef30c0732654a6d99ddc5ac5340e151530f6ce1f6a6921a8f3104fd414803a138534702843;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f56ca16e5c756426b10cc92b225c72080a1cd79e89984b34229a4d70be3afa5d5b0f46c973508ae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72eda3ea3a67b98ca763d1df2c92d55896768701f476950f56d0aaf0deb93a4a93dae05e4e31cdb99;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f2c75c43641fd3f0d0659550609810e0a63d436109d2a1769c900a3bdaff747b245d66f65ce35404;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5144c0d281ffff195022d896d2262729c524fa5a53c955c570184697b0d4cbd8d124aafdd269dae10;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbf3f172d4efea2c4de364bf62b31099019bda8b371f3d44a1e6d1130ae9e6cd019ab1a52c5a200f6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2de6cbc95d01f8073441891cf5a1520681e6d4a7bbef324882e74c5ac4c4b0938f4b2acee10d818c0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7949712ee269461de1dab1a82021befe08096eab6abb684307f3a0c07cce8073469184e1ead92e6e7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h548c9d0cbee80a5f5addc59f27ffa274f83d306e5aedde77a03b62e8ff0e7366f6990a6dc5fdd63d7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5263f0198d3edac47ed111941e17bbb500b7300b819f9ba0a755fdbc7ed3fa0da46e0966a4e0e9e62;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48466eb969f5c6bd0e79d990d895a5378e11f626847c0d94ae7c03c95aa09c7ff2253624898f6383f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4602aeedcd088c7d0eceb358e49ac3013077f57ab9e2ef1029c8e18535fa178ccff90dfdbb86564aa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c007f3cb129433535cab8a1bdedc39af11677226cfab74aa1e45e69124c8b4074de94bdf1fa9662e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hddd2c874a44f66af8f5ccfa15561a298ee65db1cad0385ccf73b897228b18664cffe3e409fe0ebcb8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdf853a84b4fda74c6d3dde9fc88cff80b78037531bc2c036a7d86a4af4dc96fd5975b72944a6f38cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha134273531bde1be1089d5df9df6d08b5466d5b9a79bff6ec3e9762cf028f53ced53da18974cddc53;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he5078fa277dc550e396a8881ef5860c90c542761099cb3178310f1557855d0cb03b2f311a0973d421;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30039aaf3795d011ae1498d546227e81c61dd03a2eb2a9c9ecc85730c57e3ba80ed67db62071a50d0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8f07bf2d16d56eba4bdbe83cf271442f229439646cfeedeacf31107c5ef428d9fa90f3bd85fb17fd7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8309bc43920252597c7a588efa6fa655c046b0aa7d13dbcdeba1309c90cd01768f9926ca4e3df9d08;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2f12801cfa84f56f04e2824c130927f1ca5cb32983bf4f8e8783a8fc6f0e293f4ebeec8cd94e9e5a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3be93abc5c3e1566d92f875eae9e905e338207930bcbf3d674975b6bb0f0af94eb7b2c581da7c3e63;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h705f443e7323c99fe58aee6d3123eacbc612c769e92ffecb4d824bf7e21c5c7721e87bdcd911ce92c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h14929968543a2a7392b20a874bea1aa3bc5a28278b96e590670c11758757b1674c96e21e8311a84bd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb6b1e160fae074846a6321e91b378b92b270b9a2ef9528d5c21b9a5c47f8648616ffe13b397e0ce50;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h26237cf7d010f7d4492e184a80f47bcbe4fd300f5a4ccdd036cd7c65b0b24c4b4b2e33adc501b8517;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h322b16fed9d06710fdbb40288467a3151cd5d0fd6dc08db2243b1588367d9457eab7d6da9a43ac3ce;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h636c6b4cfe192134f64a4f121b9846d971514fdf9bbcc2ff1384129a259b77668b9a78136139b0da6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ec2beff26ffbc80e10f0891ce8e5361f13ffbbb16cee0c83c479bae5af145864b127e0e065bf65c0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb173302faa2c66e03e6a0e7ebb00ddab5c88d3dc5c699de05762f2223956e1bab96c34574ab22f9e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h353889724b412d52a6775fc46613f83a82d1e2384ae305fbb3e42b2bc7a0d59543800657cbdc2f314;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e9ebebe2df2de6c740eeadacf53f989f0ed683e71e8ae0498fc101276f668e2311d91a105041cbc9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36ea42bb85f1c597eb56f50eee541c051e287b536bfbeae16cafcad15e17fd01143de03cd1a985985;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h64ba24315c600c736666b28967480ff3e5f638063797b970600b189c23653f4bae4a23af9c4cab2dc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30abf4ba728bd74d0888fc6780a5d4bac03eedd4fa385bb745e6e22bdfdc777c94416c3d1428068a9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hced359ec15dede7fe2a77e10ee378bff556c857f857743ff5dc0200c83e28734cc2ff67435a1de65e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ec06f13259b90c31f4950691bbb2bfc3afcc2f6d7aa0a73508ffc74f0185ba8c73d2d37bc590de9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82df2fb3f69e6b2225243ab129e07cb95d59f0c5b1e3dc72c6760f7155b0a4913309e0b666b586618;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hba1e50ef7172dc9d5daeb402010d32c9af33a3b6fa4af0963755ecaddaff319383512bbabd5d7b71a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hef04e07a257cffa8c53026d9505bfdc72d2a7324420b7ceb69c54f1562b0340412ea67d38b313460d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9951e347f32093a6d1dc10b6a5f64ffa1d6cd70fca2e7ccc8a4de4f8b6b3ccf20af874727430f2354;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7240befec429da101b6312bb62d582f7d8ab7b5e0639bc637ece47a6e60badc2ca8317b4c26106a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd0a1c642d7f633a4852ecb9f2fb33bfa04841a3500b051adca2259cbb84809c0681b2766cef23e00;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h80c304af3843bf78d2dd4301123adbfbf6ae58e249fd87ac322062134ff5cdd6ccac447af6b17beb4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab0bb6a06e9689c174b46011cac4f6e604d150e761dfa104fb208187288332ba75cffb6e54a5b65a7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h963d2645869eb633384c0362a93cebbd9ec5984b93315c34bcacaa8b929980b06c6a827955a0a5335;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9adb5bdf41a800d09f1dbbf84ef08def4bd3772b61261c13120f019a6ed9535b4979fa4632d723fd5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5b66d646303c857c33ee0ecc4b612a0be3df45b8719a91a49f0ab98a06fc04bd7d8ffe7562ffe8d6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf057533ff2fa6671616cc99c8d638df7adada5435515c9e215cc827f6465bb0ab4aa389a6e6f2820f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3ff371101db3b2ce328a131bf1cf4ccbc7c7f7d69b146ebdd258209395290badc3146c4667ab1584;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc23c2be91c91598873d3287bfab33d902f2569b9b184b6fa6ab118975f9706377dd3dfe84ab06e3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha4bb522b232ebac1068aab66a29d584fd44e4c13af831bdc3ac176a48d788d7dc3d6dfd8017a6594;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hff5d95eef0f14a51d59fade2e99fcb871f23467d4d233e109ba7016ba51f63026bee366c8efa387;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha6feb4f5905db4655a8772717085687bbe20e5565781f2a37e6464149cd9e249a2c6618cc59ba70b5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7338d6f3ad33fabc0562219ddaffd52adf717d6b91492727c7908d866e5b2c2756cb8de4514daaebd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75fd15058abf5885df3fc6de9ece6acb47c2dec5e49e5697550d15fad6083a10481016a0a5081d0e9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22c98f8336e570d07de6d93ff8b11cc8131b54970a2111b31b01431588e7ee97f31099f564b316221;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha82e80fed0f1519fc2a02c8670702ce2141f66ce46478d341307fbe6118929802bc1d54d65da52b96;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h670d79a2e61d8b9117e506633d3e0776be3d032d680b13724c68d721f24f03266edd046a604fb4252;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h648fd425eba495a0c40e4254eb4d2b4ba9de455f3b52e95aa5d388f6cf9499d105d9a54b038dda8a2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b760b4e4c07a290a0fee5e8f834f9f29e3188ce9688e3e5447a7ed4a5bd86ced570bdf0a2fb20cb1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h919377facae957dbcd4ecf0a8e3fc96a42311a91018f92e7756784c662d497cf48b9e342c2e78842;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd22fb934e4fe91ad12c173f1c313963de16bdb1eace54e69bd3c14878424c2297f45fb743c35d9970;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9fdcc6b078e51118d3b56bf138077f01cf13077cd8a8fe3431b053fddddd3327adeecaa51f2bfc637;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc201324e5fc8fc91933bbc86aa0a190d5eb7adb0f03c5c3c7401ed4884e41e3363706145502bebb4e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4bca8eb20651321d7672f52344b7dfc4b3882d3a4b1866a281a2a90ba959dcc62d97ef06f89f59f0d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb8f4b3daf46cc05e6e2545ed656cb52f76b2da687932fb5fd44dcc9da161312e568c08056219638e9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcacee859308ba47e577a6f98bb9c8bd993bd141088e59c3d94656359075760c0698610e0f738a1756;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hab9c7836d14b2f39546380d9c117478b16dd9bcb4a41f8b515239333b01fdd345d3d3d275167fea2e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98e98f1dfd84bbe6d5ba8e940a4dcb4f1e745d6f30c23444e57339a190e2dcb0578ca20f23a0892e8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12093f636c3d3bcedd433eac75eda8481afeb0001e00417d3bd7fede63f42d8b42a2df534f8519a47;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e5d0f76e49fcca68d83f2e95702ce0397f9808e4008ce7f555e06bac64b39bf5c316e9bfd15868aa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdefe9342177d033f25cb31f929cd3423539a57172ebff1464e69db5c4ab9194dd3dc19b56ae8b081e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4b682d314989114101a4afdc198f715c160e3e80b0f382e9a98813555123ba40e16bc802e54e0e0f4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h221203ecc1ee6e8ba57038cf907dadc2db001d360a9dc7a080ecb3f9bfd9c311f75e4b4a1f0e69a01;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf6a8365b4d74db050f95f5248274d6303f69a60e1a09b45309222702f6dcd9f9a1120001f338fc55f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hda3a0ac991b946bb7bdcc2fede031bed3a8181ce35f821dd8b273f17f384a8ee23c07dc4ff197d0a3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb2bc23d09eb6944f8b1ad10b9c1b9cdce666bd82328f151d65ce9aad66d8f99804699e2cd7e93d3a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5b3468809e4454aafe22428cdb0e4574a75aa3244e5caa22bed6bbd74ad62a403909475eecbe29cf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h172984ea50d9044f25360b0f8c652f65f80898f8eae7fc13c4edbd2413ad80189e22f600f65e6d0f4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h967d5a592b942005cacb65fcf2b50302e32702717e427fa6494067616981564382328fa4c1adf2202;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h257a8bfe5234509d5138ac71661d73ab36e4b2ff0067bcafafa7e7d8eb69ac1955747bc41c0d1e1e6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf1cbe816ecb4d1781d047331fd718f84d52bd9820afb8deeaca1499bbcfc077739f9b83fe4a893bda;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5af0018fd3870c57f4a5a2630faecb8937def2f0a8396ac4138b83a093793f672041e5f7c6f9b55b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47752a8669f780a5c548811b0f8c453ae643fd13957d1312b228f1c0f71c19c59cfdf54bce457d1a5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h684743f2e5910739cb41b52ed2e8adf4aba180251b5ac902602c3c42eb6391b55bd1184667b6b1f75;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9e1098b27908bfd05ddfcb115963cd609908b3e7da36ca75d95db72d54bc028b4c2cf95fff44ba13b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbfb6736480797b481c7e9d835cb376c7e43a8d780fe5bfefd550c46559a472cf62373abf39d978c6a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75bf024a92e8e4d2b1d6574325d2ccb9f3025b85c816171533c3b999448cd6778e52dd712a24c5ab6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf0d9bc40d24a647882f109d8d28c78eff22e9e4cb238d2cb637fec3b5a0457a67f2c24dd641d69b03;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f9aa6a19d99327de680ee7fa942283d0d69bd2869ed4aa1189caa598b7d7d17404f660363d07b3c7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h477fa3f4cd010963ff4de62833dec474df8b25dcb2ff8381f19a38b150cce8b720d5855b31c4a080a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h920643526b30301e333977b0eb8a4c9103f9e0b64f766e2f588a01e4aa530ade49f9e1abb3ba9d340;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76bd612ecaa209f2ef9cd95ba7d08e29297d45043867754ebd25a86aa0c88cc43881cd2c256ed935c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3849cc9af81c58a1b56a7b654247a3d5465d96072e56b63e884795d142b660cd3f0320ab419de3e21;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd5c2061020e83c40d57edd62efa2ab9cadc6592ba3801a24e47acd4ebeddbb72040ed77dcf849c4e9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcb62c0b056e838c808c00316fd9de92afb8b48ff62b4b3b46c3a89c41fa223063a4913e109283b100;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h401f0466487a7e95cb17542bab73526bf56c26a2e59146e556a39f52491b31c0030d93539384f94e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3859b4775f7bd13f7c54fb70bbb8d99e2dabd9ce59e7d9876a0df86133cc7979a13faa367c7af1996;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h285aa16de6103c1db01a3fa3ee88a8aa5e320a2cdf3f81d5bc89c2718fa373ca2f95f26c97e471614;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ef8437de2c9ff4cfa72df25d0a30428fc83e91ce3fbf6a6cb5aec56b80d9b4217f3087398e3f533c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a794152a3236626aec373f8c4eea003c212813d99d53ebed29986476b9fbe359ef18e2bfd63ce918;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h208bf8513f10a8805e20abe44cfe1fecd0c907a6981194629e85657884026448cb91c02aabbd5a84a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h978c2edd3e53fea8e748befdde2820402d66d72db3717d4de938b7baf44775f49da5154da1fde3984;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h84a3bc43d336d1c6ec5c3eb81d874b0efda8cc7dc848797d54ae7f863dbf8b550018ff409eca78af4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hacb3127de38aac92ee3a424106553e05c02ee8dd41629c6870887a04d96106049c757c7df525d2593;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a8a1040215a1186b7171a7fdf0c2eeae1e1820e5d7b6742f237bb7b31d36b63d1fca53a9a36600ef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5e57d629b4b0073f3bfa6cd0e7e7a5f4762648595c60bbf999ecc8ac314663573b3b9b0b46fd046d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb56f6245178ca7c731ee0ece18a5ceb0fdc9d638e779f25f9286b5bfa92c467042beff5b42850f842;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1adbcbe769a6fa545ae37a349c92dabbd18e49cdfd84b4b95ce4a205db9a3cea261aa113772b6eb96;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6b2bee897b13e12568cf02810ff07bfa5393f48146361411c9a5fec32a536e59c103820720f22bff;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha76945fd33300386189d62f1babb2e9110b41dc36ddf61b9fa390a61bd437473f25b2a41d5108ede0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf3f93b586dfde545c1e9feb89913aabf8ec34588a9b3cb201a160479c9c63fd9032d5e87369d949d7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b7a10a074118b194d5b726d063b88ffb4ed987ffbf0eb841ef027b17f828f6919d5aae3e41473bd0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h726756ea04b0376c4af20ac8a85f614734eceff3b2406d3bdc90e25a6f4f98250d51fb026f556ed0e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f72e3185637da3343a837f15dcd7880acf81ab6fd91bdcaa63e46c2544c664243241e2deeacbfe65;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3fe53f3d6409bf61dcdd5bee9ac577ed2f756c44144dfa9affbf701ca371eede711a667c62cb764b7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68eda8cdaf9cd6a718973d9eb08d9eb1f61f832f3cad849bc7f01cfe8c68e8fe66945d1c59d62625a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h65b6d80b3592b7424c163e52d28a666e784d9233ad5122e4394f4b0e604f52f15a1d3c6340b8e5499;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h488bba552bb67946cb539b18b9c9d9752e344539e09a35e931fe9af0a5bfc4033824d0b79a51bddb1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h843676646ee809be48826608c4be1b010100bfcd4baed6aee86b206f61cbb207922fe4f63be223ac9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5efd39f0abc8060440f28f3c339dcb9b22b6ccc541c10c2a7b2bb30aca2672e7a59331d5acd2f17de;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5d14816517b6fde0e521fdf2bfe71fc4b7bd808c46488e0361200855016d019a590b60749c03a487c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79c9d4d850af07e183405b03685ee4620c1a6ed44cb0db1604672542c5b75925363bc5e674b1240a3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc13a0ffe3a20cbce94171dae4127615dd8ed2f61e38cb93b39f7e9ad12efb90dbe3c023bf71056682;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16786e495bd8829d912ba83aae23b882c0f7301a8fb85fc169e64e470aef80cd346493653b73cfe4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9aa9fc605247b8140ee8e158aff6e30ff8d239b5cf778e21c46df05e3803bcb681ee81ff9fc01cae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d94d747504335b5917241d0fd6d20e66906493eeeba867aedf4557d33d0da6b81b1b21c0d7b874c7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd923524eeaa8a745d9f93d3f0790bcfa71419eb731871585f7be9bd5a352bcedeebae591d488f93a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h42b74b4b52ea80f0d4294c94962ec5202ce49e5e234a59cfa3406ff423583993cf5fe17439cfda9b4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9381ba60054f5f5d0acb2b2c222593706fe0a9048776dd42071acf2e7db2ed5cfddbb3445efd2a1f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfd8bc2d35dc70b5e1600f91d691d2a42a3d54826ee8f416cacd7a7f51248011826212159fa0449881;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h71127d9d87aa9389090e6019491f98db24b3944236d1e98a3bb4ae69680926fb76419c1a82fee20b9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5753a5d981464fbfaab3a531db7c461fe8e594aeb096b91f26682cc50a078b8d9f6f03f74a070628f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfbbcf700d247ec16c17fac2591d665acc9029f342bd2d7f4f7ac2027d1115e15000d9c125a0ad111b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3624db6f3610eba1dfb9b3c0ca7698767d26aba0b65933297504811cf1c5850b86bb60f3456bda337;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf55349c0954d06a9e63dbfb9ec37ea25f7601f9398c60e13595250866fb38b9cb8a6be3817c813f13;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdeb667db1bf41c46c776b8fa86541ae721fedcf0c92cba487404262aa3e2bcd2b12522a0ee670f0c7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86a5162a063ba137125bfc99e09e85f55277cd694a841569d3f348b3bad9c9feb640b86580f2c0bd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe85957ff81a94b6afb56faa436e82c05f3857157b0a5c18648be06506f70f4fa5a01b98cf01b145a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h255a79fc8ac3b11fa7228b1a29a224f02f5547e83d85259cb36220c6c1277f0f72efd09e40a1bf389;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50d4335897e0549873088554642164fee67007f7bcb14e69443f07e99400e5d680b7951a96030f030;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h443e1997f47a160a30a842bb2567582e7d70f80ef05a7492265b33da39b896ff605377a5b8654ed74;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h66c9f713b3169838ad5332360fdf12412c93b05f20d4a1a7c63d96e036f1f5e42b714bdd0c05120ae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd59cbc6f305318476e4022e333a81134022a0090b6c76f1ef227ab84dcb903b94a9d85c227a4f1244;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he676ad2ad68fa91ca32baccda3403d7c4e243a595bee6d16b0aaf36188d75b25435647b53b9005547;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfcec0c664536830aab0ae5ac7f84a39203642ea3416c9ba02ad4188130ef706a7cae0e42fc2ecab00;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h459752f4b6f44e50217977bbf995536d1c3d6265160815fb171537bcc436980903aa8767a9e2d11d4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h970923f2ce9d55101163a8a639387cc41715f21a89ff254e21d8427664a9618ff8f9878bc080bef5d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc646476d25276d690b31472871d91897fb5ef3e3b8b01ac88b0a9e096a624d9f7fe0fc8d3475ccda8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcda788373eaf1507de5dd285e4aed3494e6778b0d940d3aca2a8d0acfe2d55c9b40b9f8cc80e153a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4aa4221ff4ea167350118395ca0ee50fadbecb832b897f1efcbfa9031b7672f2b272802eb6c137e6e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h787cb5af3340bf96237b9a8f438c4a2115d3b7189c4d5eef91d810a7502fed330e3eae9a85bcb2536;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72c256a5d64cbeb6add675bab12289cccaf885928bd7bdad968b64c63ff4cefaea4eed460f09a11e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcdc299982edae497a9d9e05e6465f9a9bcb519d943321166fb847b7fd2ef166f3c80d819699ff2136;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18eed4ae7b044f68c9ee3a252de89e461fdd786e58943b8e5f1fccdd31ac9f5cf802ef2cc9670e759;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f17add7a9337bc4ac1c3232d721f9fadb0fc2249494206f0c05dcba28cf54126eec8dfdb0514a5ae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2258315c088e06b8cd96b218c20977baede05fd095f5708110c543b76b9ab4497a75020fac9421246;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h49b893ff1950fe940412fe5d523fe80a6d59accd2b12cb5299f63e4e2bd63ed52586a1c09c7acd7ae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c8c4cceb2a38d54da92aecd0ede14f399b9c9ecccff415e48f3199c1ef637b757893918e0ef42dbc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3424e4f7185673b5688cf06f62c6b2ff93f101f8c216aed407c50b3dd84b5631c114e4006d62b3af5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h873312841a44905a9e6ace89b15e997df128ac04065db3c646e620b7419be22c8383ce848167deaee;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc8536ecba0c4ca9d160c8bde5b0e8b2e9ef9a7913533957e2c4baa42b597eb57b66befbddbac8cbe2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99f6995f37370b5208c81d55a727ac845717137defb35e5827274baf5dae1ed7b2c8e3d000b375bce;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9daec407b2414944f84704b8a95c7ed7d0168a0a126148f276dbe2991802a740f1954561df6b9af96;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h43ea1a887b05e7922d0396061302fa05a89b69771f4beeab1b115ba4f85da22f85aee6cb2f1188841;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h558120512a14ee519fe603b8942a0bd643a78d25c13d5b1d4b492ad4361cb0ebe557884bd2ddf9182;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ca0139f89680b36c318543e81f658c50b6f03baea05b35316e21773e8fdab98bbba749d6832414f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbfb4a283d8fb66e8fad5fad10afc3f5224e831c3b44e03899000ca44484670090b12742fa36a36750;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb266d9bcee33c0aa4e1c9700b526773436e827f9101066fde60235970a84477e4b0339ee78f2683c3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6954211f527ad75102f6a1ad25ca48cbdcd9898e6b8906e9794cbbb9ea1469e026a1ff705719b0b6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8aff7fbe2c72b7df8b314ed484bdeb97316c03cb5266acd731cc4156bc99245a2951cf79c4d44fcb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcdcff1362dc9bf5dce067e43bcce87333634d1c2acf4ada1c32c2d0bb056c26955fca8911c1814d8b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d1f152ebf4275cdf50b41422b2a3c6d54eb1dfdc2e6787284a9af96f69f1074a3707ccf467fd47b5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha2f8466f2d1f34a0385faeda5ee1ffc0a218c5a3225a0a61aac8dd38b5f2acfd0449fc2441d747a42;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haa7870bee91ab98cb34efe9fecf34307cc333cd861c0df8b58df1d7e8ace6d01db74aa753728f401c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6ca33306dd7d552c419a9785f88c0dd351ca9913f8f41f3b6517c6007ad61c4e03f564081cccc12f7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1558793997a03f62ab17945097e4177bdf02f1bcdd7a58cda91df9a642cbc7ed64d09b79b704b89a7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h86434caff645b9a0f157f6624c196834673a42a6e5881d68ef332031026d420b2d744ac2b94affa4a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h33c569604b33e32403bcc2d968ff2f54f0054347bf4365cff7fabd6d2056600d92dcbe6892f8f53a4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9edf947134089536fbd419b5c5e80b83efffc1501a881ca30eae3ff2c97ec1c6d5a4e725f95230ecd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8c21aacd9daf6179584f035d4e2a5bbc583c683a6efcf6c23b5500be09cde76c199cffe44bddf172b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c45cc60f018b583910966f89312b74a3ac5798028c5de57c9c56829aff96f2334234615db6efac1e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h500dfc369e80063a6367066a9ff3c8898bb3960e83fed9cfacc449864d0774d1d0981639ef682639f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9895176ac1d85ba0e1af1b004adf3d9ccaa9b023c418e3ee27364c5e8cce7b351d2fe432e1f2b9b6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h96f5b509117f569c81950d584a2f3fed01f2ebc2775b1c63381040c4e133879941f23a8d12c1bae99;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa2583a609ac080840598c8401115a3d1677624d43bf0ab5ae709a3f22bc9eb7405acac2dc8a4ca04;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39c0d8635f7c631dfa58e09c67020efec3167482127f62e16ad06d78208909f67a922864e9e26b52c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1208ae8163f45e17ce081e720befd12109cacc1e1adcf3e053aa81d50d5f99f2c4544c3851e4c525c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c62165f8f6a7e94454540ab6dec6def4fb1c54e45bc4e691ac05beb863aef9d3f21e01faf7b4a68e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44bb9d53bfd51370ffc4a1bc2d271cd7ed6cc44ebeb5be2980f016aa3792c6ddd07162471785dbe9d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd37ba4392695e13ea3fd6e4bef1f668b0c0260c7c07a005c097d9c825bcac62b3518ba420e2fee16;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h91c0e2659469d52cde15051ef618b1f56fde4a02de14aab9a591851b72f8c31bd952a2117abf83010;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44ef4ff6a3acf301cce8ec7be5b549927f92aac55fa62cd7d57f7739389bad659428c0667b0042487;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd19527b8fa19a23b4c9f579ebef9c1b7129669ae7dcec2ec15ccf626fedb173e6c93987be936f1fa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haf563241f97e38c0b78e0ee8d81ea0595f802c278027c93a83756a3fb3a7b937115382fad72986455;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf55c98258dbdddfcbcc273e6c320c7a66d4594852ba8d73508c8b2601df9c3f2a30400531f4c25d08;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5c186d160047f538b92f2f8126398806edfdd8cb7afdaa2507cbce154941cbf23f576eebc9f3d6d5d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he5c66b7368ac026b0a0a14cab77ce45e554334b70573e667d5f7705c8db3db98c03d764a3f2f939e9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec56cddab178ba00c2d905ba0f9a1daefd771f1d4169d37f90255e88672a46927d2ac93a455ab8568;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h98bd1f1769501e042144d3a7f1361a7ebb2a6d1156b42dbd87a2b905e99534e2f5a6333528c1c69c9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6c241c1f5a47f5d0f6aba1a275a96e1868ca56cd3b2872b717088cc7775976e826d0ecdf6844051a0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefa04267905e9b759d38628fc37c0b924ca1ef4e17be13144aa902164490c03787f85be59f9ad95fc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd297ae691c19786ce7c2653dc2f07bc40e39c239e3aa2da563093df2bb70b0fa228176e5a43560d1a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53d7fedaa8c6ab0bf15fd6b35fdaf76919414679da5fc7a37f7cca0c6ec75f4577d15af6032ff556f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h10e464a6265bc4b9369669cd9a7f4a9c647ce2ce10414267c6cdcac744b3556cbee9edf9f3f800660;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb036fe680eacb0e5cd40e58519502d7ac7a2df963f3f52cb34ad7ece3cf23d4462afb5af3e039d9d7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e0ed3b8fc62a640cd32e464a9563d84f2e7005869d3b11aad9f4a942a3d0959a62a75eee4bc36bf9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h16dd0df8ad3145b228a4bbe86af6342ae0874bb4f2041dbc8612f2fb35827eadf4c943c914506ae7e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48d3ce5d4e87948440c9fedf1b38c7de081a05e1ca4c7c54d6c3e9a81cb3b150ae635b1a95b5bc1f3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ecb22c4602999caff6714bb06c2841127964ffa1d01f3f7249c3d0d21d74d7a09190064b2cfa64f3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a439fae3176d365ab4bdca6fa845ead90311f973e6ca206513292f84d8d5dd19c7dffb61eeee4aea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h55450438c05931dbedcced8696195e2326188293763eec92786c9ec466d3a08752a165ffce3192388;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbba4102eec11e56b15f674b6227f7fb105d9c1298c7dd21fa12e8be026f86bc3405c2a45615969be0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5bb783d144258040a4a2e804989017908cabeac26eed9bd490e41ade19c74679c18d8f5f89d1bf1d2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h21f2efdc62aa9b4953e621c1ba368c658cda484a7453aa40bb73d670c75b87e0995aefb04446cec0e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e9f1fb9050cd3e764d0255ca660f91c9d1824e1e1c59a6cb2635dfbb28ef087c5b5da498ed28550e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h33ee4c6eb62afcd0072c0848fad8f910da4478df306167f4d46f426052d2234b3c614ac8297451c29;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heec9d97b3fb1e77cebd653406129ebb7fe36a7ae50f00da159f43ea5633b09c12af2904f392ca954;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he5a2159f51e69d63e1f8cdb5a44312d429f3d4a7a7762f5a7f654daf9b8d450566489a0e7667caec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57d82a49fb0fa679db28709643c49c702f6d222e7acd5433e05c474913d8465bc1911896cb9441675;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4de173e2650257000bd95dae410a94b1f905d3c08afeb16a7e8773aa724a97556599b8548a2bf3c8b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4169837cc48521be753b4f85e9a851823a8e3cc8c4154b2a16b1935fa5253fc7b4fa7ef1a3677587;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8109aedc26a7df3d3090cb210c5250063338096345f7f148d61fe62ac411ab3936a71a6863e8be208;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9bae986ae8390646a17434f6084ac964e2932f9424db386eccf52fa5798a6fc5e84ec4b9a0bb7339;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3050e74cacb67e5b6533927bb52d3cf3758dcb4704649ad408a77ee10dd6c5121147dc6e72f6e5ffd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5ad4be7927754c22d5e0f970ce01893122500d7e058e785842b80bc3211ad3078b702d59d4e98455;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c2b0c1353fd4ed82e007c158ace10e28519c03e48984fb42a3232e0f6041991706f0f8c325d5604;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha11b8839fbd57d23ff38e7bee3c58e723c2b94a0513373449297800677e74066b66cc28ca6cd93ac1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h251728c8ba6c05721272979755d222fb813f1590c60900b6daac9190fe00c7ff0d038b3f0df08ae65;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3df174472ee60f59e704016fc9dabdc24d64fa7c8793c6537a8ec3f611dd459e9993cce1232a39cfd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1d193788fd06325646da5a662ea5019c1db1ebe96b711228c9f60d25d3a9587887f61dcbaf783221c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha814073e228075db3a4ccb12dc9bc0dfe507acafe2af9598a9e3c231e4fe4d3196758ecb1f3dc99f3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde3d71f3d34013d11a9d9ca09197eb2b62fc3e306cb7e232b99f8a73cd18e26dd2dab9474fcaf185;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h166d2e8d2ff9a1d510add747372d67e7655d0a563e344422c7375be9e7bff222fbd192d678151bf12;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c2dcaf790b008aad7915e56b026cb179e0ab0a5481c1c62754421c3d600b2feb8c772d26f0cc3a6e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8ee68aca7c25db9e805498052c41fcfbb9e1814e5061ba2295dae29a5dbd5f49ccff9e95367c93a05;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d5dda93853848202c1e125bb7dc1350057c50ff729a87d0fc50ae79cb861ab6b5dac1aaae463004f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f11320a91802a77492285ef9e7198c5e9b8f49c255e9f37275a666013b96216b85d97a2198a213fd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha08d88e2eca4dcfb7167cae67f9e3564982f34b97443c726f97a95be76191be53c3cf49d535844ade;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1527ac757d1b550f9a3875256b978d3072a9f4900ca5c9906663487ab0af5e903f3580c247c630dbe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heaa711f35da7dcb9fc1438e57df9ec7ea1fa547a3adcd5a343e01160b380e69acde614f77ddac6eda;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf08be3b08d0f142b2f53652b715539660c6e4a21214dbb963cc314f8771cf0aed3662180cc4e3b711;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3baeb8f2749063339a2c71b59ff2e62f6df53303d1eb4ea6ec2c167b77a72b72ca1e06298bcda332d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce66ef655274a9bd6cc3e978c21413dc9213ade18f33cf75b18f86337aaf3a357547c1e2d786d2caf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3621df50a4b82fa3418e904ad86433d44382d97bb185e004beca9663f80b6b92e3aff9eab0568b91;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9d45f7118cebda0b2752cd7921f1e1af87c69dcf4a87acf588cd3ef27a699bbd04a0f1550765dffc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h41138aa0bbeb6d71a31d079fe8c0c316defa6aea984c09b19a3ae3993c6b09347e71d2e6a9fc17a37;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c50c51b1c2471f337afd19c7a4968397f7b605f9a990e7a5acfc8fc790e5deb99fd7146128e75b05;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36e5fbbdba6898ce65ea2f1694e16dbc527897feac3a2bb492420d7ea3fadfe48d83713e6c0eec02f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4bde5eb3826995c9f332d856102905fc85b4b02dbf43e82bd14f4f56919137d44cf3df89ce50e2d25;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75f8d718c8b42e4e14bd5827c550c200c87b719b6c8706aba782e19acd14414491b7a3efe4129616d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h53003f384249dd27855ffb00d9924dc40d9b3762a84d4b1d255a244e7bfab328a8cddee1d406026c3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8b35736ffec27c8cb86fe356310bb19a199089f065aa342dd14ed8ec24de76e759eb1bfb059812e4e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h559ae4eb4f357352ace96bb7f2aef1a0350b6c45b1813323579ef2d770ed5ba3f3483bbaadf89907d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfefb136bee4aad8b58f19796799af8c0b145b6941e3665b24d200c83acd42c0cf43a0f791692708b3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfb61f04a65f267f039ffb4b58069d7f16d38bd610eab8161b8109fbc4d304ce8a0c7d11f60bd699b6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h270bf4662782b95a2d68ce286fe7c70cb35f65535f1c38ea145b80e1d3ac3396a746742e5b6f7d08e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3e9bc5f3cfe7e21703d0bb644c92023335ff1452aca009d1a63329c85a0e84f5a56dc7d37bbfd9127;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h349ea0e0a4a30564cfa7ba598e16367d7b02450c32a3fe4772b5534df9a20b06d40c56c0373aa673f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79d87084ab6375d331949f46645ceeea85a5f886931f953ad55d0a77087cfaf2cd6e5d3eef755da9b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8061365939ffa7eb1458542006f1de37f6524bf85ded394cd7f764c31c03ddd903bfa267f230387fe;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99c2739fa7c4e06c6c569b8fb8f84499a89ec38a8784aa07f98295265250754e8859af90c4f154e44;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd030dca6cf86accff16838938d653e9a477fdf0dd50efc67579d0a3231a6168a0babf53897b2f4f7a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79b5ae0c5c9803e621ec1147fa8ccdb99e1a7540942e17a07173e7de36b173d5a917fe71442b07003;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2ca3d7f420b24f882068849404c3340bef23eeddad9fd230fdced0e2b3b72271b792a33e09ab5cf65;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h671bf021d81e46560c6de029620acd0012b7331e0838908fb8ad9d9acfda657b8238142468dcd6a98;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7befc3a5058bb45be03ca86aac909297a2e9917aafa6223a21b48c3e88e609b6b780ae92f1a7db5b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8383bf298ea91a7b26bfcb8239ebc80921fdfa18a83eda35f00dcebb0ce3b2930d599191bd3999bb6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf7866c13f159f975319f93807d86415df9bd608326d08bbf1a79faa7a9a931c5126dcb51981a77133;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd35285ee825a09283f6b7222c2d4443c58ae378a7fabd2e5463ad6b7cc28851ea3521eafd262d88cd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a7b2e04ebd691bd1d316ea758eccd194a6584583769568a1808b00435bf487963eec0e947a500d91;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9572558e6f8a03ab3211ddb3c15e891179b5604bff654cc413d6fc926dd65b27a1fdf42f0175789be;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbac5ee971218225eb603038ca383c0302b18b80b8888436d6a6b6d47eba08056a08dfa40152e9a76b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf563c4f473ac7a970c37c03f23b751aa7c04be26e3ce58099f5004daf29e25abbaf73fcb8ee2d89ed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e1bc08901b6d0880f43ef1ebb655fc8cde41de62ef90e9a0dbd182b6d166ad47c950b2b85d553f3b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb7bb41cf3b44bd1ef222e7723540103ae7b20d68e515b27ace5833e39193fa75b18ad320674d00b8a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99d749acb0becf4e4ddee9958c7cfc092ebe124c2dec757742157829c5d467302476b83a169e75476;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h933a2d1f241e44c4fd25af9d2d3f43c1b24b8b8d192d124ca8994bb84e007ca3d0ec0396ae6b80629;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd429dd42277d4bc7419ebf2bbac9921b224d05f3bb4d8c14634caaf853e42e24e775e4bda30328862;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdeee630a9cace6784ae6360b6d54d8b00898a7c62a905aa1e42c0e7edab1d556064ea89c48a762e0b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81bc21f6d30bda7616e484c4aa4e4af59c5806c38282bbd5446d99eed0eeeae81566389db144d2fb7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h12220b0aaca6bbe0f4176fef974f4d320ade7cb69a2cf35ba61529d2856e80d7b1a3edad3fe39f53;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h130b7966417659dca455df3b1484832573a87496a7b840889116f81e7972c25ac392e70178944b24b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc3def34ec14a04ebe364adfd4ccbd594f29772577adf2609761816b524e1857e43fd45557edd395b9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8830f4841c0b1dde64e33bbe2d67003565df7e3a7a2067c698aec4fb3003a9b4af341c642f1194428;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb26351860a960d9803ba7fe398387a0d8cc49a6b7bbe12efebf7b0959abe0a7be7bacadc38cc860f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he4fda06d3e450b78441e01ee6c9cbbdad112a1079c3f18be92e199c6a9cc9de6ef1c321e2edcfca1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb92125707fa175d7f4cc0b96488a848308e75887a1311b087f3b464ffb098caee6eeecb8730d58f12;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he0366f2c806f3797eb0d798cfc8b5ae05860628ab8519af1f147c951b997f3a6f352cf56fef762159;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48618897b77313594dc623792c8cedcba8ddeeff974c4c637d93cb9df449b07dca8e069ae7c360d00;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd13689a5936fb96a98a207cbb5b1ad2507e373f976ccf5daf0945dd22614d3c2cd1b020a4dd12658f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1c39c640aa30865d4407f7c81acd91b6a724d85c5e870db308d2e5d6dd90eeba18390264ef6580229;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h149f75b42092d834b32a4b761560a36c7f152449986c1367ee8ebbf9cbd9d97236cbad834a7a141b9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hde0f7afb5c55b36678920b006797dcce79bae603edbba1fd685c9290eba1a8b95db635ad7bd55cce7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf47749758cf9c0396160aa6025bfbc41ab373704c6abfa752a6bca5fcc19458eae8aa2aee6288bb77;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7a6fbdba01b09867d0e34464bcaeb0f822eb2b9e5e5a230d895cf1a4a8dfd0c0a69307fea35910c8e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb19c7198443592a36c5d7aecfae6a835cb43eaaca1be6576f6681752468a219bee6d2798844306ebb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heb7c1a2fea425d1baa2a0e1f6aed0c90f62abb5e89d4669ad6ef6444533c06eb5a927bbf71d35a469;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcf50ad586451c573838abc2b87e663c448dbf1863c8792ce85108cb1075a94a81ac5b6d9668751304;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3bb245b7f1377f6c636be86850479437ce6da6283ec66e60acdd3fac3482e5237cc1dfb8d21ddb670;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h361fe0f59da745f58f6d5b10b321d3064d7e1078e42f4d1d660e845e0a7a36188cf4570c0d94a47cc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17e3449822ce73ffc0b7181a652edfa8d42a061c54e4166ab58d130dd19a80f308f26c98f3acb29ed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd51a89a50f729744ee62eeaf5c60a7bc68a97c9b74b0933f4bfb3f80b5ed27cb849053dab60a9f6c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2a343f3bb50b98d2c01318aec5d71be9c7ef54cdbbd68965f3b222fa94d6ce974c33fa71c89471af7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h82b789130c405dd6e5777163eeb2b3eab476521b091f7a0d9cf716df0b789a34a9c9b031648c3d220;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he112358ef49830dba1012b9f324bfad2f94668b3d97075eb8af0bddb4c9bcf841b47ceba2e2e7982e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h63efcb4e113d6d3ec9722441e819712f8a1b2af54d7011f3fa85dbb69ca65fc78482f9841c910dbe3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h74a02923b4a54d6063b23f404d59a96a42a825c27b1bcb65d5effb7fb2dc41ec8cb5944f086f83bdf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50d6b5b802b74a23b16692ba5d99dbc38b0738c0a7a107b3cb7ee151d71918abbec4d9dd801deebd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd9f61813df688f54b0dd10dbe18bd3329a5be312c7b0a65671354881eb1755293855177f0ec1dc2d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf63bab45f064c98e7bc6b4910d385e3abe8930c81e1be2d0367292519bf7e26e9e75824b4c28eb259;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9be4b4498846c571356032d007a11d5dfa1b683f13bc0244a73b01f4c4ee43facf22654a78a40fb1c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfdbbb5fb03e0649863c6b4102940ccdc85418f92ffea03cb38b8bf09aef4309f2e4e50362473603ef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h641582892b993fe9ee15256c39c509c95d66bcda12a6c8626285eded226b9fc7a3f9a686a384f2af0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17c7b8069867b7b8fd1d8bb7af7c5c9a022c2a4b09b68d65ae5449199b91819e2bfb5d70035894643;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48ffc252726988e74a9c7e8b0a73839b159cd397d8b970e14be3eecdfb07026ee23d1f5aafb26745a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h50bcc5569f7912ac90487b96c97847c9e48f5d427dd0c020288533b24156cbe91007fa0779685597d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbd27b358d56db3b4acae9a15a00fc6f03bfb234451d45ab8e8a196b68be8eda882b1d9ec1f7166d8d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1858bb4975236e22d6d0de8ceafee21486563a63f55c1a76cb441c1805f078d55f2c7595ccfc3be6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4352281a7aeea0628bc9d1db52e08f1b2fedc502657c7bc695755eea41b41fab7d72702c6b699ba00;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hec50b1ca3d7cafd36eefe4f417b7571c0f57debf5c3611e13f71f5eb8a9e8cbf9e434f6ba8e1bde81;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5e24c85c86798052a40aa12f3d6b7be821ed4f962a10967814952fe17be8ef5e50d1841392fa94a35;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h559c2daab245d8d12cf01eee63c63c4ba2f145256f06f0eea8e06d1753f1a812fedfc825ed1935a53;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8653d14de0083b4619811191a0881f80ce66fc5dad829b133dd01eb498d653870d336c050c5874d2c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2463c4bc1686cb7fd112a34317b0211a2bdac6ff324c782a92c87c31349ff2828fa666e9d39c765b2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h240b4c69a14de415bc6d449c0d3bf0c237e1efc9e3b420317c07daab2782d76fdd04baa394632385a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2288009ba6067688328291093587e28646e847dc94cf0fd9847e1f3addfecaac914592c2d4d9c3704;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hedde442432c38605ac3a130e1f028153912adf070a304502fb83f2f794bf619e363510f79170d1fa9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h606bd4586677e758e04e6f623b7933978598679e93547d1d2fdea463c7c5d790586c17820b52c5234;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he2374431ee9fb4bfdc7b3fe6f2d21369da87c4e2a17b00547f42106744f88b7b9ffed92fa256609b3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcfa049f6359528b9e8ed8c7acc34a4680b6e792cbda84c9dc15f645c76bcf6e0a3a6967ddbb0c4e20;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a2c235ee2d1222574764a8dd95947d22801a589b0e7e6249af5fc258c6a001dcaaea476e9dc76c93;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3248b560060efebae4311b77417cc02b72ce5f3fe0d43d14adccdf41bd777d32967c5805f8a779169;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb9a2fbc3c496d79ef33481005166caadb9e1a78a5e678d3d79ed5fdc89a429c609174c2d64d49426a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h31345b4c7385ad829241e13e70cabb8a7a6e96417f72ad0c3cb93e0aafdbcb4ea0ad3db8f85394efc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5f06979b6d6d3930475331a2d9e06f61b10dee549f3ad1676538717d3d55001c4b9c7bcc4f73caec5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h24cbb4500ef7d6dc809cb4fea03530135ee113c64700f8c3a82f0f6c7a9dfd144c23d9a46db018fd2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haa57da610bf1467b7a9832a2c700a46bc166ae1465af73659341a3ec0ade1bd5b58b8b08fd5573020;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f1e26e1ae399f4371d1aa8e5e277cd9a8f6dbd1cbddc207017ec04009c7d92e586a6156d16800eec;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha659efe4b2b03045dd9f5b6a7b4897e62c12a0d8bc56fb6403059c0759e7f761036713a271800925a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1474aa18d4d405279e495dd0b4a41dddcec9decdd5b31b6655ca3d0ee1c0ba0ae157ada478ab7587;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc67ed8b4d2f3cdcdd6711cc0d94534062e0f7de2882123afd71aa5e3638b3cd571f48c7f8f82a5634;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h66fd86299e20c03661cc3e466b6cc0e80d078aaa31749c7c9f1809eb5a71c7be2b6cf01823c86e83c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7c8ad58a8cf1317413b7a1af520f10dab60ebf8c161b3d2fec1ee4cf822ec3e96cf2f1b390201668;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22cdcbcf59d19b3e6a72bccc324a3a42a6d2126e4c5b84167e27acd78ec5c3a503b28f375db2c5878;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h20b5543ba879b8837a5b15748a39438a2b1c831e76d25d475bee8d30dfe41fadc262012ce8979d3af;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4de6faa9f4185d1266897777bc355527619d63e65dec398241dd6a6432d02c26ca02686ce98ffac65;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7887f051a4315d4ff32df57d907684f98968fe03707c98b45d03ccbef0f5e3ef9a2259c5b672f041d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h728c7799864dbdd700f54e70918ee8ef4623d8e9bb84288f6048029aaff3796fe9266afd7880fd551;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7ce60c0142d28527cd22f9fa5923d925860cfe7685814f7a525e6feff3c26e5fbbe7050f5c22b622a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h99fc330f7608dc6b4de148c83679e37e7ad888a87019ed9e0ba5f9806b167875d813a51edfe40d6a2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8854e8c98e1f80807c70c8da8900959273276d04deb69cbcdf26e198373f6b94dad495f3a8ee5d605;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39d27d1fb46a74e9efb9a1d87f67db4418f938146c7a349ac7035d29367d7925f3b971fb1260a240;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h669f3042672b5e129c71174d41ffe89be0cc59787b5ede5228e19243558284b33fa9419ac3b2da98a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4df1f4deb00dd62c755620325c5dc0221fc4ae603d96e40e7782719cfc226df69f309db81da8db584;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h597a082e4996dca58c8b33d39a27e6a01f23d02c52f020d85786e0627b694f5a0de5efb93c419783a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59a37dd429191c1e3462f03b91021e174926d5d48ef4378c7aabebaec598d011fc08d92328b7df294;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3616b29805e2695382e6cea4e8a942b8e4abdaaaacdeec2717bdbc9ee056b5d1bfb6d119415176d9d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb04384db9a6600042199f96fdea24c8dbc4d8650839251679c3ec56a5c6f2ae20c97859313a529452;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he1f7bc0793e673d169194800033dc0aff2c5a2ce2fff278523a4ba4855ff8aadf0cf4de2d5d6f8f44;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he690bf37efc70a38db6549a3bf59ffcc855d48274abca72058a7a25b5841699f3b3ddc257c02d31a7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h735c38542b2a14e40edf22ba3148c7e7456fec54279476ff4510385914fa4e37f693762f4a8a38939;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2606e3954497207bad46049e00cc94e6863a1b479608e9634423f51e566d6d56525a6a1f6146d0a3a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc147c99ae54a4898555ca60bcc3d83662b2a24a123e89a00504357f36eaa989533070cb01b48e177;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hea2f91fbd8a9421a71526f370806b9ab9d8585fa1ee352d780773b1f4ee3955f91692c0dbd624569;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hecfc3851b37778b34b243c33c65ad6c43236c55b4d07266bac0d782a10d46cae4ba041c640f7616aa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5804e25987f87a07d6968153e347f0e9460f8085bcb90322eb6ac5d9b051ccea7ea0ec9697631ad5a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1dbfdf7ad7fbc211774c712ed5d5a796f2b11dafbd8a3ddb08f309c315552be00c67364f2bb4393a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc33f9e9f619236a071ba11998b73c5e68a73b36011513571861d3f9f7649e0f9b85c315c1c134e128;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9b2e8942faef443c80f22455f80ab0172aa5c1ed4fcf91f992458f5516354e7adc7cc01dbaea714a3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h363b3c1ea28abd82529db7ec70b936efc0d4613f4657963a9b4bf9123520066e317c8c43da6934b21;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hebc273a970bf38a522182a3fea900032b2a0e1507166f7a45b9925b52ef550830599b8f6ee17c614c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30932b6ca25b461b996d2cbe580ffa2610a7182c0c94391756efc89453feb05d7df21f89b42fa6ebf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5188ea2c75cd93f2a43a39a0524a511db52158e60dc09ab38481c307df4d78d83759a7463892a19c2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5463e31779e562d7ccd5d5f7e11d1c17205199f221182b3157fc92712a52489e322d35f90ca0f10a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h57fc5e3411df1bd0109bd128ad2b12c70b9607c68139dad07eadb6fbe31c6432b98baad0bdbe55523;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha61ba1fea26cd486227ac3b0cf3ac3994084b78f694f6c5260610fbf914d022417b93df6c4ac54fbb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hce9e15da78e97f142184339a5edc5e438e370ad9d3414b6879b77c801cad1c37297d0b97952b24748;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd7a0efdeb4b26c3e0f0eee37ca1f45296c4cfff5a3b20559e0d0b5bbf76182d69e998d27f9458ba47;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he7e8e0b2f95046de42cac185fec820437e373aaa1717050e5b4788db5169a824523232c77770f7a85;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h580f4ba75280b0d984710bbba5c07e3dd0c500365e077bff3d88f21c9af9fab55328d578cd84b3332;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h94979d067d737ac0c2b1788f7b74cfc34ce15b3f05c715f5d405dba04aa3aa3b4d552e4cb9a8dcd64;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4dbe47c60727e1f8bb6280e76b323a4ef7379d0c6d85b33dde3571901bdca3493376ebcef77eeb2ae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb157d4d298a72aba5c21ce7e9ee3e0c4690faf175cd929dda3eb6d3b1d3d7052f25fece906e79068a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h76cc5e95bda57f91d0d1b4e677fee9d03550b34d92098237e04520c995dbf88e64823435d6e9d0e53;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7d280de713bfbfe65b1df88f835b768c274b12265cb80853e523f78ea4b77a806572a68f4314e954c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4d3cd0d346dd7f03f6f22df72db0a02f3f9f43e2b3641ce0d5886a7ebe46d9fc12733e6273b61aac0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3b414c213b5ada23ce0aabd7a9b3b0ba45048ce17b9948f1e02e7fce06124cf83d33705bf28f45c98;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9c06ddb8811c21590338fa77e74b73f20224c5eedc5158c80ecfae317531c3b515fd163e4498aa726;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcc21d22e08418d9cf8a043d5ba2cffc2e55045b96328a162d84234711f6404ce042c357fe2ca3106b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa55aa7bbb34e896565e51f6a8338f6ceb67713cb24881830df670d67f51af9d69e6e2181d4fd617d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ab586edc2e85edd1fec67d0d245d9aa1f49d5801dc0b424444ac02b839a698ddff6e2f3226bfc75b;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6928970b1d711daf3c307bcb2f7a1a608b31864c6918ef4fd5dceb4aff931d0b16eaee555c789b385;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc60de292ed2e4018184568b6393560d237cf1298995b8a59871a97ee33ff5b1bd21237c5c1a189239;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha9aec476bd29f760ee872b581d2cbb535e26e6a4c20f776d67d8c812d9f66a674425c28ad59dcdaea;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha7faf902753349da61c9d335a87d3d9d3c87aef9dd109b3d1b0987fd23fb5ad9553b28d5a56e9501d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h327191b53839d8668518a0bb8e1dd1a10be45721f6d83c3b636f0da71743a789d3ccf0df3a0241ac6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5bff3ecf75bb11adee2668e2e6497d528acdb8c5e89e9c86262db2280a394178b247a87683c8c3fb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc2a05aab9417e61c682d041e00a21d42b6e4a660c19d5aa0571f2f46919d7f4651324a5ce3b18b326;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13c5704e1ca330366da0e690076de1ced0cb75ae61509669d6fa26cf393e22c3f0c2e652a7843048;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1582693b5010c527d768b7770f0644f3747ad7a251bcd32d269a25bf2e669efdae4a0e8846440f1f4;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h13baa6dfa85f403e4916e4fca724c899067cdd1535b16ac923d26d37257454764ed75c4f93accad0e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h370a595ae586803532ba8e590ff4e1ce46b937d91198319e4208956cbd4f6e470fc984dc6b5d6c0aa;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdfa051f7a2bdcb3896a0aacc49d4be3264dce9d4ac6247a593d5c3304317a72befdf9193944cacc9f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h558151ce6a8fdfd715bf1d29110281b9a3623e0bec4e3cddb7d59ebbbb3cf87a27880dba7381e2866;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h11a068a43e8655bd1c9f15b3ea834eb9dd4c1b4047753fd8e106edcf8d04b0f6253c88b60e08f933f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h47029dceba07b1d0263bfcaccbeb479d02e01a5c68963d3c8ffa63db866b875f365deae549baed6df;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5aa02e7bb5650d250bbf7c4c4fc760e0dd324f9cd97b3ef67b2dfe37884d28a85b55e76aedf4ec331;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f74c34b21e85bdab27ffc6ecf89a3f024b84067e8e0ba953d7e760dea0e18f11f41eac1a7d096cfc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd51d8f703eb4f976412d1a7de5593c3116beace94bc6b2d57901b3e06ac4bbd2221089239dfab7f64;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha3185991f6e772b8aa07f1fc671ffbb176c695bca971509427e655cf35a4931fece7ec82a86c52aed;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha92af3445d7264aa0903c7b0168fa658f3af83c0f57f060e7cd43b9f0deb9767c872da3d70b16ee61;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72b7a8709cdf5537073ad456695938f0471936b33f70ee46393704a33950ef17905b023868d35e46;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he69abd0e30f98aee248029e8cbaa5fd0424a394ab99b89e97397da728a77534cbf217de6dda34e805;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he6a14ed02c81fa50ad319d93e1d45572caf3e9eef1301e212dd388052eff3cf7ad1151feedf8c2911;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h553fa583b3aece95bb1604335b629d351beb3e2393e068c76a7818c530eddc185c27b11927d39510;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he839d44357bb92e96baaf2f950984b7c164e7df805d751c4872fbbc508a8bfdaa1a5e11a50005b2e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbf1f69b056a7db4f174a7e45ace23e0568b376c8ee3481cb8824c5e1947c07bcf81259ac03857d169;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9dc97517264c149fca5ffe8604780a07f5b4a39667a09c2bdba103be95df04a8aa3a3730ec7fdd209;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h345b258578ea3d77b24e3a986504513d200122b76e0b9612966c426912e55f68a71eb1e51a2816c58;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3011bddea97f1b5b1622515dce9b9973146662c52083c1337d326184c2461ad87b7254f0bd9458ce0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6f3e07b9ad1cffff9936b5588db68d61730249f042422f1971a514b64adda71669cd86099a7b3af6e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3c74e9e3600394d90f3a566fd306ee5c41f27f9645cfb420cc831f1414fe1b687089bedaa14df64c5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h69c593f0dbce6967313ef221d480a12479ed6ed319b5e62ca65d57f4469757ef945e25225142be7b2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4f594567a67c04a785c47c13e0c08cfa773768a90d4cf046845c2b7ae307c2e9afb66f7726c789093;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h44daffb25abc5487258723525617c43b239567cb32f3a1c7d154748f102c956b54d2f73fe87c6b23d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf004f9ec5521ac0c56038163db9b9f96fae9d2da3d82dd87c6a71195e4717712f792f1d3cc77d85dd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd4b176726e0e8ab11f83923ff5fe0d315022fd3a5aff2e8785ab411e1153f464cd868447700ec5088;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha81d13d1d004d0a2c37a6ec600233777723022ffb4322a41a588e9a9f874d29d206dbf81a5ac2b5d8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf001d7795878c61e473d08cf305fc89ca0437681a02e3cab8a815b9ee6b53d7fa3b42794f67793159;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5b3ef2785de9352048ebcb481507e606fbeabb4b74d500ee2a72d79c3f14e175798fe8b065c9aa768;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1121b24adb855e1b30db6784758c7c623d37d6d5f20526667fe59f96b3697cf612fc9debf47e25576;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3f8ecaad819a7dcd0022d23f52b737239ea99f1a4f1aa70f43137e6000b36a8e1ab2764b2b3290dba;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9ecf8424c9a3e54447b1ae83561a2832c3da31f16bee247fc84d216955eb48f7715a26464d307bfba;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'had30ee184fcfb6eca390b255bddfcb573a1a8bce1853be7efcaf2309a84917fe489abd6a52db1d5d7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he99ae744ad7d7d1076af9c0fa332b8ead35a26cb85bd314ca4c74383beacadb0402b263d8127dc849;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6a5ff3e819d7bee6866af6a6db64a8e026b3b9cc2c58b1c2486665f6f410447e4d9ea9d31c243a1a1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9f6b10f0be2957c6fa8e856b0defe9efb776a78beaa38d5cbba2d584f4fb1438491aa1156e54ed8d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdb892077aa1645b4c955319451d9326f6f9d664f54a6edd29fcd87b6f31fd51058b639628ca489258;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd547b102445f0da23cc816f94935ce0a764179022f394e607346c1a938b99771217ea244e7f173cc0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8e600310828f8eb1f6187cb8ccad5a979bee4140965d1b670e9db9f1b72a63c55fea353302071dae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h135993103064ef1b48c9b08c025f59a19793c2bed023984198fcef08b337f2cdbfd101dc2d5b75631;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd8d73918efa988cb47ad119a51babdae6c947498fb58d27329b0cf5e40949fb510e671946129b8d46;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb33062e86c0af49bc3ee5856d0ad09a1f0794d35a14f9afbccca926162def206523befb9af1fa43a2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h855e262b00c2148991427ed3a7df5cbf45a7f8afc92987fb329837196dc3d92ae9aa390bb75b2da19;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h81dfaba8cdebdb50968e8ae8906db9656147651a1558cc3a12115a2aa6995577af4df310ea2775bcc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h72e9fc7509496da80b94db77762ca8976509f051d055432d32386cdff671bc9b937e77e2f3ec12d29;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hac3c661f2d6b94f38af3372dd3e46a8da07126bbe74ead8292ea9d29f66495e290a4415968ca90922;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8951d5931e82944d09c7c0259e52e26886d294bcd3682cea2c8fa3167c841099c2f582473874b46b7;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc614069e958241a151de8ca27dfbc047b13e4a8c6ad1397898033fd7814a87dc31560478094a51cbc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha8b50baf0055c0cd6bcf20abe87a32964395b555354fafc89ed49e0136bd3183a0b67434140ee1b98;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f6529753d032ab9078cd458962170c1f95cb234aaa389c686d3b394a4e3b640efd5715f12571030e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h18dbba2b0383b57d2b16d2046d63b90f66120cce0f1351dad49126aa3a98b98590734d746ccdb5fcd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfe2ade8127196e089b739c84e5ad3cbb977726f7e0b4ddf24cca221905bcaba3ecdfa46636d4971a9;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h642cc4aa424c7badb51acb74a7f5048b5ae32b8929b2f5f6f837012c5688ff7796f7f83a209f99e2f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'heabcf4c2208614cbfbab40384b7f673267e3e029ee72a6639d24e7cd37d68769042edbacfdd82d398;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h34f6d2545ceff6d2889cf1491076096df9b14d280c62d805a4c5ef7adfea5c44cb8f29326798d814e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb95831050eb717193fe4b1ace4ad365a661fe9143a9cf5f7c4e0c4885ad727f66fef8fd0acfaa40eb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hebc2ae9ade0f908a4af4302859fdf29bcaa51e0d679a4ecb7048d46b655f0c411d3e78a66a909bc46;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h52c0cc2a7c245786301f3f184c8303ca2c8d0cfe23521da4f1dc7450c2587726fce7ae0e90c0c0f72;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h30e43f2a5156a16cf3cb01d1c67519e6c89488e620328d70b094e974e47e28c7ba54e1540a73c8936;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h820e1256382381da2e6ca639d688925f08b23c6c698f6f2f460302bb64c14b019ab3eb3fbeaa98b67;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29062958f7c3606aa42a77cf00bc43b4e634a57267ae3929e4576ec8c9473152ba4bcb702b330e63c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9d9387f4298e84eaaf00cd96b5866051e876d257bcbb900fb8b763b7f7528edfd7590fe6709fe865e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5693495854bef7aaa5a642e10e65ac100226b245f4e43e33b04df07cbc7999901f3fbc3f97c741869;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h3a98b80f779b09ee7daa28dcf6e588594f8ce925b49850890398db0680ce96193980e771ba0be43e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d75adfde672ee1a19a91525cc80303c0a04243902ccd07c891cbe0fcea2e4189a09bf1d7fb0b9cbb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha4f005767333d6190bff40ccececb7a51d220735fce2e8b1dc324eb80402a31ae3e028cad57fa2ac0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hecb097d667e52d76065a326ddfc2a3cf5ba761ff098cb8c3edafd0ffb994308999e820de0e92bda93;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h9f12c55ef2e3756ae810f44a2ae9b0d0e973f62ac3d49a7a2a6130f5a9323167879dc173db5170a99;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h29f021e4c900497b5d64a4fec2cd7a3153ab9643bb70945570ec75c61c5a0fed5021749601f2d3d64;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdcf4c2015d6b60b4b1ed114fec3e356ce3db069d319890f8f30378efb7af41e22c271f72ae2bda4ac;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4936e8c8a1ded341712a74398ad92cd1f0c8cbd1f1c705216f2ab5a12b1938c931bf3050296a89917;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hbb62e75766a7521c6167f2e1c252520fcca3393b613a88f60b0e191237faede9faae8c262a790a10c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb638922af7806a025e74e1d3154cb1fcffcb74ab3f63b6305f2992066236c5bac58d9642a576e9a19;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4fc32ae4f4d1d54a6976757f6ddb5d3a224abd67b99345a274678e58146aa66c3e38d89441ce4e630;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd618ba23f148712cb2a44262549f3e5dd71eb177de6dcdb8dd2341f2ca74a51a959807d58a51934f0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h454351a96aa4374dd1c87481b6a81707b45d9afd71b6135f0b100a13d73ff5e385670f923b949e455;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h7280d4fd76d43362d944a2def5220eace2ee799c1e5923ddefac25d82ecd4d3f66440f9b12946cb6f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'habbd53b03fb4e43a3167cff21177aade96892ae02dc84cb777a7696e5bd335a1465cb521e9e755abf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he24b02f7e9c92dcc92fa40e7e61a69edecdcf4609c7f49d3d4167541fc25f8254adf8bd9611b9cebb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h949eacbc8554042c1ecadd0c445e2c9733ebed89a5e3e0d8176048839154ddb0fe1b00e87350ac844;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h22a71442f7c7f03d9b6d6bd844e722ddcb60490a00032639e6f88c8762f0df2fd630f948b44c10b3f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h135f52227dcd243c856a2d62d1a7707f3c65f88073d913f0f557b32cf92dd4842e8f8d174e1a5fb6e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2f4e2a160eb9cb67c1e8a9a23e8c458f1d219904df51ec8b90f03c5e61cb94cb1933ea68ac909030;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h5022322bc2343a5172bc4ed51e8225f07c62187020e7b4cbf689183fabceaa61c696d7b5ebac5607;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd9e44fd98501bf86cb669fe5cd3f578e1a6383f02e961009b8b8761527f3cf5ac2317ba51e5ee3fb3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he9c7a84ad54246adf3a39d63ee1e7cf51fea781cf951c533fbadcf3fac25e0284d9e1a86b0c7f7428;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8d52d6b6c6855bfc994f4fe4cd7a4488c30085c19ec0ba6069cfb43a0314f37fca6994371c7f5f4fd;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf9992c4c0a77798011a16cb3479809cf64a3f8e1e0ac608e02012fed7ebd6f0edcf1b32b54b5a31b6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd804cfa3e90244421bfcd39c08bf6f7a6c2597ddd3ae52ef880337848558f3a1feaf2aecf10c5c2d8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd66f071f80da11f659a1703c3b3a03fa8e56e44c5e2cd99cee5af6c0400c2bc7f1440d4375fbe1c5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h664c4e908cac1991bd4ee7ff6eb34d44ade46dc17fe0d55c6082ff4fb1b82973a01127c0e2cb86e83;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h56b7850bfb6f8b2f7cbcf7a36abff05594c0003b5d2de0942dadee87a353ceaf90557fb4718f7be1a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h68733e825c22498045c1b7a91ae448b60bef97c0e49c0ed58b784f60f25ef42911f65fd323a8bb8e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc47d05bc2ec3ed29bc562db10eb6dce871a16174b89d326db8cc7f01166964c8606bbf5528b0c875c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc5b1196898fa675f38558dc644945eba8a96e33ff90bd53d30bbe5802c9c822a0fb0b45200cd8aebf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2859f2bf497d25243c05b6a47399c0bb9925e5e1a53c2171a671903159f091a6b7d1a1f11c108200a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd0dfd2f7684b93aa1b89610d6f3388414cb3ab4d909ca0690d4fb3b12cad283b139a59419d6390a4c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h17c8abeabc3b807b597580d11f3f1984f5aeb0261482a72538188f477960d35a04f9a649cffafd12e;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h1ac386e600a6388f9c93f670a66a2eeeacdc0f677120fcd297183c3e4f19e290ac61d51ba1b061185;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h2018122787a52e61a89c09ffbd8b906500d608e03c13824f6db21cb60f759e06a81e15f08a28dea6;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h52ebf7765fca7050f4013372e40642d04717ebbb4dda4b6d210373281073f08846ca53321d2c170b2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8bb3294c70c95606b9da4573fee0f64096dc4940e3cbda335236097cbf14f55ef0944aaa5f6f96914;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h817865980e516b9704574f2a75e1744bba39e2ad6a54e53185b3f843f06bef36ec8166f330ee7bc0a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h584376e730794819aec26661b791bda7a875264cc88a19c7cd2a664f5168671922bb8663fadf2fe75;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hd900264c591e2066d664f83e86493253174d7e047a5a332ac8c14cf411354a981ad70c57149234f51;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d48c7c2eb872840360d71d563f37f99c5c78ffb2889b548d14bbdf99b222787de342b946ef024f5c;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdc53db470ed8278547d6d20dc4bd544bb6cfb452c3c11b226ecd6a7caec2c3d21dccd067fcbf59f41;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb3946eff6bfe90154d73b6c139ad862be8769241704b96b3e7832df38eda8757e2c60e0dd8428bfe5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h8e3fa512c24fc602ffefacdde25d52ae8e2488594b768ef5d17ec67169c41993300b69a74aef31cae;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h39faf350784b0b4a3b8e409c52f781e9cb0488ae799edd297720c6c235d5e8ab7ba7f5e1456ba6c88;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hfa0980f9e772a16a9b46b021c1421cc89ad8857df89174062cbf5ed7628bdd9687e5fcb29593694f2;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc9d45d36b774703f5c6e0f5077aa8426a238bc9c34b0ff2fc7fecb1dfd9b36d11a6c1344f2a95fdbb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h36a4db48059b28d07b32c5b4e74f643d9b8614a119aa9630e461decfa9132dcb52066472ae64762f8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h23a71df7e15135cbecb871ab853ef2d2fc2cefbcb44d1f0cdbd1ff3d99d90feefc18c8d0cbd4879f3;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdd4722f2f141672ced9d5a06c86fc9665f40300062e4c689564917334e0412fd838c9785999782ef;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h59b842a0a86b4631001e5541fd6846ae7d4965a3e6896c3aab03e2527f483fb26f9a9628668fe6feb;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4c73af8cce9c2d730078725760ef2959cfe45b9f18dee3adb26e9c746c05505ceb2ee122534d82651;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he73bdef3d323fbfd5d2bc30d9ae890dbfa510267bc5c42fb1763971ee971564e5784f9523e88b6782;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf63a5b8c0b96e6050f940912d0e55597b916dd584a69c7b4b9d8f4d608b30a25f9afa64b784ba6e08;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h79956e7b58c706279e04bfc14061aa77cc5c1ebcccac5ed5520feef9bcda440f67567a8560377d30d;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hb5bf911ae96f384e0a56bdc2c1f318a713eca9afe2c19e7d6e99713fc8150d25461e461d50bf172a0;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hdefee018a5507218e85274aae8e277e1ad845977a211da4ca2aa8e11d8ff0ad8f585fb32ea02610e5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h69db283b9541fe4f26219a4e5bbec67bf21927145c46182d2d1ea0f142ea2e6ea2a85d4c1aa6d2e85;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h226d8d42b40df431f234aee222185783b45466195611c54fd6efecbab3f67a7be473e97ac5c593c83;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'he5191eed2e13610008d991173e94ce5949fe34c1b0e129d1067e076a698d2e6d3bf01650bc3fe81f8;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h48148ea3c0dd14d9b778099f06f6e7b95e9d5f6771acf2a575dab3e7919aa2ca78a7e8f0529de472f;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6e03bcbfcb73d53c57b0a9df992784885fd3b1b3e9c2c747ca3ee19b9df9852c7d9f3f54951019311;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'haaacd2381ec89c0cddcb60ace3aea88bee665b542db5dc55cf8e8a5aa7be2d3055240dcce1a39c52a;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h75b11262c8b2009c89c4da4f3497f1ee2591cfb6a7ec5dd7ca8553c9b5d4e21cf32d63a4e1f0a0dd5;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hcfeffea2cf17d224958013e758c1d8fdba72b6bc474c0978da53db5a98b935c3c7580e91ea5065483;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hf606f0b3a44fa693952b7c5713d388e43aca3b9cfdce6b19b85425efad5e01cdb6a27643425626f92;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'ha493d841fea93acbc0a2704bc8c5595d39ae86f6a9c37a28e84ef66525e958598af7d6041e531b3bc;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hefdf9ca750ce3260c43696c9711833d953aed3a0a32b4c680ad42e7547986d7a162d4281b44e0a7e1;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'hc672cd2776383ac36e88658ba2f5e8f19f613875368647345c7cafb5fc3bbbd35c748e82de2086b33;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h6d6e1a3b9ed07e73e23d0063ce86d6674c0cf41b4f8c92acc41b6f1b71152269ef4af75d161a095cf;
        #1
        {src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 324'h4405e677874f2542ecfd595b407b2fd0d529c982602947d827715e7295920b8b672caad6fdafbec2b;
        #1
        $finish();
    end
endmodule
