module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38);
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    reg [127:0] src12;
    reg [127:0] src13;
    reg [127:0] src14;
    reg [127:0] src15;
    reg [127:0] src16;
    reg [127:0] src17;
    reg [127:0] src18;
    reg [127:0] src19;
    reg [127:0] src20;
    reg [127:0] src21;
    reg [127:0] src22;
    reg [127:0] src23;
    reg [127:0] src24;
    reg [127:0] src25;
    reg [127:0] src26;
    reg [127:0] src27;
    reg [127:0] src28;
    reg [127:0] src29;
    reg [127:0] src30;
    reg [127:0] src31;
    compressor_CLA128_32 compressor_CLA128_32(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38));
    initial begin
        src0 <= 128'h0;
        src1 <= 128'h0;
        src2 <= 128'h0;
        src3 <= 128'h0;
        src4 <= 128'h0;
        src5 <= 128'h0;
        src6 <= 128'h0;
        src7 <= 128'h0;
        src8 <= 128'h0;
        src9 <= 128'h0;
        src10 <= 128'h0;
        src11 <= 128'h0;
        src12 <= 128'h0;
        src13 <= 128'h0;
        src14 <= 128'h0;
        src15 <= 128'h0;
        src16 <= 128'h0;
        src17 <= 128'h0;
        src18 <= 128'h0;
        src19 <= 128'h0;
        src20 <= 128'h0;
        src21 <= 128'h0;
        src22 <= 128'h0;
        src23 <= 128'h0;
        src24 <= 128'h0;
        src25 <= 128'h0;
        src26 <= 128'h0;
        src27 <= 128'h0;
        src28 <= 128'h0;
        src29 <= 128'h0;
        src30 <= 128'h0;
        src31 <= 128'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
    end
endmodule
module compressor_CLA128_32(
    input [127:0]src0,
    input [127:0]src1,
    input [127:0]src2,
    input [127:0]src3,
    input [127:0]src4,
    input [127:0]src5,
    input [127:0]src6,
    input [127:0]src7,
    input [127:0]src8,
    input [127:0]src9,
    input [127:0]src10,
    input [127:0]src11,
    input [127:0]src12,
    input [127:0]src13,
    input [127:0]src14,
    input [127:0]src15,
    input [127:0]src16,
    input [127:0]src17,
    input [127:0]src18,
    input [127:0]src19,
    input [127:0]src20,
    input [127:0]src21,
    input [127:0]src22,
    input [127:0]src23,
    input [127:0]src24,
    input [127:0]src25,
    input [127:0]src26,
    input [127:0]src27,
    input [127:0]src28,
    input [127:0]src29,
    input [127:0]src30,
    input [127:0]src31,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [0:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [0:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38)
    );
    LookAheadCarryUnit64 LCU64(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out38[1], comp_out37[1], 1'h0, comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], 1'h0, comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [127:0] src0,
      input wire [127:0] src1,
      input wire [127:0] src2,
      input wire [127:0] src3,
      input wire [127:0] src4,
      input wire [127:0] src5,
      input wire [127:0] src6,
      input wire [127:0] src7,
      input wire [127:0] src8,
      input wire [127:0] src9,
      input wire [127:0] src10,
      input wire [127:0] src11,
      input wire [127:0] src12,
      input wire [127:0] src13,
      input wire [127:0] src14,
      input wire [127:0] src15,
      input wire [127:0] src16,
      input wire [127:0] src17,
      input wire [127:0] src18,
      input wire [127:0] src19,
      input wire [127:0] src20,
      input wire [127:0] src21,
      input wire [127:0] src22,
      input wire [127:0] src23,
      input wire [127:0] src24,
      input wire [127:0] src25,
      input wire [127:0] src26,
      input wire [127:0] src27,
      input wire [127:0] src28,
      input wire [127:0] src29,
      input wire [127:0] src30,
      input wire [127:0] src31,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [0:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [0:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38);

   wire [127:0] stage0_0;
   wire [127:0] stage0_1;
   wire [127:0] stage0_2;
   wire [127:0] stage0_3;
   wire [127:0] stage0_4;
   wire [127:0] stage0_5;
   wire [127:0] stage0_6;
   wire [127:0] stage0_7;
   wire [127:0] stage0_8;
   wire [127:0] stage0_9;
   wire [127:0] stage0_10;
   wire [127:0] stage0_11;
   wire [127:0] stage0_12;
   wire [127:0] stage0_13;
   wire [127:0] stage0_14;
   wire [127:0] stage0_15;
   wire [127:0] stage0_16;
   wire [127:0] stage0_17;
   wire [127:0] stage0_18;
   wire [127:0] stage0_19;
   wire [127:0] stage0_20;
   wire [127:0] stage0_21;
   wire [127:0] stage0_22;
   wire [127:0] stage0_23;
   wire [127:0] stage0_24;
   wire [127:0] stage0_25;
   wire [127:0] stage0_26;
   wire [127:0] stage0_27;
   wire [127:0] stage0_28;
   wire [127:0] stage0_29;
   wire [127:0] stage0_30;
   wire [127:0] stage0_31;
   wire [35:0] stage1_0;
   wire [39:0] stage1_1;
   wire [57:0] stage1_2;
   wire [58:0] stage1_3;
   wire [66:0] stage1_4;
   wire [62:0] stage1_5;
   wire [49:0] stage1_6;
   wire [69:0] stage1_7;
   wire [55:0] stage1_8;
   wire [60:0] stage1_9;
   wire [53:0] stage1_10;
   wire [57:0] stage1_11;
   wire [57:0] stage1_12;
   wire [60:0] stage1_13;
   wire [45:0] stage1_14;
   wire [46:0] stage1_15;
   wire [86:0] stage1_16;
   wire [62:0] stage1_17;
   wire [65:0] stage1_18;
   wire [42:0] stage1_19;
   wire [65:0] stage1_20;
   wire [64:0] stage1_21;
   wire [60:0] stage1_22;
   wire [43:0] stage1_23;
   wire [89:0] stage1_24;
   wire [69:0] stage1_25;
   wire [68:0] stage1_26;
   wire [55:0] stage1_27;
   wire [55:0] stage1_28;
   wire [56:0] stage1_29;
   wire [60:0] stage1_30;
   wire [70:0] stage1_31;
   wire [33:0] stage1_32;
   wire [15:0] stage1_33;
   wire [35:0] stage2_0;
   wire [19:0] stage2_1;
   wire [26:0] stage2_2;
   wire [33:0] stage2_3;
   wire [25:0] stage2_4;
   wire [30:0] stage2_5;
   wire [47:0] stage2_6;
   wire [19:0] stage2_7;
   wire [38:0] stage2_8;
   wire [22:0] stage2_9;
   wire [21:0] stage2_10;
   wire [26:0] stage2_11;
   wire [20:0] stage2_12;
   wire [34:0] stage2_13;
   wire [26:0] stage2_14;
   wire [22:0] stage2_15;
   wire [22:0] stage2_16;
   wire [48:0] stage2_17;
   wire [37:0] stage2_18;
   wire [20:0] stage2_19;
   wire [55:0] stage2_20;
   wire [20:0] stage2_21;
   wire [26:0] stage2_22;
   wire [33:0] stage2_23;
   wire [32:0] stage2_24;
   wire [46:0] stage2_25;
   wire [36:0] stage2_26;
   wire [30:0] stage2_27;
   wire [35:0] stage2_28;
   wire [31:0] stage2_29;
   wire [18:0] stage2_30;
   wire [33:0] stage2_31;
   wire [28:0] stage2_32;
   wire [17:0] stage2_33;
   wire [5:0] stage2_34;
   wire [1:0] stage2_35;
   wire [6:0] stage3_0;
   wire [12:0] stage3_1;
   wire [7:0] stage3_2;
   wire [12:0] stage3_3;
   wire [17:0] stage3_4;
   wire [8:0] stage3_5;
   wire [33:0] stage3_6;
   wire [12:0] stage3_7;
   wire [16:0] stage3_8;
   wire [8:0] stage3_9;
   wire [12:0] stage3_10;
   wire [13:0] stage3_11;
   wire [18:0] stage3_12;
   wire [10:0] stage3_13;
   wire [21:0] stage3_14;
   wire [11:0] stage3_15;
   wire [12:0] stage3_16;
   wire [24:0] stage3_17;
   wire [13:0] stage3_18;
   wire [25:0] stage3_19;
   wire [15:0] stage3_20;
   wire [13:0] stage3_21;
   wire [15:0] stage3_22;
   wire [10:0] stage3_23;
   wire [18:0] stage3_24;
   wire [13:0] stage3_25;
   wire [18:0] stage3_26;
   wire [13:0] stage3_27;
   wire [10:0] stage3_28;
   wire [17:0] stage3_29;
   wire [14:0] stage3_30;
   wire [8:0] stage3_31;
   wire [14:0] stage3_32;
   wire [20:0] stage3_33;
   wire [8:0] stage3_34;
   wire [1:0] stage3_35;
   wire [0:0] stage3_36;
   wire [1:0] stage4_0;
   wire [7:0] stage4_1;
   wire [3:0] stage4_2;
   wire [6:0] stage4_3;
   wire [7:0] stage4_4;
   wire [8:0] stage4_5;
   wire [10:0] stage4_6;
   wire [10:0] stage4_7;
   wire [10:0] stage4_8;
   wire [5:0] stage4_9;
   wire [6:0] stage4_10;
   wire [3:0] stage4_11;
   wire [8:0] stage4_12;
   wire [6:0] stage4_13;
   wire [5:0] stage4_14;
   wire [8:0] stage4_15;
   wire [6:0] stage4_16;
   wire [6:0] stage4_17;
   wire [11:0] stage4_18;
   wire [7:0] stage4_19;
   wire [6:0] stage4_20;
   wire [9:0] stage4_21;
   wire [6:0] stage4_22;
   wire [7:0] stage4_23;
   wire [10:0] stage4_24;
   wire [5:0] stage4_25;
   wire [12:0] stage4_26;
   wire [5:0] stage4_27;
   wire [6:0] stage4_28;
   wire [5:0] stage4_29;
   wire [4:0] stage4_30;
   wire [5:0] stage4_31;
   wire [6:0] stage4_32;
   wire [12:0] stage4_33;
   wire [11:0] stage4_34;
   wire [2:0] stage4_35;
   wire [1:0] stage4_36;
   wire [1:0] stage5_0;
   wire [1:0] stage5_1;
   wire [1:0] stage5_2;
   wire [4:0] stage5_3;
   wire [2:0] stage5_4;
   wire [3:0] stage5_5;
   wire [3:0] stage5_6;
   wire [3:0] stage5_7;
   wire [7:0] stage5_8;
   wire [2:0] stage5_9;
   wire [2:0] stage5_10;
   wire [5:0] stage5_11;
   wire [2:0] stage5_12;
   wire [2:0] stage5_13;
   wire [1:0] stage5_14;
   wire [6:0] stage5_15;
   wire [2:0] stage5_16;
   wire [2:0] stage5_17;
   wire [3:0] stage5_18;
   wire [5:0] stage5_19;
   wire [2:0] stage5_20;
   wire [5:0] stage5_21;
   wire [2:0] stage5_22;
   wire [5:0] stage5_23;
   wire [4:0] stage5_24;
   wire [2:0] stage5_25;
   wire [3:0] stage5_26;
   wire [3:0] stage5_27;
   wire [3:0] stage5_28;
   wire [1:0] stage5_29;
   wire [6:0] stage5_30;
   wire [1:0] stage5_31;
   wire [2:0] stage5_32;
   wire [3:0] stage5_33;
   wire [3:0] stage5_34;
   wire [3:0] stage5_35;
   wire [2:0] stage5_36;
   wire [1:0] stage5_37;
   wire [0:0] stage5_38;
   wire [1:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [0:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [1:0] stage6_19;
   wire [1:0] stage6_20;
   wire [1:0] stage6_21;
   wire [1:0] stage6_22;
   wire [1:0] stage6_23;
   wire [1:0] stage6_24;
   wire [1:0] stage6_25;
   wire [1:0] stage6_26;
   wire [1:0] stage6_27;
   wire [1:0] stage6_28;
   wire [1:0] stage6_29;
   wire [1:0] stage6_30;
   wire [1:0] stage6_31;
   wire [1:0] stage6_32;
   wire [1:0] stage6_33;
   wire [1:0] stage6_34;
   wire [1:0] stage6_35;
   wire [0:0] stage6_36;
   wire [1:0] stage6_37;
   wire [1:0] stage6_38;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;
   assign dst20 = stage6_20;
   assign dst21 = stage6_21;
   assign dst22 = stage6_22;
   assign dst23 = stage6_23;
   assign dst24 = stage6_24;
   assign dst25 = stage6_25;
   assign dst26 = stage6_26;
   assign dst27 = stage6_27;
   assign dst28 = stage6_28;
   assign dst29 = stage6_29;
   assign dst30 = stage6_30;
   assign dst31 = stage6_31;
   assign dst32 = stage6_32;
   assign dst33 = stage6_33;
   assign dst34 = stage6_34;
   assign dst35 = stage6_35;
   assign dst36 = stage6_36;
   assign dst37 = stage6_37;
   assign dst38 = stage6_38;

   gpc1163_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2]},
      {stage0_1[0], stage0_1[1], stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5]},
      {stage0_2[0]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc1163_5 gpc1 (
      {stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_1[6], stage0_1[7], stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11]},
      {stage0_2[1]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[6], stage0_0[7], stage0_0[8]},
      {stage0_1[12], stage0_1[13], stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17]},
      {stage0_2[2]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1163_5 gpc3 (
      {stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_1[18], stage0_1[19], stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23]},
      {stage0_2[3]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc1163_5 gpc4 (
      {stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[24], stage0_1[25], stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29]},
      {stage0_2[4]},
      {stage0_3[4]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc1163_5 gpc5 (
      {stage0_0[15], stage0_0[16], stage0_0[17]},
      {stage0_1[30], stage0_1[31], stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35]},
      {stage0_2[5]},
      {stage0_3[5]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc1163_5 gpc6 (
      {stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_1[36], stage0_1[37], stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41]},
      {stage0_2[6]},
      {stage0_3[6]},
      {stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc1163_5 gpc7 (
      {stage0_0[21], stage0_0[22], stage0_0[23]},
      {stage0_1[42], stage0_1[43], stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47]},
      {stage0_2[7]},
      {stage0_3[7]},
      {stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc606_5 gpc8 (
      {stage0_0[24], stage0_0[25], stage0_0[26], stage0_0[27], stage0_0[28], stage0_0[29]},
      {stage0_2[8], stage0_2[9], stage0_2[10], stage0_2[11], stage0_2[12], stage0_2[13]},
      {stage1_4[8],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc606_5 gpc9 (
      {stage0_0[30], stage0_0[31], stage0_0[32], stage0_0[33], stage0_0[34], stage0_0[35]},
      {stage0_2[14], stage0_2[15], stage0_2[16], stage0_2[17], stage0_2[18], stage0_2[19]},
      {stage1_4[9],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc606_5 gpc10 (
      {stage0_0[36], stage0_0[37], stage0_0[38], stage0_0[39], stage0_0[40], stage0_0[41]},
      {stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25]},
      {stage1_4[10],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc606_5 gpc11 (
      {stage0_0[42], stage0_0[43], stage0_0[44], stage0_0[45], stage0_0[46], stage0_0[47]},
      {stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31]},
      {stage1_4[11],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc606_5 gpc12 (
      {stage0_0[48], stage0_0[49], stage0_0[50], stage0_0[51], stage0_0[52], stage0_0[53]},
      {stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37]},
      {stage1_4[12],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc606_5 gpc13 (
      {stage0_0[54], stage0_0[55], stage0_0[56], stage0_0[57], stage0_0[58], stage0_0[59]},
      {stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43]},
      {stage1_4[13],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc606_5 gpc14 (
      {stage0_0[60], stage0_0[61], stage0_0[62], stage0_0[63], stage0_0[64], stage0_0[65]},
      {stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49]},
      {stage1_4[14],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc606_5 gpc15 (
      {stage0_0[66], stage0_0[67], stage0_0[68], stage0_0[69], stage0_0[70], stage0_0[71]},
      {stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55]},
      {stage1_4[15],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc606_5 gpc16 (
      {stage0_0[72], stage0_0[73], stage0_0[74], stage0_0[75], stage0_0[76], stage0_0[77]},
      {stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61]},
      {stage1_4[16],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc606_5 gpc17 (
      {stage0_0[78], stage0_0[79], stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83]},
      {stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67]},
      {stage1_4[17],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc606_5 gpc18 (
      {stage0_0[84], stage0_0[85], stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89]},
      {stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73]},
      {stage1_4[18],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc606_5 gpc19 (
      {stage0_0[90], stage0_0[91], stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95]},
      {stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79]},
      {stage1_4[19],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc615_5 gpc20 (
      {stage0_0[96], stage0_0[97], stage0_0[98], stage0_0[99], stage0_0[100]},
      {stage0_1[48]},
      {stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85]},
      {stage1_4[20],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc615_5 gpc21 (
      {stage0_0[101], stage0_0[102], stage0_0[103], stage0_0[104], stage0_0[105]},
      {stage0_1[49]},
      {stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91]},
      {stage1_4[21],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc615_5 gpc22 (
      {stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109], stage0_0[110]},
      {stage0_1[50]},
      {stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97]},
      {stage1_4[22],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc615_5 gpc23 (
      {stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115]},
      {stage0_1[51]},
      {stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103]},
      {stage1_4[23],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55], stage0_1[56], stage0_1[57]},
      {stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12], stage0_3[13]},
      {stage1_5[0],stage1_4[24],stage1_3[24],stage1_2[24],stage1_1[24]}
   );
   gpc606_5 gpc25 (
      {stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61], stage0_1[62], stage0_1[63]},
      {stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18], stage0_3[19]},
      {stage1_5[1],stage1_4[25],stage1_3[25],stage1_2[25],stage1_1[25]}
   );
   gpc606_5 gpc26 (
      {stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67], stage0_1[68], stage0_1[69]},
      {stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24], stage0_3[25]},
      {stage1_5[2],stage1_4[26],stage1_3[26],stage1_2[26],stage1_1[26]}
   );
   gpc606_5 gpc27 (
      {stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73], stage0_1[74], stage0_1[75]},
      {stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29], stage0_3[30], stage0_3[31]},
      {stage1_5[3],stage1_4[27],stage1_3[27],stage1_2[27],stage1_1[27]}
   );
   gpc606_5 gpc28 (
      {stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79], stage0_1[80], stage0_1[81]},
      {stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35], stage0_3[36], stage0_3[37]},
      {stage1_5[4],stage1_4[28],stage1_3[28],stage1_2[28],stage1_1[28]}
   );
   gpc606_5 gpc29 (
      {stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85], stage0_1[86], stage0_1[87]},
      {stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41], stage0_3[42], stage0_3[43]},
      {stage1_5[5],stage1_4[29],stage1_3[29],stage1_2[29],stage1_1[29]}
   );
   gpc606_5 gpc30 (
      {stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91], stage0_1[92], stage0_1[93]},
      {stage0_3[44], stage0_3[45], stage0_3[46], stage0_3[47], stage0_3[48], stage0_3[49]},
      {stage1_5[6],stage1_4[30],stage1_3[30],stage1_2[30],stage1_1[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97], stage0_1[98], stage0_1[99]},
      {stage0_3[50], stage0_3[51], stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55]},
      {stage1_5[7],stage1_4[31],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103], stage0_1[104], stage0_1[105]},
      {stage0_3[56], stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61]},
      {stage1_5[8],stage1_4[32],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109], stage0_1[110], stage0_1[111]},
      {stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66], stage0_3[67]},
      {stage1_5[9],stage1_4[33],stage1_3[33],stage1_2[33],stage1_1[33]}
   );
   gpc606_5 gpc34 (
      {stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115], stage0_1[116], stage0_1[117]},
      {stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71], stage0_3[72], stage0_3[73]},
      {stage1_5[10],stage1_4[34],stage1_3[34],stage1_2[34],stage1_1[34]}
   );
   gpc606_5 gpc35 (
      {stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121], stage0_1[122], stage0_1[123]},
      {stage0_3[74], stage0_3[75], stage0_3[76], stage0_3[77], stage0_3[78], stage0_3[79]},
      {stage1_5[11],stage1_4[35],stage1_3[35],stage1_2[35],stage1_1[35]}
   );
   gpc1343_5 gpc36 (
      {stage0_2[104], stage0_2[105], stage0_2[106]},
      {stage0_3[80], stage0_3[81], stage0_3[82], stage0_3[83]},
      {stage0_4[0], stage0_4[1], stage0_4[2]},
      {stage0_5[0]},
      {stage1_6[0],stage1_5[12],stage1_4[36],stage1_3[36],stage1_2[36]}
   );
   gpc1163_5 gpc37 (
      {stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage0_4[3], stage0_4[4], stage0_4[5], stage0_4[6], stage0_4[7], stage0_4[8]},
      {stage0_5[1]},
      {stage0_6[0]},
      {stage1_7[0],stage1_6[1],stage1_5[13],stage1_4[37],stage1_3[37]}
   );
   gpc615_5 gpc38 (
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91]},
      {stage0_4[9]},
      {stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5], stage0_5[6], stage0_5[7]},
      {stage1_7[1],stage1_6[2],stage1_5[14],stage1_4[38],stage1_3[38]}
   );
   gpc615_5 gpc39 (
      {stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96]},
      {stage0_4[10]},
      {stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12], stage0_5[13]},
      {stage1_7[2],stage1_6[3],stage1_5[15],stage1_4[39],stage1_3[39]}
   );
   gpc615_5 gpc40 (
      {stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101]},
      {stage0_4[11]},
      {stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18], stage0_5[19]},
      {stage1_7[3],stage1_6[4],stage1_5[16],stage1_4[40],stage1_3[40]}
   );
   gpc615_5 gpc41 (
      {stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106]},
      {stage0_4[12]},
      {stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24], stage0_5[25]},
      {stage1_7[4],stage1_6[5],stage1_5[17],stage1_4[41],stage1_3[41]}
   );
   gpc615_5 gpc42 (
      {stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111]},
      {stage0_4[13]},
      {stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29], stage0_5[30], stage0_5[31]},
      {stage1_7[5],stage1_6[6],stage1_5[18],stage1_4[42],stage1_3[42]}
   );
   gpc606_5 gpc43 (
      {stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17], stage0_4[18], stage0_4[19]},
      {stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5], stage0_6[6]},
      {stage1_8[0],stage1_7[6],stage1_6[7],stage1_5[19],stage1_4[43]}
   );
   gpc606_5 gpc44 (
      {stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23], stage0_4[24], stage0_4[25]},
      {stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11], stage0_6[12]},
      {stage1_8[1],stage1_7[7],stage1_6[8],stage1_5[20],stage1_4[44]}
   );
   gpc606_5 gpc45 (
      {stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29], stage0_4[30], stage0_4[31]},
      {stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17], stage0_6[18]},
      {stage1_8[2],stage1_7[8],stage1_6[9],stage1_5[21],stage1_4[45]}
   );
   gpc606_5 gpc46 (
      {stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35], stage0_4[36], stage0_4[37]},
      {stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23], stage0_6[24]},
      {stage1_8[3],stage1_7[9],stage1_6[10],stage1_5[22],stage1_4[46]}
   );
   gpc606_5 gpc47 (
      {stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41], stage0_4[42], stage0_4[43]},
      {stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29], stage0_6[30]},
      {stage1_8[4],stage1_7[10],stage1_6[11],stage1_5[23],stage1_4[47]}
   );
   gpc606_5 gpc48 (
      {stage0_4[44], stage0_4[45], stage0_4[46], stage0_4[47], stage0_4[48], stage0_4[49]},
      {stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35], stage0_6[36]},
      {stage1_8[5],stage1_7[11],stage1_6[12],stage1_5[24],stage1_4[48]}
   );
   gpc606_5 gpc49 (
      {stage0_4[50], stage0_4[51], stage0_4[52], stage0_4[53], stage0_4[54], stage0_4[55]},
      {stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41], stage0_6[42]},
      {stage1_8[6],stage1_7[12],stage1_6[13],stage1_5[25],stage1_4[49]}
   );
   gpc606_5 gpc50 (
      {stage0_4[56], stage0_4[57], stage0_4[58], stage0_4[59], stage0_4[60], stage0_4[61]},
      {stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47], stage0_6[48]},
      {stage1_8[7],stage1_7[13],stage1_6[14],stage1_5[26],stage1_4[50]}
   );
   gpc606_5 gpc51 (
      {stage0_4[62], stage0_4[63], stage0_4[64], stage0_4[65], stage0_4[66], stage0_4[67]},
      {stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53], stage0_6[54]},
      {stage1_8[8],stage1_7[14],stage1_6[15],stage1_5[27],stage1_4[51]}
   );
   gpc606_5 gpc52 (
      {stage0_4[68], stage0_4[69], stage0_4[70], stage0_4[71], stage0_4[72], stage0_4[73]},
      {stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59], stage0_6[60]},
      {stage1_8[9],stage1_7[15],stage1_6[16],stage1_5[28],stage1_4[52]}
   );
   gpc606_5 gpc53 (
      {stage0_4[74], stage0_4[75], stage0_4[76], stage0_4[77], stage0_4[78], stage0_4[79]},
      {stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65], stage0_6[66]},
      {stage1_8[10],stage1_7[16],stage1_6[17],stage1_5[29],stage1_4[53]}
   );
   gpc606_5 gpc54 (
      {stage0_4[80], stage0_4[81], stage0_4[82], stage0_4[83], stage0_4[84], stage0_4[85]},
      {stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71], stage0_6[72]},
      {stage1_8[11],stage1_7[17],stage1_6[18],stage1_5[30],stage1_4[54]}
   );
   gpc606_5 gpc55 (
      {stage0_4[86], stage0_4[87], stage0_4[88], stage0_4[89], stage0_4[90], stage0_4[91]},
      {stage0_6[73], stage0_6[74], stage0_6[75], stage0_6[76], stage0_6[77], stage0_6[78]},
      {stage1_8[12],stage1_7[18],stage1_6[19],stage1_5[31],stage1_4[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[92], stage0_4[93], stage0_4[94], stage0_4[95], stage0_4[96], stage0_4[97]},
      {stage0_6[79], stage0_6[80], stage0_6[81], stage0_6[82], stage0_6[83], stage0_6[84]},
      {stage1_8[13],stage1_7[19],stage1_6[20],stage1_5[32],stage1_4[56]}
   );
   gpc606_5 gpc57 (
      {stage0_4[98], stage0_4[99], stage0_4[100], stage0_4[101], stage0_4[102], stage0_4[103]},
      {stage0_6[85], stage0_6[86], stage0_6[87], stage0_6[88], stage0_6[89], stage0_6[90]},
      {stage1_8[14],stage1_7[20],stage1_6[21],stage1_5[33],stage1_4[57]}
   );
   gpc606_5 gpc58 (
      {stage0_4[104], stage0_4[105], stage0_4[106], stage0_4[107], stage0_4[108], stage0_4[109]},
      {stage0_6[91], stage0_6[92], stage0_6[93], stage0_6[94], stage0_6[95], stage0_6[96]},
      {stage1_8[15],stage1_7[21],stage1_6[22],stage1_5[34],stage1_4[58]}
   );
   gpc606_5 gpc59 (
      {stage0_4[110], stage0_4[111], stage0_4[112], stage0_4[113], stage0_4[114], stage0_4[115]},
      {stage0_6[97], stage0_6[98], stage0_6[99], stage0_6[100], stage0_6[101], stage0_6[102]},
      {stage1_8[16],stage1_7[22],stage1_6[23],stage1_5[35],stage1_4[59]}
   );
   gpc606_5 gpc60 (
      {stage0_4[116], stage0_4[117], stage0_4[118], stage0_4[119], stage0_4[120], stage0_4[121]},
      {stage0_6[103], stage0_6[104], stage0_6[105], stage0_6[106], stage0_6[107], stage0_6[108]},
      {stage1_8[17],stage1_7[23],stage1_6[24],stage1_5[36],stage1_4[60]}
   );
   gpc606_5 gpc61 (
      {stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35], stage0_5[36], stage0_5[37]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[18],stage1_7[24],stage1_6[25],stage1_5[37]}
   );
   gpc606_5 gpc62 (
      {stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41], stage0_5[42], stage0_5[43]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[19],stage1_7[25],stage1_6[26],stage1_5[38]}
   );
   gpc606_5 gpc63 (
      {stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47], stage0_5[48], stage0_5[49]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[20],stage1_7[26],stage1_6[27],stage1_5[39]}
   );
   gpc606_5 gpc64 (
      {stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53], stage0_5[54], stage0_5[55]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[21],stage1_7[27],stage1_6[28],stage1_5[40]}
   );
   gpc606_5 gpc65 (
      {stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59], stage0_5[60], stage0_5[61]},
      {stage0_7[24], stage0_7[25], stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29]},
      {stage1_9[4],stage1_8[22],stage1_7[28],stage1_6[29],stage1_5[41]}
   );
   gpc606_5 gpc66 (
      {stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65], stage0_5[66], stage0_5[67]},
      {stage0_7[30], stage0_7[31], stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35]},
      {stage1_9[5],stage1_8[23],stage1_7[29],stage1_6[30],stage1_5[42]}
   );
   gpc606_5 gpc67 (
      {stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71], stage0_5[72], stage0_5[73]},
      {stage0_7[36], stage0_7[37], stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41]},
      {stage1_9[6],stage1_8[24],stage1_7[30],stage1_6[31],stage1_5[43]}
   );
   gpc606_5 gpc68 (
      {stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77], stage0_5[78], stage0_5[79]},
      {stage0_7[42], stage0_7[43], stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47]},
      {stage1_9[7],stage1_8[25],stage1_7[31],stage1_6[32],stage1_5[44]}
   );
   gpc606_5 gpc69 (
      {stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83], stage0_5[84], stage0_5[85]},
      {stage0_7[48], stage0_7[49], stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53]},
      {stage1_9[8],stage1_8[26],stage1_7[32],stage1_6[33],stage1_5[45]}
   );
   gpc606_5 gpc70 (
      {stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89], stage0_5[90], stage0_5[91]},
      {stage0_7[54], stage0_7[55], stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59]},
      {stage1_9[9],stage1_8[27],stage1_7[33],stage1_6[34],stage1_5[46]}
   );
   gpc606_5 gpc71 (
      {stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95], stage0_5[96], stage0_5[97]},
      {stage0_7[60], stage0_7[61], stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65]},
      {stage1_9[10],stage1_8[28],stage1_7[34],stage1_6[35],stage1_5[47]}
   );
   gpc606_5 gpc72 (
      {stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101], stage0_5[102], stage0_5[103]},
      {stage0_7[66], stage0_7[67], stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71]},
      {stage1_9[11],stage1_8[29],stage1_7[35],stage1_6[36],stage1_5[48]}
   );
   gpc606_5 gpc73 (
      {stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107], stage0_5[108], stage0_5[109]},
      {stage0_7[72], stage0_7[73], stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77]},
      {stage1_9[12],stage1_8[30],stage1_7[36],stage1_6[37],stage1_5[49]}
   );
   gpc606_5 gpc74 (
      {stage0_5[110], stage0_5[111], stage0_5[112], stage0_5[113], stage0_5[114], stage0_5[115]},
      {stage0_7[78], stage0_7[79], stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83]},
      {stage1_9[13],stage1_8[31],stage1_7[37],stage1_6[38],stage1_5[50]}
   );
   gpc615_5 gpc75 (
      {stage0_6[109], stage0_6[110], stage0_6[111], stage0_6[112], stage0_6[113]},
      {stage0_7[84]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[14],stage1_8[32],stage1_7[38],stage1_6[39]}
   );
   gpc615_5 gpc76 (
      {stage0_6[114], stage0_6[115], stage0_6[116], stage0_6[117], stage0_6[118]},
      {stage0_7[85]},
      {stage0_8[6], stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11]},
      {stage1_10[1],stage1_9[15],stage1_8[33],stage1_7[39],stage1_6[40]}
   );
   gpc615_5 gpc77 (
      {stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89], stage0_7[90]},
      {stage0_8[12]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[2],stage1_9[16],stage1_8[34],stage1_7[40]}
   );
   gpc615_5 gpc78 (
      {stage0_7[91], stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95]},
      {stage0_8[13]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[3],stage1_9[17],stage1_8[35],stage1_7[41]}
   );
   gpc615_5 gpc79 (
      {stage0_7[96], stage0_7[97], stage0_7[98], stage0_7[99], stage0_7[100]},
      {stage0_8[14]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[4],stage1_9[18],stage1_8[36],stage1_7[42]}
   );
   gpc207_4 gpc80 (
      {stage0_8[15], stage0_8[16], stage0_8[17], stage0_8[18], stage0_8[19], stage0_8[20], stage0_8[21]},
      {stage0_10[0], stage0_10[1]},
      {stage1_11[3],stage1_10[5],stage1_9[19],stage1_8[37]}
   );
   gpc606_5 gpc81 (
      {stage0_8[22], stage0_8[23], stage0_8[24], stage0_8[25], stage0_8[26], stage0_8[27]},
      {stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5], stage0_10[6], stage0_10[7]},
      {stage1_12[0],stage1_11[4],stage1_10[6],stage1_9[20],stage1_8[38]}
   );
   gpc606_5 gpc82 (
      {stage0_8[28], stage0_8[29], stage0_8[30], stage0_8[31], stage0_8[32], stage0_8[33]},
      {stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11], stage0_10[12], stage0_10[13]},
      {stage1_12[1],stage1_11[5],stage1_10[7],stage1_9[21],stage1_8[39]}
   );
   gpc606_5 gpc83 (
      {stage0_8[34], stage0_8[35], stage0_8[36], stage0_8[37], stage0_8[38], stage0_8[39]},
      {stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17], stage0_10[18], stage0_10[19]},
      {stage1_12[2],stage1_11[6],stage1_10[8],stage1_9[22],stage1_8[40]}
   );
   gpc606_5 gpc84 (
      {stage0_8[40], stage0_8[41], stage0_8[42], stage0_8[43], stage0_8[44], stage0_8[45]},
      {stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23], stage0_10[24], stage0_10[25]},
      {stage1_12[3],stage1_11[7],stage1_10[9],stage1_9[23],stage1_8[41]}
   );
   gpc606_5 gpc85 (
      {stage0_8[46], stage0_8[47], stage0_8[48], stage0_8[49], stage0_8[50], stage0_8[51]},
      {stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29], stage0_10[30], stage0_10[31]},
      {stage1_12[4],stage1_11[8],stage1_10[10],stage1_9[24],stage1_8[42]}
   );
   gpc606_5 gpc86 (
      {stage0_8[52], stage0_8[53], stage0_8[54], stage0_8[55], stage0_8[56], stage0_8[57]},
      {stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35], stage0_10[36], stage0_10[37]},
      {stage1_12[5],stage1_11[9],stage1_10[11],stage1_9[25],stage1_8[43]}
   );
   gpc606_5 gpc87 (
      {stage0_8[58], stage0_8[59], stage0_8[60], stage0_8[61], stage0_8[62], stage0_8[63]},
      {stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41], stage0_10[42], stage0_10[43]},
      {stage1_12[6],stage1_11[10],stage1_10[12],stage1_9[26],stage1_8[44]}
   );
   gpc606_5 gpc88 (
      {stage0_8[64], stage0_8[65], stage0_8[66], stage0_8[67], stage0_8[68], stage0_8[69]},
      {stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47], stage0_10[48], stage0_10[49]},
      {stage1_12[7],stage1_11[11],stage1_10[13],stage1_9[27],stage1_8[45]}
   );
   gpc606_5 gpc89 (
      {stage0_8[70], stage0_8[71], stage0_8[72], stage0_8[73], stage0_8[74], stage0_8[75]},
      {stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53], stage0_10[54], stage0_10[55]},
      {stage1_12[8],stage1_11[12],stage1_10[14],stage1_9[28],stage1_8[46]}
   );
   gpc606_5 gpc90 (
      {stage0_8[76], stage0_8[77], stage0_8[78], stage0_8[79], stage0_8[80], stage0_8[81]},
      {stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59], stage0_10[60], stage0_10[61]},
      {stage1_12[9],stage1_11[13],stage1_10[15],stage1_9[29],stage1_8[47]}
   );
   gpc606_5 gpc91 (
      {stage0_8[82], stage0_8[83], stage0_8[84], stage0_8[85], stage0_8[86], stage0_8[87]},
      {stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65], stage0_10[66], stage0_10[67]},
      {stage1_12[10],stage1_11[14],stage1_10[16],stage1_9[30],stage1_8[48]}
   );
   gpc606_5 gpc92 (
      {stage0_8[88], stage0_8[89], stage0_8[90], stage0_8[91], stage0_8[92], stage0_8[93]},
      {stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71], stage0_10[72], stage0_10[73]},
      {stage1_12[11],stage1_11[15],stage1_10[17],stage1_9[31],stage1_8[49]}
   );
   gpc606_5 gpc93 (
      {stage0_8[94], stage0_8[95], stage0_8[96], stage0_8[97], stage0_8[98], stage0_8[99]},
      {stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77], stage0_10[78], stage0_10[79]},
      {stage1_12[12],stage1_11[16],stage1_10[18],stage1_9[32],stage1_8[50]}
   );
   gpc606_5 gpc94 (
      {stage0_8[100], stage0_8[101], stage0_8[102], stage0_8[103], stage0_8[104], stage0_8[105]},
      {stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83], stage0_10[84], stage0_10[85]},
      {stage1_12[13],stage1_11[17],stage1_10[19],stage1_9[33],stage1_8[51]}
   );
   gpc606_5 gpc95 (
      {stage0_8[106], stage0_8[107], stage0_8[108], stage0_8[109], stage0_8[110], stage0_8[111]},
      {stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89], stage0_10[90], stage0_10[91]},
      {stage1_12[14],stage1_11[18],stage1_10[20],stage1_9[34],stage1_8[52]}
   );
   gpc606_5 gpc96 (
      {stage0_8[112], stage0_8[113], stage0_8[114], stage0_8[115], stage0_8[116], stage0_8[117]},
      {stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95], stage0_10[96], stage0_10[97]},
      {stage1_12[15],stage1_11[19],stage1_10[21],stage1_9[35],stage1_8[53]}
   );
   gpc615_5 gpc97 (
      {stage0_8[118], stage0_8[119], stage0_8[120], stage0_8[121], stage0_8[122]},
      {stage0_9[18]},
      {stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101], stage0_10[102], stage0_10[103]},
      {stage1_12[16],stage1_11[20],stage1_10[22],stage1_9[36],stage1_8[54]}
   );
   gpc615_5 gpc98 (
      {stage0_8[123], stage0_8[124], stage0_8[125], stage0_8[126], stage0_8[127]},
      {stage0_9[19]},
      {stage0_10[104], stage0_10[105], stage0_10[106], stage0_10[107], stage0_10[108], stage0_10[109]},
      {stage1_12[17],stage1_11[21],stage1_10[23],stage1_9[37],stage1_8[55]}
   );
   gpc606_5 gpc99 (
      {stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23], stage0_9[24], stage0_9[25]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[18],stage1_11[22],stage1_10[24],stage1_9[38]}
   );
   gpc606_5 gpc100 (
      {stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29], stage0_9[30], stage0_9[31]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[19],stage1_11[23],stage1_10[25],stage1_9[39]}
   );
   gpc606_5 gpc101 (
      {stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35], stage0_9[36], stage0_9[37]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[20],stage1_11[24],stage1_10[26],stage1_9[40]}
   );
   gpc606_5 gpc102 (
      {stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41], stage0_9[42], stage0_9[43]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[21],stage1_11[25],stage1_10[27],stage1_9[41]}
   );
   gpc606_5 gpc103 (
      {stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47], stage0_9[48], stage0_9[49]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[22],stage1_11[26],stage1_10[28],stage1_9[42]}
   );
   gpc606_5 gpc104 (
      {stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53], stage0_9[54], stage0_9[55]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[23],stage1_11[27],stage1_10[29],stage1_9[43]}
   );
   gpc606_5 gpc105 (
      {stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59], stage0_9[60], stage0_9[61]},
      {stage0_11[36], stage0_11[37], stage0_11[38], stage0_11[39], stage0_11[40], stage0_11[41]},
      {stage1_13[6],stage1_12[24],stage1_11[28],stage1_10[30],stage1_9[44]}
   );
   gpc606_5 gpc106 (
      {stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65], stage0_9[66], stage0_9[67]},
      {stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46], stage0_11[47]},
      {stage1_13[7],stage1_12[25],stage1_11[29],stage1_10[31],stage1_9[45]}
   );
   gpc606_5 gpc107 (
      {stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71], stage0_9[72], stage0_9[73]},
      {stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage1_13[8],stage1_12[26],stage1_11[30],stage1_10[32],stage1_9[46]}
   );
   gpc606_5 gpc108 (
      {stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77], stage0_9[78], stage0_9[79]},
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59]},
      {stage1_13[9],stage1_12[27],stage1_11[31],stage1_10[33],stage1_9[47]}
   );
   gpc606_5 gpc109 (
      {stage0_9[80], stage0_9[81], stage0_9[82], stage0_9[83], stage0_9[84], stage0_9[85]},
      {stage0_11[60], stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65]},
      {stage1_13[10],stage1_12[28],stage1_11[32],stage1_10[34],stage1_9[48]}
   );
   gpc606_5 gpc110 (
      {stage0_9[86], stage0_9[87], stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91]},
      {stage0_11[66], stage0_11[67], stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71]},
      {stage1_13[11],stage1_12[29],stage1_11[33],stage1_10[35],stage1_9[49]}
   );
   gpc606_5 gpc111 (
      {stage0_9[92], stage0_9[93], stage0_9[94], stage0_9[95], stage0_9[96], stage0_9[97]},
      {stage0_11[72], stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage1_13[12],stage1_12[30],stage1_11[34],stage1_10[36],stage1_9[50]}
   );
   gpc606_5 gpc112 (
      {stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101], stage0_9[102], stage0_9[103]},
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82], stage0_11[83]},
      {stage1_13[13],stage1_12[31],stage1_11[35],stage1_10[37],stage1_9[51]}
   );
   gpc606_5 gpc113 (
      {stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107], stage0_9[108], stage0_9[109]},
      {stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87], stage0_11[88], stage0_11[89]},
      {stage1_13[14],stage1_12[32],stage1_11[36],stage1_10[38],stage1_9[52]}
   );
   gpc606_5 gpc114 (
      {stage0_9[110], stage0_9[111], stage0_9[112], stage0_9[113], stage0_9[114], stage0_9[115]},
      {stage0_11[90], stage0_11[91], stage0_11[92], stage0_11[93], stage0_11[94], stage0_11[95]},
      {stage1_13[15],stage1_12[33],stage1_11[37],stage1_10[39],stage1_9[53]}
   );
   gpc606_5 gpc115 (
      {stage0_9[116], stage0_9[117], stage0_9[118], stage0_9[119], stage0_9[120], stage0_9[121]},
      {stage0_11[96], stage0_11[97], stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101]},
      {stage1_13[16],stage1_12[34],stage1_11[38],stage1_10[40],stage1_9[54]}
   );
   gpc606_5 gpc116 (
      {stage0_10[110], stage0_10[111], stage0_10[112], stage0_10[113], stage0_10[114], stage0_10[115]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[17],stage1_12[35],stage1_11[39],stage1_10[41]}
   );
   gpc615_5 gpc117 (
      {stage0_11[102], stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106]},
      {stage0_12[6]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[1],stage1_13[18],stage1_12[36],stage1_11[40]}
   );
   gpc615_5 gpc118 (
      {stage0_11[107], stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111]},
      {stage0_12[7]},
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage1_15[1],stage1_14[2],stage1_13[19],stage1_12[37],stage1_11[41]}
   );
   gpc606_5 gpc119 (
      {stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11], stage0_12[12], stage0_12[13]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[2],stage1_14[3],stage1_13[20],stage1_12[38]}
   );
   gpc606_5 gpc120 (
      {stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17], stage0_12[18], stage0_12[19]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[3],stage1_14[4],stage1_13[21],stage1_12[39]}
   );
   gpc606_5 gpc121 (
      {stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23], stage0_12[24], stage0_12[25]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[4],stage1_14[5],stage1_13[22],stage1_12[40]}
   );
   gpc606_5 gpc122 (
      {stage0_12[26], stage0_12[27], stage0_12[28], stage0_12[29], stage0_12[30], stage0_12[31]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[5],stage1_14[6],stage1_13[23],stage1_12[41]}
   );
   gpc606_5 gpc123 (
      {stage0_12[32], stage0_12[33], stage0_12[34], stage0_12[35], stage0_12[36], stage0_12[37]},
      {stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27], stage0_14[28], stage0_14[29]},
      {stage1_16[4],stage1_15[6],stage1_14[7],stage1_13[24],stage1_12[42]}
   );
   gpc606_5 gpc124 (
      {stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41], stage0_12[42], stage0_12[43]},
      {stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33], stage0_14[34], stage0_14[35]},
      {stage1_16[5],stage1_15[7],stage1_14[8],stage1_13[25],stage1_12[43]}
   );
   gpc606_5 gpc125 (
      {stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47], stage0_12[48], stage0_12[49]},
      {stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39], stage0_14[40], stage0_14[41]},
      {stage1_16[6],stage1_15[8],stage1_14[9],stage1_13[26],stage1_12[44]}
   );
   gpc606_5 gpc126 (
      {stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53], stage0_12[54], stage0_12[55]},
      {stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45], stage0_14[46], stage0_14[47]},
      {stage1_16[7],stage1_15[9],stage1_14[10],stage1_13[27],stage1_12[45]}
   );
   gpc606_5 gpc127 (
      {stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59], stage0_12[60], stage0_12[61]},
      {stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51], stage0_14[52], stage0_14[53]},
      {stage1_16[8],stage1_15[10],stage1_14[11],stage1_13[28],stage1_12[46]}
   );
   gpc606_5 gpc128 (
      {stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65], stage0_12[66], stage0_12[67]},
      {stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57], stage0_14[58], stage0_14[59]},
      {stage1_16[9],stage1_15[11],stage1_14[12],stage1_13[29],stage1_12[47]}
   );
   gpc606_5 gpc129 (
      {stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71], stage0_12[72], stage0_12[73]},
      {stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63], stage0_14[64], stage0_14[65]},
      {stage1_16[10],stage1_15[12],stage1_14[13],stage1_13[30],stage1_12[48]}
   );
   gpc606_5 gpc130 (
      {stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77], stage0_12[78], stage0_12[79]},
      {stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69], stage0_14[70], stage0_14[71]},
      {stage1_16[11],stage1_15[13],stage1_14[14],stage1_13[31],stage1_12[49]}
   );
   gpc606_5 gpc131 (
      {stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83], stage0_12[84], stage0_12[85]},
      {stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75], stage0_14[76], stage0_14[77]},
      {stage1_16[12],stage1_15[14],stage1_14[15],stage1_13[32],stage1_12[50]}
   );
   gpc606_5 gpc132 (
      {stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89], stage0_12[90], stage0_12[91]},
      {stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81], stage0_14[82], stage0_14[83]},
      {stage1_16[13],stage1_15[15],stage1_14[16],stage1_13[33],stage1_12[51]}
   );
   gpc606_5 gpc133 (
      {stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95], stage0_12[96], stage0_12[97]},
      {stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87], stage0_14[88], stage0_14[89]},
      {stage1_16[14],stage1_15[16],stage1_14[17],stage1_13[34],stage1_12[52]}
   );
   gpc606_5 gpc134 (
      {stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101], stage0_12[102], stage0_12[103]},
      {stage0_14[90], stage0_14[91], stage0_14[92], stage0_14[93], stage0_14[94], stage0_14[95]},
      {stage1_16[15],stage1_15[17],stage1_14[18],stage1_13[35],stage1_12[53]}
   );
   gpc606_5 gpc135 (
      {stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107], stage0_12[108], stage0_12[109]},
      {stage0_14[96], stage0_14[97], stage0_14[98], stage0_14[99], stage0_14[100], stage0_14[101]},
      {stage1_16[16],stage1_15[18],stage1_14[19],stage1_13[36],stage1_12[54]}
   );
   gpc606_5 gpc136 (
      {stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113], stage0_12[114], stage0_12[115]},
      {stage0_14[102], stage0_14[103], stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107]},
      {stage1_16[17],stage1_15[19],stage1_14[20],stage1_13[37],stage1_12[55]}
   );
   gpc606_5 gpc137 (
      {stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121]},
      {stage0_14[108], stage0_14[109], stage0_14[110], stage0_14[111], stage0_14[112], stage0_14[113]},
      {stage1_16[18],stage1_15[20],stage1_14[21],stage1_13[38],stage1_12[56]}
   );
   gpc606_5 gpc138 (
      {stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127]},
      {stage0_14[114], stage0_14[115], stage0_14[116], stage0_14[117], stage0_14[118], stage0_14[119]},
      {stage1_16[19],stage1_15[21],stage1_14[22],stage1_13[39],stage1_12[57]}
   );
   gpc606_5 gpc139 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[20],stage1_15[22],stage1_14[23],stage1_13[40]}
   );
   gpc606_5 gpc140 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[21],stage1_15[23],stage1_14[24],stage1_13[41]}
   );
   gpc606_5 gpc141 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[22],stage1_15[24],stage1_14[25],stage1_13[42]}
   );
   gpc606_5 gpc142 (
      {stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33], stage0_13[34], stage0_13[35]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[23],stage1_15[25],stage1_14[26],stage1_13[43]}
   );
   gpc606_5 gpc143 (
      {stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39], stage0_13[40], stage0_13[41]},
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29]},
      {stage1_17[4],stage1_16[24],stage1_15[26],stage1_14[27],stage1_13[44]}
   );
   gpc606_5 gpc144 (
      {stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45], stage0_13[46], stage0_13[47]},
      {stage0_15[30], stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35]},
      {stage1_17[5],stage1_16[25],stage1_15[27],stage1_14[28],stage1_13[45]}
   );
   gpc606_5 gpc145 (
      {stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51], stage0_13[52], stage0_13[53]},
      {stage0_15[36], stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41]},
      {stage1_17[6],stage1_16[26],stage1_15[28],stage1_14[29],stage1_13[46]}
   );
   gpc606_5 gpc146 (
      {stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57], stage0_13[58], stage0_13[59]},
      {stage0_15[42], stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47]},
      {stage1_17[7],stage1_16[27],stage1_15[29],stage1_14[30],stage1_13[47]}
   );
   gpc606_5 gpc147 (
      {stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63], stage0_13[64], stage0_13[65]},
      {stage0_15[48], stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53]},
      {stage1_17[8],stage1_16[28],stage1_15[30],stage1_14[31],stage1_13[48]}
   );
   gpc606_5 gpc148 (
      {stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69], stage0_13[70], stage0_13[71]},
      {stage0_15[54], stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59]},
      {stage1_17[9],stage1_16[29],stage1_15[31],stage1_14[32],stage1_13[49]}
   );
   gpc606_5 gpc149 (
      {stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75], stage0_13[76], stage0_13[77]},
      {stage0_15[60], stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65]},
      {stage1_17[10],stage1_16[30],stage1_15[32],stage1_14[33],stage1_13[50]}
   );
   gpc606_5 gpc150 (
      {stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81], stage0_13[82], stage0_13[83]},
      {stage0_15[66], stage0_15[67], stage0_15[68], stage0_15[69], stage0_15[70], stage0_15[71]},
      {stage1_17[11],stage1_16[31],stage1_15[33],stage1_14[34],stage1_13[51]}
   );
   gpc606_5 gpc151 (
      {stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87], stage0_13[88], stage0_13[89]},
      {stage0_15[72], stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77]},
      {stage1_17[12],stage1_16[32],stage1_15[34],stage1_14[35],stage1_13[52]}
   );
   gpc606_5 gpc152 (
      {stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93], stage0_13[94], stage0_13[95]},
      {stage0_15[78], stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83]},
      {stage1_17[13],stage1_16[33],stage1_15[35],stage1_14[36],stage1_13[53]}
   );
   gpc606_5 gpc153 (
      {stage0_13[96], stage0_13[97], stage0_13[98], stage0_13[99], stage0_13[100], stage0_13[101]},
      {stage0_15[84], stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89]},
      {stage1_17[14],stage1_16[34],stage1_15[36],stage1_14[37],stage1_13[54]}
   );
   gpc606_5 gpc154 (
      {stage0_13[102], stage0_13[103], stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107]},
      {stage0_15[90], stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage1_17[15],stage1_16[35],stage1_15[37],stage1_14[38],stage1_13[55]}
   );
   gpc606_5 gpc155 (
      {stage0_13[108], stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100], stage0_15[101]},
      {stage1_17[16],stage1_16[36],stage1_15[38],stage1_14[39],stage1_13[56]}
   );
   gpc606_5 gpc156 (
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118], stage0_13[119]},
      {stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105], stage0_15[106], stage0_15[107]},
      {stage1_17[17],stage1_16[37],stage1_15[39],stage1_14[40],stage1_13[57]}
   );
   gpc606_5 gpc157 (
      {stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123], stage0_13[124], stage0_13[125]},
      {stage0_15[108], stage0_15[109], stage0_15[110], stage0_15[111], stage0_15[112], stage0_15[113]},
      {stage1_17[18],stage1_16[38],stage1_15[40],stage1_14[41],stage1_13[58]}
   );
   gpc615_5 gpc158 (
      {stage0_14[120], stage0_14[121], stage0_14[122], stage0_14[123], stage0_14[124]},
      {stage0_15[114]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[19],stage1_16[39],stage1_15[41],stage1_14[42]}
   );
   gpc615_5 gpc159 (
      {stage0_15[115], stage0_15[116], stage0_15[117], stage0_15[118], stage0_15[119]},
      {stage0_16[6]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[1],stage1_17[20],stage1_16[40],stage1_15[42]}
   );
   gpc615_5 gpc160 (
      {stage0_15[120], stage0_15[121], stage0_15[122], stage0_15[123], stage0_15[124]},
      {stage0_16[7]},
      {stage0_17[6], stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11]},
      {stage1_19[1],stage1_18[2],stage1_17[21],stage1_16[41],stage1_15[43]}
   );
   gpc606_5 gpc161 (
      {stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11], stage0_16[12], stage0_16[13]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[2],stage1_18[3],stage1_17[22],stage1_16[42]}
   );
   gpc606_5 gpc162 (
      {stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17], stage0_16[18], stage0_16[19]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[3],stage1_18[4],stage1_17[23],stage1_16[43]}
   );
   gpc606_5 gpc163 (
      {stage0_16[20], stage0_16[21], stage0_16[22], stage0_16[23], stage0_16[24], stage0_16[25]},
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage1_20[2],stage1_19[4],stage1_18[5],stage1_17[24],stage1_16[44]}
   );
   gpc606_5 gpc164 (
      {stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29], stage0_16[30], stage0_16[31]},
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage1_20[3],stage1_19[5],stage1_18[6],stage1_17[25],stage1_16[45]}
   );
   gpc606_5 gpc165 (
      {stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35], stage0_16[36], stage0_16[37]},
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29]},
      {stage1_20[4],stage1_19[6],stage1_18[7],stage1_17[26],stage1_16[46]}
   );
   gpc606_5 gpc166 (
      {stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41], stage0_16[42], stage0_16[43]},
      {stage0_18[30], stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35]},
      {stage1_20[5],stage1_19[7],stage1_18[8],stage1_17[27],stage1_16[47]}
   );
   gpc606_5 gpc167 (
      {stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47], stage0_16[48], stage0_16[49]},
      {stage0_18[36], stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41]},
      {stage1_20[6],stage1_19[8],stage1_18[9],stage1_17[28],stage1_16[48]}
   );
   gpc606_5 gpc168 (
      {stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53], stage0_16[54], stage0_16[55]},
      {stage0_18[42], stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47]},
      {stage1_20[7],stage1_19[9],stage1_18[10],stage1_17[29],stage1_16[49]}
   );
   gpc606_5 gpc169 (
      {stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59], stage0_16[60], stage0_16[61]},
      {stage0_18[48], stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53]},
      {stage1_20[8],stage1_19[10],stage1_18[11],stage1_17[30],stage1_16[50]}
   );
   gpc606_5 gpc170 (
      {stage0_16[62], stage0_16[63], stage0_16[64], stage0_16[65], stage0_16[66], stage0_16[67]},
      {stage0_18[54], stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59]},
      {stage1_20[9],stage1_19[11],stage1_18[12],stage1_17[31],stage1_16[51]}
   );
   gpc606_5 gpc171 (
      {stage0_16[68], stage0_16[69], stage0_16[70], stage0_16[71], stage0_16[72], stage0_16[73]},
      {stage0_18[60], stage0_18[61], stage0_18[62], stage0_18[63], stage0_18[64], stage0_18[65]},
      {stage1_20[10],stage1_19[12],stage1_18[13],stage1_17[32],stage1_16[52]}
   );
   gpc606_5 gpc172 (
      {stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77], stage0_16[78], stage0_16[79]},
      {stage0_18[66], stage0_18[67], stage0_18[68], stage0_18[69], stage0_18[70], stage0_18[71]},
      {stage1_20[11],stage1_19[13],stage1_18[14],stage1_17[33],stage1_16[53]}
   );
   gpc606_5 gpc173 (
      {stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83], stage0_16[84], stage0_16[85]},
      {stage0_18[72], stage0_18[73], stage0_18[74], stage0_18[75], stage0_18[76], stage0_18[77]},
      {stage1_20[12],stage1_19[14],stage1_18[15],stage1_17[34],stage1_16[54]}
   );
   gpc606_5 gpc174 (
      {stage0_16[86], stage0_16[87], stage0_16[88], stage0_16[89], stage0_16[90], stage0_16[91]},
      {stage0_18[78], stage0_18[79], stage0_18[80], stage0_18[81], stage0_18[82], stage0_18[83]},
      {stage1_20[13],stage1_19[15],stage1_18[16],stage1_17[35],stage1_16[55]}
   );
   gpc606_5 gpc175 (
      {stage0_16[92], stage0_16[93], stage0_16[94], stage0_16[95], stage0_16[96], stage0_16[97]},
      {stage0_18[84], stage0_18[85], stage0_18[86], stage0_18[87], stage0_18[88], stage0_18[89]},
      {stage1_20[14],stage1_19[16],stage1_18[17],stage1_17[36],stage1_16[56]}
   );
   gpc606_5 gpc176 (
      {stage0_17[12], stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[15],stage1_19[17],stage1_18[18],stage1_17[37]}
   );
   gpc606_5 gpc177 (
      {stage0_17[18], stage0_17[19], stage0_17[20], stage0_17[21], stage0_17[22], stage0_17[23]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[16],stage1_19[18],stage1_18[19],stage1_17[38]}
   );
   gpc606_5 gpc178 (
      {stage0_17[24], stage0_17[25], stage0_17[26], stage0_17[27], stage0_17[28], stage0_17[29]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[17],stage1_19[19],stage1_18[20],stage1_17[39]}
   );
   gpc606_5 gpc179 (
      {stage0_17[30], stage0_17[31], stage0_17[32], stage0_17[33], stage0_17[34], stage0_17[35]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[18],stage1_19[20],stage1_18[21],stage1_17[40]}
   );
   gpc606_5 gpc180 (
      {stage0_17[36], stage0_17[37], stage0_17[38], stage0_17[39], stage0_17[40], stage0_17[41]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[19],stage1_19[21],stage1_18[22],stage1_17[41]}
   );
   gpc606_5 gpc181 (
      {stage0_17[42], stage0_17[43], stage0_17[44], stage0_17[45], stage0_17[46], stage0_17[47]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[20],stage1_19[22],stage1_18[23],stage1_17[42]}
   );
   gpc606_5 gpc182 (
      {stage0_17[48], stage0_17[49], stage0_17[50], stage0_17[51], stage0_17[52], stage0_17[53]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[21],stage1_19[23],stage1_18[24],stage1_17[43]}
   );
   gpc606_5 gpc183 (
      {stage0_17[54], stage0_17[55], stage0_17[56], stage0_17[57], stage0_17[58], stage0_17[59]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[22],stage1_19[24],stage1_18[25],stage1_17[44]}
   );
   gpc606_5 gpc184 (
      {stage0_17[60], stage0_17[61], stage0_17[62], stage0_17[63], stage0_17[64], stage0_17[65]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[23],stage1_19[25],stage1_18[26],stage1_17[45]}
   );
   gpc606_5 gpc185 (
      {stage0_17[66], stage0_17[67], stage0_17[68], stage0_17[69], stage0_17[70], stage0_17[71]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[24],stage1_19[26],stage1_18[27],stage1_17[46]}
   );
   gpc606_5 gpc186 (
      {stage0_17[72], stage0_17[73], stage0_17[74], stage0_17[75], stage0_17[76], stage0_17[77]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[25],stage1_19[27],stage1_18[28],stage1_17[47]}
   );
   gpc606_5 gpc187 (
      {stage0_17[78], stage0_17[79], stage0_17[80], stage0_17[81], stage0_17[82], stage0_17[83]},
      {stage0_19[66], stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71]},
      {stage1_21[11],stage1_20[26],stage1_19[28],stage1_18[29],stage1_17[48]}
   );
   gpc606_5 gpc188 (
      {stage0_17[84], stage0_17[85], stage0_17[86], stage0_17[87], stage0_17[88], stage0_17[89]},
      {stage0_19[72], stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage1_21[12],stage1_20[27],stage1_19[29],stage1_18[30],stage1_17[49]}
   );
   gpc606_5 gpc189 (
      {stage0_17[90], stage0_17[91], stage0_17[92], stage0_17[93], stage0_17[94], stage0_17[95]},
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82], stage0_19[83]},
      {stage1_21[13],stage1_20[28],stage1_19[30],stage1_18[31],stage1_17[50]}
   );
   gpc606_5 gpc190 (
      {stage0_17[96], stage0_17[97], stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101]},
      {stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87], stage0_19[88], stage0_19[89]},
      {stage1_21[14],stage1_20[29],stage1_19[31],stage1_18[32],stage1_17[51]}
   );
   gpc606_5 gpc191 (
      {stage0_17[102], stage0_17[103], stage0_17[104], stage0_17[105], stage0_17[106], stage0_17[107]},
      {stage0_19[90], stage0_19[91], stage0_19[92], stage0_19[93], stage0_19[94], stage0_19[95]},
      {stage1_21[15],stage1_20[30],stage1_19[32],stage1_18[33],stage1_17[52]}
   );
   gpc606_5 gpc192 (
      {stage0_17[108], stage0_17[109], stage0_17[110], stage0_17[111], stage0_17[112], stage0_17[113]},
      {stage0_19[96], stage0_19[97], stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101]},
      {stage1_21[16],stage1_20[31],stage1_19[33],stage1_18[34],stage1_17[53]}
   );
   gpc606_5 gpc193 (
      {stage0_17[114], stage0_17[115], stage0_17[116], stage0_17[117], stage0_17[118], stage0_17[119]},
      {stage0_19[102], stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage1_21[17],stage1_20[32],stage1_19[34],stage1_18[35],stage1_17[54]}
   );
   gpc615_5 gpc194 (
      {stage0_18[90], stage0_18[91], stage0_18[92], stage0_18[93], stage0_18[94]},
      {stage0_19[108]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[18],stage1_20[33],stage1_19[35],stage1_18[36]}
   );
   gpc615_5 gpc195 (
      {stage0_18[95], stage0_18[96], stage0_18[97], stage0_18[98], stage0_18[99]},
      {stage0_19[109]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[19],stage1_20[34],stage1_19[36],stage1_18[37]}
   );
   gpc615_5 gpc196 (
      {stage0_19[110], stage0_19[111], stage0_19[112], stage0_19[113], stage0_19[114]},
      {stage0_20[12]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[2],stage1_21[20],stage1_20[35],stage1_19[37]}
   );
   gpc615_5 gpc197 (
      {stage0_19[115], stage0_19[116], stage0_19[117], stage0_19[118], stage0_19[119]},
      {stage0_20[13]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[3],stage1_21[21],stage1_20[36],stage1_19[38]}
   );
   gpc615_5 gpc198 (
      {stage0_19[120], stage0_19[121], stage0_19[122], stage0_19[123], stage0_19[124]},
      {stage0_20[14]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[4],stage1_21[22],stage1_20[37],stage1_19[39]}
   );
   gpc606_5 gpc199 (
      {stage0_20[15], stage0_20[16], stage0_20[17], stage0_20[18], stage0_20[19], stage0_20[20]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[3],stage1_22[5],stage1_21[23],stage1_20[38]}
   );
   gpc606_5 gpc200 (
      {stage0_20[21], stage0_20[22], stage0_20[23], stage0_20[24], stage0_20[25], stage0_20[26]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[4],stage1_22[6],stage1_21[24],stage1_20[39]}
   );
   gpc606_5 gpc201 (
      {stage0_20[27], stage0_20[28], stage0_20[29], stage0_20[30], stage0_20[31], stage0_20[32]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[5],stage1_22[7],stage1_21[25],stage1_20[40]}
   );
   gpc606_5 gpc202 (
      {stage0_20[33], stage0_20[34], stage0_20[35], stage0_20[36], stage0_20[37], stage0_20[38]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[6],stage1_22[8],stage1_21[26],stage1_20[41]}
   );
   gpc606_5 gpc203 (
      {stage0_20[39], stage0_20[40], stage0_20[41], stage0_20[42], stage0_20[43], stage0_20[44]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[7],stage1_22[9],stage1_21[27],stage1_20[42]}
   );
   gpc606_5 gpc204 (
      {stage0_20[45], stage0_20[46], stage0_20[47], stage0_20[48], stage0_20[49], stage0_20[50]},
      {stage0_22[30], stage0_22[31], stage0_22[32], stage0_22[33], stage0_22[34], stage0_22[35]},
      {stage1_24[5],stage1_23[8],stage1_22[10],stage1_21[28],stage1_20[43]}
   );
   gpc606_5 gpc205 (
      {stage0_20[51], stage0_20[52], stage0_20[53], stage0_20[54], stage0_20[55], stage0_20[56]},
      {stage0_22[36], stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41]},
      {stage1_24[6],stage1_23[9],stage1_22[11],stage1_21[29],stage1_20[44]}
   );
   gpc606_5 gpc206 (
      {stage0_20[57], stage0_20[58], stage0_20[59], stage0_20[60], stage0_20[61], stage0_20[62]},
      {stage0_22[42], stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47]},
      {stage1_24[7],stage1_23[10],stage1_22[12],stage1_21[30],stage1_20[45]}
   );
   gpc606_5 gpc207 (
      {stage0_20[63], stage0_20[64], stage0_20[65], stage0_20[66], stage0_20[67], stage0_20[68]},
      {stage0_22[48], stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53]},
      {stage1_24[8],stage1_23[11],stage1_22[13],stage1_21[31],stage1_20[46]}
   );
   gpc606_5 gpc208 (
      {stage0_20[69], stage0_20[70], stage0_20[71], stage0_20[72], stage0_20[73], stage0_20[74]},
      {stage0_22[54], stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59]},
      {stage1_24[9],stage1_23[12],stage1_22[14],stage1_21[32],stage1_20[47]}
   );
   gpc606_5 gpc209 (
      {stage0_20[75], stage0_20[76], stage0_20[77], stage0_20[78], stage0_20[79], stage0_20[80]},
      {stage0_22[60], stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65]},
      {stage1_24[10],stage1_23[13],stage1_22[15],stage1_21[33],stage1_20[48]}
   );
   gpc606_5 gpc210 (
      {stage0_20[81], stage0_20[82], stage0_20[83], stage0_20[84], stage0_20[85], stage0_20[86]},
      {stage0_22[66], stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71]},
      {stage1_24[11],stage1_23[14],stage1_22[16],stage1_21[34],stage1_20[49]}
   );
   gpc606_5 gpc211 (
      {stage0_20[87], stage0_20[88], stage0_20[89], stage0_20[90], stage0_20[91], stage0_20[92]},
      {stage0_22[72], stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77]},
      {stage1_24[12],stage1_23[15],stage1_22[17],stage1_21[35],stage1_20[50]}
   );
   gpc606_5 gpc212 (
      {stage0_20[93], stage0_20[94], stage0_20[95], stage0_20[96], stage0_20[97], stage0_20[98]},
      {stage0_22[78], stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83]},
      {stage1_24[13],stage1_23[16],stage1_22[18],stage1_21[36],stage1_20[51]}
   );
   gpc606_5 gpc213 (
      {stage0_20[99], stage0_20[100], stage0_20[101], stage0_20[102], stage0_20[103], stage0_20[104]},
      {stage0_22[84], stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89]},
      {stage1_24[14],stage1_23[17],stage1_22[19],stage1_21[37],stage1_20[52]}
   );
   gpc606_5 gpc214 (
      {stage0_20[105], stage0_20[106], stage0_20[107], stage0_20[108], stage0_20[109], stage0_20[110]},
      {stage0_22[90], stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage1_24[15],stage1_23[18],stage1_22[20],stage1_21[38],stage1_20[53]}
   );
   gpc606_5 gpc215 (
      {stage0_20[111], stage0_20[112], stage0_20[113], stage0_20[114], stage0_20[115], stage0_20[116]},
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100], stage0_22[101]},
      {stage1_24[16],stage1_23[19],stage1_22[21],stage1_21[39],stage1_20[54]}
   );
   gpc606_5 gpc216 (
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[17],stage1_23[20],stage1_22[22],stage1_21[40]}
   );
   gpc606_5 gpc217 (
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[18],stage1_23[21],stage1_22[23],stage1_21[41]}
   );
   gpc606_5 gpc218 (
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[19],stage1_23[22],stage1_22[24],stage1_21[42]}
   );
   gpc606_5 gpc219 (
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[20],stage1_23[23],stage1_22[25],stage1_21[43]}
   );
   gpc606_5 gpc220 (
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[21],stage1_23[24],stage1_22[26],stage1_21[44]}
   );
   gpc606_5 gpc221 (
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[22],stage1_23[25],stage1_22[27],stage1_21[45]}
   );
   gpc606_5 gpc222 (
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59]},
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage1_25[6],stage1_24[23],stage1_23[26],stage1_22[28],stage1_21[46]}
   );
   gpc606_5 gpc223 (
      {stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65]},
      {stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage1_25[7],stage1_24[24],stage1_23[27],stage1_22[29],stage1_21[47]}
   );
   gpc606_5 gpc224 (
      {stage0_21[66], stage0_21[67], stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71]},
      {stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53]},
      {stage1_25[8],stage1_24[25],stage1_23[28],stage1_22[30],stage1_21[48]}
   );
   gpc606_5 gpc225 (
      {stage0_21[72], stage0_21[73], stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77]},
      {stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59]},
      {stage1_25[9],stage1_24[26],stage1_23[29],stage1_22[31],stage1_21[49]}
   );
   gpc606_5 gpc226 (
      {stage0_21[78], stage0_21[79], stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83]},
      {stage0_23[60], stage0_23[61], stage0_23[62], stage0_23[63], stage0_23[64], stage0_23[65]},
      {stage1_25[10],stage1_24[27],stage1_23[30],stage1_22[32],stage1_21[50]}
   );
   gpc606_5 gpc227 (
      {stage0_21[84], stage0_21[85], stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89]},
      {stage0_23[66], stage0_23[67], stage0_23[68], stage0_23[69], stage0_23[70], stage0_23[71]},
      {stage1_25[11],stage1_24[28],stage1_23[31],stage1_22[33],stage1_21[51]}
   );
   gpc606_5 gpc228 (
      {stage0_21[90], stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95]},
      {stage0_23[72], stage0_23[73], stage0_23[74], stage0_23[75], stage0_23[76], stage0_23[77]},
      {stage1_25[12],stage1_24[29],stage1_23[32],stage1_22[34],stage1_21[52]}
   );
   gpc606_5 gpc229 (
      {stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100], stage0_21[101]},
      {stage0_23[78], stage0_23[79], stage0_23[80], stage0_23[81], stage0_23[82], stage0_23[83]},
      {stage1_25[13],stage1_24[30],stage1_23[33],stage1_22[35],stage1_21[53]}
   );
   gpc606_5 gpc230 (
      {stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105], stage0_21[106], stage0_21[107]},
      {stage0_23[84], stage0_23[85], stage0_23[86], stage0_23[87], stage0_23[88], stage0_23[89]},
      {stage1_25[14],stage1_24[31],stage1_23[34],stage1_22[36],stage1_21[54]}
   );
   gpc606_5 gpc231 (
      {stage0_21[108], stage0_21[109], stage0_21[110], stage0_21[111], stage0_21[112], stage0_21[113]},
      {stage0_23[90], stage0_23[91], stage0_23[92], stage0_23[93], stage0_23[94], stage0_23[95]},
      {stage1_25[15],stage1_24[32],stage1_23[35],stage1_22[37],stage1_21[55]}
   );
   gpc606_5 gpc232 (
      {stage0_21[114], stage0_21[115], stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119]},
      {stage0_23[96], stage0_23[97], stage0_23[98], stage0_23[99], stage0_23[100], stage0_23[101]},
      {stage1_25[16],stage1_24[33],stage1_23[36],stage1_22[38],stage1_21[56]}
   );
   gpc615_5 gpc233 (
      {stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105], stage0_22[106]},
      {stage0_23[102]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[17],stage1_24[34],stage1_23[37],stage1_22[39]}
   );
   gpc606_5 gpc234 (
      {stage0_23[103], stage0_23[104], stage0_23[105], stage0_23[106], stage0_23[107], stage0_23[108]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[1],stage1_25[18],stage1_24[35],stage1_23[38]}
   );
   gpc606_5 gpc235 (
      {stage0_23[109], stage0_23[110], stage0_23[111], stage0_23[112], stage0_23[113], stage0_23[114]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[2],stage1_25[19],stage1_24[36],stage1_23[39]}
   );
   gpc606_5 gpc236 (
      {stage0_23[115], stage0_23[116], stage0_23[117], stage0_23[118], stage0_23[119], stage0_23[120]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[3],stage1_25[20],stage1_24[37],stage1_23[40]}
   );
   gpc615_5 gpc237 (
      {stage0_23[121], stage0_23[122], stage0_23[123], stage0_23[124], stage0_23[125]},
      {stage0_24[6]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[4],stage1_25[21],stage1_24[38],stage1_23[41]}
   );
   gpc606_5 gpc238 (
      {stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11], stage0_24[12]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[4],stage1_26[5],stage1_25[22],stage1_24[39]}
   );
   gpc606_5 gpc239 (
      {stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17], stage0_24[18]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[5],stage1_26[6],stage1_25[23],stage1_24[40]}
   );
   gpc606_5 gpc240 (
      {stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23], stage0_24[24]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[6],stage1_26[7],stage1_25[24],stage1_24[41]}
   );
   gpc606_5 gpc241 (
      {stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29], stage0_24[30]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[7],stage1_26[8],stage1_25[25],stage1_24[42]}
   );
   gpc606_5 gpc242 (
      {stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35], stage0_24[36]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[8],stage1_26[9],stage1_25[26],stage1_24[43]}
   );
   gpc606_5 gpc243 (
      {stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41], stage0_24[42]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[9],stage1_26[10],stage1_25[27],stage1_24[44]}
   );
   gpc606_5 gpc244 (
      {stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47], stage0_24[48]},
      {stage0_26[36], stage0_26[37], stage0_26[38], stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage1_28[6],stage1_27[10],stage1_26[11],stage1_25[28],stage1_24[45]}
   );
   gpc606_5 gpc245 (
      {stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53], stage0_24[54]},
      {stage0_26[42], stage0_26[43], stage0_26[44], stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage1_28[7],stage1_27[11],stage1_26[12],stage1_25[29],stage1_24[46]}
   );
   gpc606_5 gpc246 (
      {stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59], stage0_24[60]},
      {stage0_26[48], stage0_26[49], stage0_26[50], stage0_26[51], stage0_26[52], stage0_26[53]},
      {stage1_28[8],stage1_27[12],stage1_26[13],stage1_25[30],stage1_24[47]}
   );
   gpc606_5 gpc247 (
      {stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65], stage0_24[66]},
      {stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57], stage0_26[58], stage0_26[59]},
      {stage1_28[9],stage1_27[13],stage1_26[14],stage1_25[31],stage1_24[48]}
   );
   gpc606_5 gpc248 (
      {stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71], stage0_24[72]},
      {stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63], stage0_26[64], stage0_26[65]},
      {stage1_28[10],stage1_27[14],stage1_26[15],stage1_25[32],stage1_24[49]}
   );
   gpc606_5 gpc249 (
      {stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77], stage0_24[78]},
      {stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69], stage0_26[70], stage0_26[71]},
      {stage1_28[11],stage1_27[15],stage1_26[16],stage1_25[33],stage1_24[50]}
   );
   gpc606_5 gpc250 (
      {stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83], stage0_24[84]},
      {stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75], stage0_26[76], stage0_26[77]},
      {stage1_28[12],stage1_27[16],stage1_26[17],stage1_25[34],stage1_24[51]}
   );
   gpc606_5 gpc251 (
      {stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89], stage0_24[90]},
      {stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81], stage0_26[82], stage0_26[83]},
      {stage1_28[13],stage1_27[17],stage1_26[18],stage1_25[35],stage1_24[52]}
   );
   gpc606_5 gpc252 (
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[14],stage1_27[18],stage1_26[19],stage1_25[36]}
   );
   gpc606_5 gpc253 (
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[15],stage1_27[19],stage1_26[20],stage1_25[37]}
   );
   gpc606_5 gpc254 (
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[16],stage1_27[20],stage1_26[21],stage1_25[38]}
   );
   gpc606_5 gpc255 (
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[17],stage1_27[21],stage1_26[22],stage1_25[39]}
   );
   gpc606_5 gpc256 (
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[18],stage1_27[22],stage1_26[23],stage1_25[40]}
   );
   gpc606_5 gpc257 (
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[19],stage1_27[23],stage1_26[24],stage1_25[41]}
   );
   gpc606_5 gpc258 (
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[20],stage1_27[24],stage1_26[25],stage1_25[42]}
   );
   gpc606_5 gpc259 (
      {stage0_25[66], stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[21],stage1_27[25],stage1_26[26],stage1_25[43]}
   );
   gpc606_5 gpc260 (
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[22],stage1_27[26],stage1_26[27],stage1_25[44]}
   );
   gpc606_5 gpc261 (
      {stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage1_29[9],stage1_28[23],stage1_27[27],stage1_26[28],stage1_25[45]}
   );
   gpc606_5 gpc262 (
      {stage0_25[84], stage0_25[85], stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage1_29[10],stage1_28[24],stage1_27[28],stage1_26[29],stage1_25[46]}
   );
   gpc606_5 gpc263 (
      {stage0_25[90], stage0_25[91], stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage1_29[11],stage1_28[25],stage1_27[29],stage1_26[30],stage1_25[47]}
   );
   gpc606_5 gpc264 (
      {stage0_25[96], stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage1_29[12],stage1_28[26],stage1_27[30],stage1_26[31],stage1_25[48]}
   );
   gpc606_5 gpc265 (
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage1_29[13],stage1_28[27],stage1_27[31],stage1_26[32],stage1_25[49]}
   );
   gpc615_5 gpc266 (
      {stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87], stage0_26[88]},
      {stage0_27[84]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[14],stage1_28[28],stage1_27[32],stage1_26[33]}
   );
   gpc615_5 gpc267 (
      {stage0_26[89], stage0_26[90], stage0_26[91], stage0_26[92], stage0_26[93]},
      {stage0_27[85]},
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage1_30[1],stage1_29[15],stage1_28[29],stage1_27[33],stage1_26[34]}
   );
   gpc615_5 gpc268 (
      {stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89], stage0_27[90]},
      {stage0_28[12]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[2],stage1_29[16],stage1_28[30],stage1_27[34]}
   );
   gpc615_5 gpc269 (
      {stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage0_28[13]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[3],stage1_29[17],stage1_28[31],stage1_27[35]}
   );
   gpc615_5 gpc270 (
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100]},
      {stage0_28[14]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[4],stage1_29[18],stage1_28[32],stage1_27[36]}
   );
   gpc615_5 gpc271 (
      {stage0_27[101], stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105]},
      {stage0_28[15]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[5],stage1_29[19],stage1_28[33],stage1_27[37]}
   );
   gpc615_5 gpc272 (
      {stage0_27[106], stage0_27[107], stage0_27[108], stage0_27[109], stage0_27[110]},
      {stage0_28[16]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[6],stage1_29[20],stage1_28[34],stage1_27[38]}
   );
   gpc606_5 gpc273 (
      {stage0_28[17], stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[5],stage1_30[7],stage1_29[21],stage1_28[35]}
   );
   gpc606_5 gpc274 (
      {stage0_28[23], stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[6],stage1_30[8],stage1_29[22],stage1_28[36]}
   );
   gpc606_5 gpc275 (
      {stage0_28[29], stage0_28[30], stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[7],stage1_30[9],stage1_29[23],stage1_28[37]}
   );
   gpc606_5 gpc276 (
      {stage0_28[35], stage0_28[36], stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[8],stage1_30[10],stage1_29[24],stage1_28[38]}
   );
   gpc606_5 gpc277 (
      {stage0_28[41], stage0_28[42], stage0_28[43], stage0_28[44], stage0_28[45], stage0_28[46]},
      {stage0_30[24], stage0_30[25], stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29]},
      {stage1_32[4],stage1_31[9],stage1_30[11],stage1_29[25],stage1_28[39]}
   );
   gpc606_5 gpc278 (
      {stage0_28[47], stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51], stage0_28[52]},
      {stage0_30[30], stage0_30[31], stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35]},
      {stage1_32[5],stage1_31[10],stage1_30[12],stage1_29[26],stage1_28[40]}
   );
   gpc606_5 gpc279 (
      {stage0_28[53], stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57], stage0_28[58]},
      {stage0_30[36], stage0_30[37], stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41]},
      {stage1_32[6],stage1_31[11],stage1_30[13],stage1_29[27],stage1_28[41]}
   );
   gpc606_5 gpc280 (
      {stage0_28[59], stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63], stage0_28[64]},
      {stage0_30[42], stage0_30[43], stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47]},
      {stage1_32[7],stage1_31[12],stage1_30[14],stage1_29[28],stage1_28[42]}
   );
   gpc606_5 gpc281 (
      {stage0_28[65], stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69], stage0_28[70]},
      {stage0_30[48], stage0_30[49], stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53]},
      {stage1_32[8],stage1_31[13],stage1_30[15],stage1_29[29],stage1_28[43]}
   );
   gpc606_5 gpc282 (
      {stage0_28[71], stage0_28[72], stage0_28[73], stage0_28[74], stage0_28[75], stage0_28[76]},
      {stage0_30[54], stage0_30[55], stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59]},
      {stage1_32[9],stage1_31[14],stage1_30[16],stage1_29[30],stage1_28[44]}
   );
   gpc606_5 gpc283 (
      {stage0_28[77], stage0_28[78], stage0_28[79], stage0_28[80], stage0_28[81], stage0_28[82]},
      {stage0_30[60], stage0_30[61], stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65]},
      {stage1_32[10],stage1_31[15],stage1_30[17],stage1_29[31],stage1_28[45]}
   );
   gpc606_5 gpc284 (
      {stage0_28[83], stage0_28[84], stage0_28[85], stage0_28[86], stage0_28[87], stage0_28[88]},
      {stage0_30[66], stage0_30[67], stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71]},
      {stage1_32[11],stage1_31[16],stage1_30[18],stage1_29[32],stage1_28[46]}
   );
   gpc606_5 gpc285 (
      {stage0_28[89], stage0_28[90], stage0_28[91], stage0_28[92], stage0_28[93], stage0_28[94]},
      {stage0_30[72], stage0_30[73], stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77]},
      {stage1_32[12],stage1_31[17],stage1_30[19],stage1_29[33],stage1_28[47]}
   );
   gpc606_5 gpc286 (
      {stage0_28[95], stage0_28[96], stage0_28[97], stage0_28[98], stage0_28[99], stage0_28[100]},
      {stage0_30[78], stage0_30[79], stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83]},
      {stage1_32[13],stage1_31[18],stage1_30[20],stage1_29[34],stage1_28[48]}
   );
   gpc606_5 gpc287 (
      {stage0_28[101], stage0_28[102], stage0_28[103], stage0_28[104], stage0_28[105], stage0_28[106]},
      {stage0_30[84], stage0_30[85], stage0_30[86], stage0_30[87], stage0_30[88], stage0_30[89]},
      {stage1_32[14],stage1_31[19],stage1_30[21],stage1_29[35],stage1_28[49]}
   );
   gpc606_5 gpc288 (
      {stage0_28[107], stage0_28[108], stage0_28[109], stage0_28[110], stage0_28[111], stage0_28[112]},
      {stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93], stage0_30[94], stage0_30[95]},
      {stage1_32[15],stage1_31[20],stage1_30[22],stage1_29[36],stage1_28[50]}
   );
   gpc606_5 gpc289 (
      {stage0_28[113], stage0_28[114], stage0_28[115], stage0_28[116], stage0_28[117], stage0_28[118]},
      {stage0_30[96], stage0_30[97], stage0_30[98], stage0_30[99], stage0_30[100], stage0_30[101]},
      {stage1_32[16],stage1_31[21],stage1_30[23],stage1_29[37],stage1_28[51]}
   );
   gpc606_5 gpc290 (
      {stage0_28[119], stage0_28[120], stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124]},
      {stage0_30[102], stage0_30[103], stage0_30[104], stage0_30[105], stage0_30[106], stage0_30[107]},
      {stage1_32[17],stage1_31[22],stage1_30[24],stage1_29[38],stage1_28[52]}
   );
   gpc606_5 gpc291 (
      {stage0_29[30], stage0_29[31], stage0_29[32], stage0_29[33], stage0_29[34], stage0_29[35]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[18],stage1_31[23],stage1_30[25],stage1_29[39]}
   );
   gpc606_5 gpc292 (
      {stage0_29[36], stage0_29[37], stage0_29[38], stage0_29[39], stage0_29[40], stage0_29[41]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[19],stage1_31[24],stage1_30[26],stage1_29[40]}
   );
   gpc606_5 gpc293 (
      {stage0_29[42], stage0_29[43], stage0_29[44], stage0_29[45], stage0_29[46], stage0_29[47]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[20],stage1_31[25],stage1_30[27],stage1_29[41]}
   );
   gpc606_5 gpc294 (
      {stage0_29[48], stage0_29[49], stage0_29[50], stage0_29[51], stage0_29[52], stage0_29[53]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[21],stage1_31[26],stage1_30[28],stage1_29[42]}
   );
   gpc606_5 gpc295 (
      {stage0_29[54], stage0_29[55], stage0_29[56], stage0_29[57], stage0_29[58], stage0_29[59]},
      {stage0_31[24], stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29]},
      {stage1_33[4],stage1_32[22],stage1_31[27],stage1_30[29],stage1_29[43]}
   );
   gpc606_5 gpc296 (
      {stage0_29[60], stage0_29[61], stage0_29[62], stage0_29[63], stage0_29[64], stage0_29[65]},
      {stage0_31[30], stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35]},
      {stage1_33[5],stage1_32[23],stage1_31[28],stage1_30[30],stage1_29[44]}
   );
   gpc606_5 gpc297 (
      {stage0_29[66], stage0_29[67], stage0_29[68], stage0_29[69], stage0_29[70], stage0_29[71]},
      {stage0_31[36], stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41]},
      {stage1_33[6],stage1_32[24],stage1_31[29],stage1_30[31],stage1_29[45]}
   );
   gpc606_5 gpc298 (
      {stage0_29[72], stage0_29[73], stage0_29[74], stage0_29[75], stage0_29[76], stage0_29[77]},
      {stage0_31[42], stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47]},
      {stage1_33[7],stage1_32[25],stage1_31[30],stage1_30[32],stage1_29[46]}
   );
   gpc606_5 gpc299 (
      {stage0_29[78], stage0_29[79], stage0_29[80], stage0_29[81], stage0_29[82], stage0_29[83]},
      {stage0_31[48], stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53]},
      {stage1_33[8],stage1_32[26],stage1_31[31],stage1_30[33],stage1_29[47]}
   );
   gpc606_5 gpc300 (
      {stage0_29[84], stage0_29[85], stage0_29[86], stage0_29[87], stage0_29[88], stage0_29[89]},
      {stage0_31[54], stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59]},
      {stage1_33[9],stage1_32[27],stage1_31[32],stage1_30[34],stage1_29[48]}
   );
   gpc606_5 gpc301 (
      {stage0_29[90], stage0_29[91], stage0_29[92], stage0_29[93], stage0_29[94], stage0_29[95]},
      {stage0_31[60], stage0_31[61], stage0_31[62], stage0_31[63], stage0_31[64], stage0_31[65]},
      {stage1_33[10],stage1_32[28],stage1_31[33],stage1_30[35],stage1_29[49]}
   );
   gpc606_5 gpc302 (
      {stage0_29[96], stage0_29[97], stage0_29[98], stage0_29[99], stage0_29[100], stage0_29[101]},
      {stage0_31[66], stage0_31[67], stage0_31[68], stage0_31[69], stage0_31[70], stage0_31[71]},
      {stage1_33[11],stage1_32[29],stage1_31[34],stage1_30[36],stage1_29[50]}
   );
   gpc606_5 gpc303 (
      {stage0_29[102], stage0_29[103], stage0_29[104], stage0_29[105], stage0_29[106], stage0_29[107]},
      {stage0_31[72], stage0_31[73], stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77]},
      {stage1_33[12],stage1_32[30],stage1_31[35],stage1_30[37],stage1_29[51]}
   );
   gpc606_5 gpc304 (
      {stage0_29[108], stage0_29[109], stage0_29[110], stage0_29[111], stage0_29[112], stage0_29[113]},
      {stage0_31[78], stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage1_33[13],stage1_32[31],stage1_31[36],stage1_30[38],stage1_29[52]}
   );
   gpc606_5 gpc305 (
      {stage0_29[114], stage0_29[115], stage0_29[116], stage0_29[117], stage0_29[118], stage0_29[119]},
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88], stage0_31[89]},
      {stage1_33[14],stage1_32[32],stage1_31[37],stage1_30[39],stage1_29[53]}
   );
   gpc606_5 gpc306 (
      {stage0_29[120], stage0_29[121], stage0_29[122], stage0_29[123], stage0_29[124], stage0_29[125]},
      {stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93], stage0_31[94], stage0_31[95]},
      {stage1_33[15],stage1_32[33],stage1_31[38],stage1_30[40],stage1_29[54]}
   );
   gpc1_1 gpc307 (
      {stage0_0[116]},
      {stage1_0[24]}
   );
   gpc1_1 gpc308 (
      {stage0_0[117]},
      {stage1_0[25]}
   );
   gpc1_1 gpc309 (
      {stage0_0[118]},
      {stage1_0[26]}
   );
   gpc1_1 gpc310 (
      {stage0_0[119]},
      {stage1_0[27]}
   );
   gpc1_1 gpc311 (
      {stage0_0[120]},
      {stage1_0[28]}
   );
   gpc1_1 gpc312 (
      {stage0_0[121]},
      {stage1_0[29]}
   );
   gpc1_1 gpc313 (
      {stage0_0[122]},
      {stage1_0[30]}
   );
   gpc1_1 gpc314 (
      {stage0_0[123]},
      {stage1_0[31]}
   );
   gpc1_1 gpc315 (
      {stage0_0[124]},
      {stage1_0[32]}
   );
   gpc1_1 gpc316 (
      {stage0_0[125]},
      {stage1_0[33]}
   );
   gpc1_1 gpc317 (
      {stage0_0[126]},
      {stage1_0[34]}
   );
   gpc1_1 gpc318 (
      {stage0_0[127]},
      {stage1_0[35]}
   );
   gpc1_1 gpc319 (
      {stage0_1[124]},
      {stage1_1[36]}
   );
   gpc1_1 gpc320 (
      {stage0_1[125]},
      {stage1_1[37]}
   );
   gpc1_1 gpc321 (
      {stage0_1[126]},
      {stage1_1[38]}
   );
   gpc1_1 gpc322 (
      {stage0_1[127]},
      {stage1_1[39]}
   );
   gpc1_1 gpc323 (
      {stage0_2[107]},
      {stage1_2[37]}
   );
   gpc1_1 gpc324 (
      {stage0_2[108]},
      {stage1_2[38]}
   );
   gpc1_1 gpc325 (
      {stage0_2[109]},
      {stage1_2[39]}
   );
   gpc1_1 gpc326 (
      {stage0_2[110]},
      {stage1_2[40]}
   );
   gpc1_1 gpc327 (
      {stage0_2[111]},
      {stage1_2[41]}
   );
   gpc1_1 gpc328 (
      {stage0_2[112]},
      {stage1_2[42]}
   );
   gpc1_1 gpc329 (
      {stage0_2[113]},
      {stage1_2[43]}
   );
   gpc1_1 gpc330 (
      {stage0_2[114]},
      {stage1_2[44]}
   );
   gpc1_1 gpc331 (
      {stage0_2[115]},
      {stage1_2[45]}
   );
   gpc1_1 gpc332 (
      {stage0_2[116]},
      {stage1_2[46]}
   );
   gpc1_1 gpc333 (
      {stage0_2[117]},
      {stage1_2[47]}
   );
   gpc1_1 gpc334 (
      {stage0_2[118]},
      {stage1_2[48]}
   );
   gpc1_1 gpc335 (
      {stage0_2[119]},
      {stage1_2[49]}
   );
   gpc1_1 gpc336 (
      {stage0_2[120]},
      {stage1_2[50]}
   );
   gpc1_1 gpc337 (
      {stage0_2[121]},
      {stage1_2[51]}
   );
   gpc1_1 gpc338 (
      {stage0_2[122]},
      {stage1_2[52]}
   );
   gpc1_1 gpc339 (
      {stage0_2[123]},
      {stage1_2[53]}
   );
   gpc1_1 gpc340 (
      {stage0_2[124]},
      {stage1_2[54]}
   );
   gpc1_1 gpc341 (
      {stage0_2[125]},
      {stage1_2[55]}
   );
   gpc1_1 gpc342 (
      {stage0_2[126]},
      {stage1_2[56]}
   );
   gpc1_1 gpc343 (
      {stage0_2[127]},
      {stage1_2[57]}
   );
   gpc1_1 gpc344 (
      {stage0_3[112]},
      {stage1_3[43]}
   );
   gpc1_1 gpc345 (
      {stage0_3[113]},
      {stage1_3[44]}
   );
   gpc1_1 gpc346 (
      {stage0_3[114]},
      {stage1_3[45]}
   );
   gpc1_1 gpc347 (
      {stage0_3[115]},
      {stage1_3[46]}
   );
   gpc1_1 gpc348 (
      {stage0_3[116]},
      {stage1_3[47]}
   );
   gpc1_1 gpc349 (
      {stage0_3[117]},
      {stage1_3[48]}
   );
   gpc1_1 gpc350 (
      {stage0_3[118]},
      {stage1_3[49]}
   );
   gpc1_1 gpc351 (
      {stage0_3[119]},
      {stage1_3[50]}
   );
   gpc1_1 gpc352 (
      {stage0_3[120]},
      {stage1_3[51]}
   );
   gpc1_1 gpc353 (
      {stage0_3[121]},
      {stage1_3[52]}
   );
   gpc1_1 gpc354 (
      {stage0_3[122]},
      {stage1_3[53]}
   );
   gpc1_1 gpc355 (
      {stage0_3[123]},
      {stage1_3[54]}
   );
   gpc1_1 gpc356 (
      {stage0_3[124]},
      {stage1_3[55]}
   );
   gpc1_1 gpc357 (
      {stage0_3[125]},
      {stage1_3[56]}
   );
   gpc1_1 gpc358 (
      {stage0_3[126]},
      {stage1_3[57]}
   );
   gpc1_1 gpc359 (
      {stage0_3[127]},
      {stage1_3[58]}
   );
   gpc1_1 gpc360 (
      {stage0_4[122]},
      {stage1_4[61]}
   );
   gpc1_1 gpc361 (
      {stage0_4[123]},
      {stage1_4[62]}
   );
   gpc1_1 gpc362 (
      {stage0_4[124]},
      {stage1_4[63]}
   );
   gpc1_1 gpc363 (
      {stage0_4[125]},
      {stage1_4[64]}
   );
   gpc1_1 gpc364 (
      {stage0_4[126]},
      {stage1_4[65]}
   );
   gpc1_1 gpc365 (
      {stage0_4[127]},
      {stage1_4[66]}
   );
   gpc1_1 gpc366 (
      {stage0_5[116]},
      {stage1_5[51]}
   );
   gpc1_1 gpc367 (
      {stage0_5[117]},
      {stage1_5[52]}
   );
   gpc1_1 gpc368 (
      {stage0_5[118]},
      {stage1_5[53]}
   );
   gpc1_1 gpc369 (
      {stage0_5[119]},
      {stage1_5[54]}
   );
   gpc1_1 gpc370 (
      {stage0_5[120]},
      {stage1_5[55]}
   );
   gpc1_1 gpc371 (
      {stage0_5[121]},
      {stage1_5[56]}
   );
   gpc1_1 gpc372 (
      {stage0_5[122]},
      {stage1_5[57]}
   );
   gpc1_1 gpc373 (
      {stage0_5[123]},
      {stage1_5[58]}
   );
   gpc1_1 gpc374 (
      {stage0_5[124]},
      {stage1_5[59]}
   );
   gpc1_1 gpc375 (
      {stage0_5[125]},
      {stage1_5[60]}
   );
   gpc1_1 gpc376 (
      {stage0_5[126]},
      {stage1_5[61]}
   );
   gpc1_1 gpc377 (
      {stage0_5[127]},
      {stage1_5[62]}
   );
   gpc1_1 gpc378 (
      {stage0_6[119]},
      {stage1_6[41]}
   );
   gpc1_1 gpc379 (
      {stage0_6[120]},
      {stage1_6[42]}
   );
   gpc1_1 gpc380 (
      {stage0_6[121]},
      {stage1_6[43]}
   );
   gpc1_1 gpc381 (
      {stage0_6[122]},
      {stage1_6[44]}
   );
   gpc1_1 gpc382 (
      {stage0_6[123]},
      {stage1_6[45]}
   );
   gpc1_1 gpc383 (
      {stage0_6[124]},
      {stage1_6[46]}
   );
   gpc1_1 gpc384 (
      {stage0_6[125]},
      {stage1_6[47]}
   );
   gpc1_1 gpc385 (
      {stage0_6[126]},
      {stage1_6[48]}
   );
   gpc1_1 gpc386 (
      {stage0_6[127]},
      {stage1_6[49]}
   );
   gpc1_1 gpc387 (
      {stage0_7[101]},
      {stage1_7[43]}
   );
   gpc1_1 gpc388 (
      {stage0_7[102]},
      {stage1_7[44]}
   );
   gpc1_1 gpc389 (
      {stage0_7[103]},
      {stage1_7[45]}
   );
   gpc1_1 gpc390 (
      {stage0_7[104]},
      {stage1_7[46]}
   );
   gpc1_1 gpc391 (
      {stage0_7[105]},
      {stage1_7[47]}
   );
   gpc1_1 gpc392 (
      {stage0_7[106]},
      {stage1_7[48]}
   );
   gpc1_1 gpc393 (
      {stage0_7[107]},
      {stage1_7[49]}
   );
   gpc1_1 gpc394 (
      {stage0_7[108]},
      {stage1_7[50]}
   );
   gpc1_1 gpc395 (
      {stage0_7[109]},
      {stage1_7[51]}
   );
   gpc1_1 gpc396 (
      {stage0_7[110]},
      {stage1_7[52]}
   );
   gpc1_1 gpc397 (
      {stage0_7[111]},
      {stage1_7[53]}
   );
   gpc1_1 gpc398 (
      {stage0_7[112]},
      {stage1_7[54]}
   );
   gpc1_1 gpc399 (
      {stage0_7[113]},
      {stage1_7[55]}
   );
   gpc1_1 gpc400 (
      {stage0_7[114]},
      {stage1_7[56]}
   );
   gpc1_1 gpc401 (
      {stage0_7[115]},
      {stage1_7[57]}
   );
   gpc1_1 gpc402 (
      {stage0_7[116]},
      {stage1_7[58]}
   );
   gpc1_1 gpc403 (
      {stage0_7[117]},
      {stage1_7[59]}
   );
   gpc1_1 gpc404 (
      {stage0_7[118]},
      {stage1_7[60]}
   );
   gpc1_1 gpc405 (
      {stage0_7[119]},
      {stage1_7[61]}
   );
   gpc1_1 gpc406 (
      {stage0_7[120]},
      {stage1_7[62]}
   );
   gpc1_1 gpc407 (
      {stage0_7[121]},
      {stage1_7[63]}
   );
   gpc1_1 gpc408 (
      {stage0_7[122]},
      {stage1_7[64]}
   );
   gpc1_1 gpc409 (
      {stage0_7[123]},
      {stage1_7[65]}
   );
   gpc1_1 gpc410 (
      {stage0_7[124]},
      {stage1_7[66]}
   );
   gpc1_1 gpc411 (
      {stage0_7[125]},
      {stage1_7[67]}
   );
   gpc1_1 gpc412 (
      {stage0_7[126]},
      {stage1_7[68]}
   );
   gpc1_1 gpc413 (
      {stage0_7[127]},
      {stage1_7[69]}
   );
   gpc1_1 gpc414 (
      {stage0_9[122]},
      {stage1_9[55]}
   );
   gpc1_1 gpc415 (
      {stage0_9[123]},
      {stage1_9[56]}
   );
   gpc1_1 gpc416 (
      {stage0_9[124]},
      {stage1_9[57]}
   );
   gpc1_1 gpc417 (
      {stage0_9[125]},
      {stage1_9[58]}
   );
   gpc1_1 gpc418 (
      {stage0_9[126]},
      {stage1_9[59]}
   );
   gpc1_1 gpc419 (
      {stage0_9[127]},
      {stage1_9[60]}
   );
   gpc1_1 gpc420 (
      {stage0_10[116]},
      {stage1_10[42]}
   );
   gpc1_1 gpc421 (
      {stage0_10[117]},
      {stage1_10[43]}
   );
   gpc1_1 gpc422 (
      {stage0_10[118]},
      {stage1_10[44]}
   );
   gpc1_1 gpc423 (
      {stage0_10[119]},
      {stage1_10[45]}
   );
   gpc1_1 gpc424 (
      {stage0_10[120]},
      {stage1_10[46]}
   );
   gpc1_1 gpc425 (
      {stage0_10[121]},
      {stage1_10[47]}
   );
   gpc1_1 gpc426 (
      {stage0_10[122]},
      {stage1_10[48]}
   );
   gpc1_1 gpc427 (
      {stage0_10[123]},
      {stage1_10[49]}
   );
   gpc1_1 gpc428 (
      {stage0_10[124]},
      {stage1_10[50]}
   );
   gpc1_1 gpc429 (
      {stage0_10[125]},
      {stage1_10[51]}
   );
   gpc1_1 gpc430 (
      {stage0_10[126]},
      {stage1_10[52]}
   );
   gpc1_1 gpc431 (
      {stage0_10[127]},
      {stage1_10[53]}
   );
   gpc1_1 gpc432 (
      {stage0_11[112]},
      {stage1_11[42]}
   );
   gpc1_1 gpc433 (
      {stage0_11[113]},
      {stage1_11[43]}
   );
   gpc1_1 gpc434 (
      {stage0_11[114]},
      {stage1_11[44]}
   );
   gpc1_1 gpc435 (
      {stage0_11[115]},
      {stage1_11[45]}
   );
   gpc1_1 gpc436 (
      {stage0_11[116]},
      {stage1_11[46]}
   );
   gpc1_1 gpc437 (
      {stage0_11[117]},
      {stage1_11[47]}
   );
   gpc1_1 gpc438 (
      {stage0_11[118]},
      {stage1_11[48]}
   );
   gpc1_1 gpc439 (
      {stage0_11[119]},
      {stage1_11[49]}
   );
   gpc1_1 gpc440 (
      {stage0_11[120]},
      {stage1_11[50]}
   );
   gpc1_1 gpc441 (
      {stage0_11[121]},
      {stage1_11[51]}
   );
   gpc1_1 gpc442 (
      {stage0_11[122]},
      {stage1_11[52]}
   );
   gpc1_1 gpc443 (
      {stage0_11[123]},
      {stage1_11[53]}
   );
   gpc1_1 gpc444 (
      {stage0_11[124]},
      {stage1_11[54]}
   );
   gpc1_1 gpc445 (
      {stage0_11[125]},
      {stage1_11[55]}
   );
   gpc1_1 gpc446 (
      {stage0_11[126]},
      {stage1_11[56]}
   );
   gpc1_1 gpc447 (
      {stage0_11[127]},
      {stage1_11[57]}
   );
   gpc1_1 gpc448 (
      {stage0_13[126]},
      {stage1_13[59]}
   );
   gpc1_1 gpc449 (
      {stage0_13[127]},
      {stage1_13[60]}
   );
   gpc1_1 gpc450 (
      {stage0_14[125]},
      {stage1_14[43]}
   );
   gpc1_1 gpc451 (
      {stage0_14[126]},
      {stage1_14[44]}
   );
   gpc1_1 gpc452 (
      {stage0_14[127]},
      {stage1_14[45]}
   );
   gpc1_1 gpc453 (
      {stage0_15[125]},
      {stage1_15[44]}
   );
   gpc1_1 gpc454 (
      {stage0_15[126]},
      {stage1_15[45]}
   );
   gpc1_1 gpc455 (
      {stage0_15[127]},
      {stage1_15[46]}
   );
   gpc1_1 gpc456 (
      {stage0_16[98]},
      {stage1_16[57]}
   );
   gpc1_1 gpc457 (
      {stage0_16[99]},
      {stage1_16[58]}
   );
   gpc1_1 gpc458 (
      {stage0_16[100]},
      {stage1_16[59]}
   );
   gpc1_1 gpc459 (
      {stage0_16[101]},
      {stage1_16[60]}
   );
   gpc1_1 gpc460 (
      {stage0_16[102]},
      {stage1_16[61]}
   );
   gpc1_1 gpc461 (
      {stage0_16[103]},
      {stage1_16[62]}
   );
   gpc1_1 gpc462 (
      {stage0_16[104]},
      {stage1_16[63]}
   );
   gpc1_1 gpc463 (
      {stage0_16[105]},
      {stage1_16[64]}
   );
   gpc1_1 gpc464 (
      {stage0_16[106]},
      {stage1_16[65]}
   );
   gpc1_1 gpc465 (
      {stage0_16[107]},
      {stage1_16[66]}
   );
   gpc1_1 gpc466 (
      {stage0_16[108]},
      {stage1_16[67]}
   );
   gpc1_1 gpc467 (
      {stage0_16[109]},
      {stage1_16[68]}
   );
   gpc1_1 gpc468 (
      {stage0_16[110]},
      {stage1_16[69]}
   );
   gpc1_1 gpc469 (
      {stage0_16[111]},
      {stage1_16[70]}
   );
   gpc1_1 gpc470 (
      {stage0_16[112]},
      {stage1_16[71]}
   );
   gpc1_1 gpc471 (
      {stage0_16[113]},
      {stage1_16[72]}
   );
   gpc1_1 gpc472 (
      {stage0_16[114]},
      {stage1_16[73]}
   );
   gpc1_1 gpc473 (
      {stage0_16[115]},
      {stage1_16[74]}
   );
   gpc1_1 gpc474 (
      {stage0_16[116]},
      {stage1_16[75]}
   );
   gpc1_1 gpc475 (
      {stage0_16[117]},
      {stage1_16[76]}
   );
   gpc1_1 gpc476 (
      {stage0_16[118]},
      {stage1_16[77]}
   );
   gpc1_1 gpc477 (
      {stage0_16[119]},
      {stage1_16[78]}
   );
   gpc1_1 gpc478 (
      {stage0_16[120]},
      {stage1_16[79]}
   );
   gpc1_1 gpc479 (
      {stage0_16[121]},
      {stage1_16[80]}
   );
   gpc1_1 gpc480 (
      {stage0_16[122]},
      {stage1_16[81]}
   );
   gpc1_1 gpc481 (
      {stage0_16[123]},
      {stage1_16[82]}
   );
   gpc1_1 gpc482 (
      {stage0_16[124]},
      {stage1_16[83]}
   );
   gpc1_1 gpc483 (
      {stage0_16[125]},
      {stage1_16[84]}
   );
   gpc1_1 gpc484 (
      {stage0_16[126]},
      {stage1_16[85]}
   );
   gpc1_1 gpc485 (
      {stage0_16[127]},
      {stage1_16[86]}
   );
   gpc1_1 gpc486 (
      {stage0_17[120]},
      {stage1_17[55]}
   );
   gpc1_1 gpc487 (
      {stage0_17[121]},
      {stage1_17[56]}
   );
   gpc1_1 gpc488 (
      {stage0_17[122]},
      {stage1_17[57]}
   );
   gpc1_1 gpc489 (
      {stage0_17[123]},
      {stage1_17[58]}
   );
   gpc1_1 gpc490 (
      {stage0_17[124]},
      {stage1_17[59]}
   );
   gpc1_1 gpc491 (
      {stage0_17[125]},
      {stage1_17[60]}
   );
   gpc1_1 gpc492 (
      {stage0_17[126]},
      {stage1_17[61]}
   );
   gpc1_1 gpc493 (
      {stage0_17[127]},
      {stage1_17[62]}
   );
   gpc1_1 gpc494 (
      {stage0_18[100]},
      {stage1_18[38]}
   );
   gpc1_1 gpc495 (
      {stage0_18[101]},
      {stage1_18[39]}
   );
   gpc1_1 gpc496 (
      {stage0_18[102]},
      {stage1_18[40]}
   );
   gpc1_1 gpc497 (
      {stage0_18[103]},
      {stage1_18[41]}
   );
   gpc1_1 gpc498 (
      {stage0_18[104]},
      {stage1_18[42]}
   );
   gpc1_1 gpc499 (
      {stage0_18[105]},
      {stage1_18[43]}
   );
   gpc1_1 gpc500 (
      {stage0_18[106]},
      {stage1_18[44]}
   );
   gpc1_1 gpc501 (
      {stage0_18[107]},
      {stage1_18[45]}
   );
   gpc1_1 gpc502 (
      {stage0_18[108]},
      {stage1_18[46]}
   );
   gpc1_1 gpc503 (
      {stage0_18[109]},
      {stage1_18[47]}
   );
   gpc1_1 gpc504 (
      {stage0_18[110]},
      {stage1_18[48]}
   );
   gpc1_1 gpc505 (
      {stage0_18[111]},
      {stage1_18[49]}
   );
   gpc1_1 gpc506 (
      {stage0_18[112]},
      {stage1_18[50]}
   );
   gpc1_1 gpc507 (
      {stage0_18[113]},
      {stage1_18[51]}
   );
   gpc1_1 gpc508 (
      {stage0_18[114]},
      {stage1_18[52]}
   );
   gpc1_1 gpc509 (
      {stage0_18[115]},
      {stage1_18[53]}
   );
   gpc1_1 gpc510 (
      {stage0_18[116]},
      {stage1_18[54]}
   );
   gpc1_1 gpc511 (
      {stage0_18[117]},
      {stage1_18[55]}
   );
   gpc1_1 gpc512 (
      {stage0_18[118]},
      {stage1_18[56]}
   );
   gpc1_1 gpc513 (
      {stage0_18[119]},
      {stage1_18[57]}
   );
   gpc1_1 gpc514 (
      {stage0_18[120]},
      {stage1_18[58]}
   );
   gpc1_1 gpc515 (
      {stage0_18[121]},
      {stage1_18[59]}
   );
   gpc1_1 gpc516 (
      {stage0_18[122]},
      {stage1_18[60]}
   );
   gpc1_1 gpc517 (
      {stage0_18[123]},
      {stage1_18[61]}
   );
   gpc1_1 gpc518 (
      {stage0_18[124]},
      {stage1_18[62]}
   );
   gpc1_1 gpc519 (
      {stage0_18[125]},
      {stage1_18[63]}
   );
   gpc1_1 gpc520 (
      {stage0_18[126]},
      {stage1_18[64]}
   );
   gpc1_1 gpc521 (
      {stage0_18[127]},
      {stage1_18[65]}
   );
   gpc1_1 gpc522 (
      {stage0_19[125]},
      {stage1_19[40]}
   );
   gpc1_1 gpc523 (
      {stage0_19[126]},
      {stage1_19[41]}
   );
   gpc1_1 gpc524 (
      {stage0_19[127]},
      {stage1_19[42]}
   );
   gpc1_1 gpc525 (
      {stage0_20[117]},
      {stage1_20[55]}
   );
   gpc1_1 gpc526 (
      {stage0_20[118]},
      {stage1_20[56]}
   );
   gpc1_1 gpc527 (
      {stage0_20[119]},
      {stage1_20[57]}
   );
   gpc1_1 gpc528 (
      {stage0_20[120]},
      {stage1_20[58]}
   );
   gpc1_1 gpc529 (
      {stage0_20[121]},
      {stage1_20[59]}
   );
   gpc1_1 gpc530 (
      {stage0_20[122]},
      {stage1_20[60]}
   );
   gpc1_1 gpc531 (
      {stage0_20[123]},
      {stage1_20[61]}
   );
   gpc1_1 gpc532 (
      {stage0_20[124]},
      {stage1_20[62]}
   );
   gpc1_1 gpc533 (
      {stage0_20[125]},
      {stage1_20[63]}
   );
   gpc1_1 gpc534 (
      {stage0_20[126]},
      {stage1_20[64]}
   );
   gpc1_1 gpc535 (
      {stage0_20[127]},
      {stage1_20[65]}
   );
   gpc1_1 gpc536 (
      {stage0_21[120]},
      {stage1_21[57]}
   );
   gpc1_1 gpc537 (
      {stage0_21[121]},
      {stage1_21[58]}
   );
   gpc1_1 gpc538 (
      {stage0_21[122]},
      {stage1_21[59]}
   );
   gpc1_1 gpc539 (
      {stage0_21[123]},
      {stage1_21[60]}
   );
   gpc1_1 gpc540 (
      {stage0_21[124]},
      {stage1_21[61]}
   );
   gpc1_1 gpc541 (
      {stage0_21[125]},
      {stage1_21[62]}
   );
   gpc1_1 gpc542 (
      {stage0_21[126]},
      {stage1_21[63]}
   );
   gpc1_1 gpc543 (
      {stage0_21[127]},
      {stage1_21[64]}
   );
   gpc1_1 gpc544 (
      {stage0_22[107]},
      {stage1_22[40]}
   );
   gpc1_1 gpc545 (
      {stage0_22[108]},
      {stage1_22[41]}
   );
   gpc1_1 gpc546 (
      {stage0_22[109]},
      {stage1_22[42]}
   );
   gpc1_1 gpc547 (
      {stage0_22[110]},
      {stage1_22[43]}
   );
   gpc1_1 gpc548 (
      {stage0_22[111]},
      {stage1_22[44]}
   );
   gpc1_1 gpc549 (
      {stage0_22[112]},
      {stage1_22[45]}
   );
   gpc1_1 gpc550 (
      {stage0_22[113]},
      {stage1_22[46]}
   );
   gpc1_1 gpc551 (
      {stage0_22[114]},
      {stage1_22[47]}
   );
   gpc1_1 gpc552 (
      {stage0_22[115]},
      {stage1_22[48]}
   );
   gpc1_1 gpc553 (
      {stage0_22[116]},
      {stage1_22[49]}
   );
   gpc1_1 gpc554 (
      {stage0_22[117]},
      {stage1_22[50]}
   );
   gpc1_1 gpc555 (
      {stage0_22[118]},
      {stage1_22[51]}
   );
   gpc1_1 gpc556 (
      {stage0_22[119]},
      {stage1_22[52]}
   );
   gpc1_1 gpc557 (
      {stage0_22[120]},
      {stage1_22[53]}
   );
   gpc1_1 gpc558 (
      {stage0_22[121]},
      {stage1_22[54]}
   );
   gpc1_1 gpc559 (
      {stage0_22[122]},
      {stage1_22[55]}
   );
   gpc1_1 gpc560 (
      {stage0_22[123]},
      {stage1_22[56]}
   );
   gpc1_1 gpc561 (
      {stage0_22[124]},
      {stage1_22[57]}
   );
   gpc1_1 gpc562 (
      {stage0_22[125]},
      {stage1_22[58]}
   );
   gpc1_1 gpc563 (
      {stage0_22[126]},
      {stage1_22[59]}
   );
   gpc1_1 gpc564 (
      {stage0_22[127]},
      {stage1_22[60]}
   );
   gpc1_1 gpc565 (
      {stage0_23[126]},
      {stage1_23[42]}
   );
   gpc1_1 gpc566 (
      {stage0_23[127]},
      {stage1_23[43]}
   );
   gpc1_1 gpc567 (
      {stage0_24[91]},
      {stage1_24[53]}
   );
   gpc1_1 gpc568 (
      {stage0_24[92]},
      {stage1_24[54]}
   );
   gpc1_1 gpc569 (
      {stage0_24[93]},
      {stage1_24[55]}
   );
   gpc1_1 gpc570 (
      {stage0_24[94]},
      {stage1_24[56]}
   );
   gpc1_1 gpc571 (
      {stage0_24[95]},
      {stage1_24[57]}
   );
   gpc1_1 gpc572 (
      {stage0_24[96]},
      {stage1_24[58]}
   );
   gpc1_1 gpc573 (
      {stage0_24[97]},
      {stage1_24[59]}
   );
   gpc1_1 gpc574 (
      {stage0_24[98]},
      {stage1_24[60]}
   );
   gpc1_1 gpc575 (
      {stage0_24[99]},
      {stage1_24[61]}
   );
   gpc1_1 gpc576 (
      {stage0_24[100]},
      {stage1_24[62]}
   );
   gpc1_1 gpc577 (
      {stage0_24[101]},
      {stage1_24[63]}
   );
   gpc1_1 gpc578 (
      {stage0_24[102]},
      {stage1_24[64]}
   );
   gpc1_1 gpc579 (
      {stage0_24[103]},
      {stage1_24[65]}
   );
   gpc1_1 gpc580 (
      {stage0_24[104]},
      {stage1_24[66]}
   );
   gpc1_1 gpc581 (
      {stage0_24[105]},
      {stage1_24[67]}
   );
   gpc1_1 gpc582 (
      {stage0_24[106]},
      {stage1_24[68]}
   );
   gpc1_1 gpc583 (
      {stage0_24[107]},
      {stage1_24[69]}
   );
   gpc1_1 gpc584 (
      {stage0_24[108]},
      {stage1_24[70]}
   );
   gpc1_1 gpc585 (
      {stage0_24[109]},
      {stage1_24[71]}
   );
   gpc1_1 gpc586 (
      {stage0_24[110]},
      {stage1_24[72]}
   );
   gpc1_1 gpc587 (
      {stage0_24[111]},
      {stage1_24[73]}
   );
   gpc1_1 gpc588 (
      {stage0_24[112]},
      {stage1_24[74]}
   );
   gpc1_1 gpc589 (
      {stage0_24[113]},
      {stage1_24[75]}
   );
   gpc1_1 gpc590 (
      {stage0_24[114]},
      {stage1_24[76]}
   );
   gpc1_1 gpc591 (
      {stage0_24[115]},
      {stage1_24[77]}
   );
   gpc1_1 gpc592 (
      {stage0_24[116]},
      {stage1_24[78]}
   );
   gpc1_1 gpc593 (
      {stage0_24[117]},
      {stage1_24[79]}
   );
   gpc1_1 gpc594 (
      {stage0_24[118]},
      {stage1_24[80]}
   );
   gpc1_1 gpc595 (
      {stage0_24[119]},
      {stage1_24[81]}
   );
   gpc1_1 gpc596 (
      {stage0_24[120]},
      {stage1_24[82]}
   );
   gpc1_1 gpc597 (
      {stage0_24[121]},
      {stage1_24[83]}
   );
   gpc1_1 gpc598 (
      {stage0_24[122]},
      {stage1_24[84]}
   );
   gpc1_1 gpc599 (
      {stage0_24[123]},
      {stage1_24[85]}
   );
   gpc1_1 gpc600 (
      {stage0_24[124]},
      {stage1_24[86]}
   );
   gpc1_1 gpc601 (
      {stage0_24[125]},
      {stage1_24[87]}
   );
   gpc1_1 gpc602 (
      {stage0_24[126]},
      {stage1_24[88]}
   );
   gpc1_1 gpc603 (
      {stage0_24[127]},
      {stage1_24[89]}
   );
   gpc1_1 gpc604 (
      {stage0_25[108]},
      {stage1_25[50]}
   );
   gpc1_1 gpc605 (
      {stage0_25[109]},
      {stage1_25[51]}
   );
   gpc1_1 gpc606 (
      {stage0_25[110]},
      {stage1_25[52]}
   );
   gpc1_1 gpc607 (
      {stage0_25[111]},
      {stage1_25[53]}
   );
   gpc1_1 gpc608 (
      {stage0_25[112]},
      {stage1_25[54]}
   );
   gpc1_1 gpc609 (
      {stage0_25[113]},
      {stage1_25[55]}
   );
   gpc1_1 gpc610 (
      {stage0_25[114]},
      {stage1_25[56]}
   );
   gpc1_1 gpc611 (
      {stage0_25[115]},
      {stage1_25[57]}
   );
   gpc1_1 gpc612 (
      {stage0_25[116]},
      {stage1_25[58]}
   );
   gpc1_1 gpc613 (
      {stage0_25[117]},
      {stage1_25[59]}
   );
   gpc1_1 gpc614 (
      {stage0_25[118]},
      {stage1_25[60]}
   );
   gpc1_1 gpc615 (
      {stage0_25[119]},
      {stage1_25[61]}
   );
   gpc1_1 gpc616 (
      {stage0_25[120]},
      {stage1_25[62]}
   );
   gpc1_1 gpc617 (
      {stage0_25[121]},
      {stage1_25[63]}
   );
   gpc1_1 gpc618 (
      {stage0_25[122]},
      {stage1_25[64]}
   );
   gpc1_1 gpc619 (
      {stage0_25[123]},
      {stage1_25[65]}
   );
   gpc1_1 gpc620 (
      {stage0_25[124]},
      {stage1_25[66]}
   );
   gpc1_1 gpc621 (
      {stage0_25[125]},
      {stage1_25[67]}
   );
   gpc1_1 gpc622 (
      {stage0_25[126]},
      {stage1_25[68]}
   );
   gpc1_1 gpc623 (
      {stage0_25[127]},
      {stage1_25[69]}
   );
   gpc1_1 gpc624 (
      {stage0_26[94]},
      {stage1_26[35]}
   );
   gpc1_1 gpc625 (
      {stage0_26[95]},
      {stage1_26[36]}
   );
   gpc1_1 gpc626 (
      {stage0_26[96]},
      {stage1_26[37]}
   );
   gpc1_1 gpc627 (
      {stage0_26[97]},
      {stage1_26[38]}
   );
   gpc1_1 gpc628 (
      {stage0_26[98]},
      {stage1_26[39]}
   );
   gpc1_1 gpc629 (
      {stage0_26[99]},
      {stage1_26[40]}
   );
   gpc1_1 gpc630 (
      {stage0_26[100]},
      {stage1_26[41]}
   );
   gpc1_1 gpc631 (
      {stage0_26[101]},
      {stage1_26[42]}
   );
   gpc1_1 gpc632 (
      {stage0_26[102]},
      {stage1_26[43]}
   );
   gpc1_1 gpc633 (
      {stage0_26[103]},
      {stage1_26[44]}
   );
   gpc1_1 gpc634 (
      {stage0_26[104]},
      {stage1_26[45]}
   );
   gpc1_1 gpc635 (
      {stage0_26[105]},
      {stage1_26[46]}
   );
   gpc1_1 gpc636 (
      {stage0_26[106]},
      {stage1_26[47]}
   );
   gpc1_1 gpc637 (
      {stage0_26[107]},
      {stage1_26[48]}
   );
   gpc1_1 gpc638 (
      {stage0_26[108]},
      {stage1_26[49]}
   );
   gpc1_1 gpc639 (
      {stage0_26[109]},
      {stage1_26[50]}
   );
   gpc1_1 gpc640 (
      {stage0_26[110]},
      {stage1_26[51]}
   );
   gpc1_1 gpc641 (
      {stage0_26[111]},
      {stage1_26[52]}
   );
   gpc1_1 gpc642 (
      {stage0_26[112]},
      {stage1_26[53]}
   );
   gpc1_1 gpc643 (
      {stage0_26[113]},
      {stage1_26[54]}
   );
   gpc1_1 gpc644 (
      {stage0_26[114]},
      {stage1_26[55]}
   );
   gpc1_1 gpc645 (
      {stage0_26[115]},
      {stage1_26[56]}
   );
   gpc1_1 gpc646 (
      {stage0_26[116]},
      {stage1_26[57]}
   );
   gpc1_1 gpc647 (
      {stage0_26[117]},
      {stage1_26[58]}
   );
   gpc1_1 gpc648 (
      {stage0_26[118]},
      {stage1_26[59]}
   );
   gpc1_1 gpc649 (
      {stage0_26[119]},
      {stage1_26[60]}
   );
   gpc1_1 gpc650 (
      {stage0_26[120]},
      {stage1_26[61]}
   );
   gpc1_1 gpc651 (
      {stage0_26[121]},
      {stage1_26[62]}
   );
   gpc1_1 gpc652 (
      {stage0_26[122]},
      {stage1_26[63]}
   );
   gpc1_1 gpc653 (
      {stage0_26[123]},
      {stage1_26[64]}
   );
   gpc1_1 gpc654 (
      {stage0_26[124]},
      {stage1_26[65]}
   );
   gpc1_1 gpc655 (
      {stage0_26[125]},
      {stage1_26[66]}
   );
   gpc1_1 gpc656 (
      {stage0_26[126]},
      {stage1_26[67]}
   );
   gpc1_1 gpc657 (
      {stage0_26[127]},
      {stage1_26[68]}
   );
   gpc1_1 gpc658 (
      {stage0_27[111]},
      {stage1_27[39]}
   );
   gpc1_1 gpc659 (
      {stage0_27[112]},
      {stage1_27[40]}
   );
   gpc1_1 gpc660 (
      {stage0_27[113]},
      {stage1_27[41]}
   );
   gpc1_1 gpc661 (
      {stage0_27[114]},
      {stage1_27[42]}
   );
   gpc1_1 gpc662 (
      {stage0_27[115]},
      {stage1_27[43]}
   );
   gpc1_1 gpc663 (
      {stage0_27[116]},
      {stage1_27[44]}
   );
   gpc1_1 gpc664 (
      {stage0_27[117]},
      {stage1_27[45]}
   );
   gpc1_1 gpc665 (
      {stage0_27[118]},
      {stage1_27[46]}
   );
   gpc1_1 gpc666 (
      {stage0_27[119]},
      {stage1_27[47]}
   );
   gpc1_1 gpc667 (
      {stage0_27[120]},
      {stage1_27[48]}
   );
   gpc1_1 gpc668 (
      {stage0_27[121]},
      {stage1_27[49]}
   );
   gpc1_1 gpc669 (
      {stage0_27[122]},
      {stage1_27[50]}
   );
   gpc1_1 gpc670 (
      {stage0_27[123]},
      {stage1_27[51]}
   );
   gpc1_1 gpc671 (
      {stage0_27[124]},
      {stage1_27[52]}
   );
   gpc1_1 gpc672 (
      {stage0_27[125]},
      {stage1_27[53]}
   );
   gpc1_1 gpc673 (
      {stage0_27[126]},
      {stage1_27[54]}
   );
   gpc1_1 gpc674 (
      {stage0_27[127]},
      {stage1_27[55]}
   );
   gpc1_1 gpc675 (
      {stage0_28[125]},
      {stage1_28[53]}
   );
   gpc1_1 gpc676 (
      {stage0_28[126]},
      {stage1_28[54]}
   );
   gpc1_1 gpc677 (
      {stage0_28[127]},
      {stage1_28[55]}
   );
   gpc1_1 gpc678 (
      {stage0_29[126]},
      {stage1_29[55]}
   );
   gpc1_1 gpc679 (
      {stage0_29[127]},
      {stage1_29[56]}
   );
   gpc1_1 gpc680 (
      {stage0_30[108]},
      {stage1_30[41]}
   );
   gpc1_1 gpc681 (
      {stage0_30[109]},
      {stage1_30[42]}
   );
   gpc1_1 gpc682 (
      {stage0_30[110]},
      {stage1_30[43]}
   );
   gpc1_1 gpc683 (
      {stage0_30[111]},
      {stage1_30[44]}
   );
   gpc1_1 gpc684 (
      {stage0_30[112]},
      {stage1_30[45]}
   );
   gpc1_1 gpc685 (
      {stage0_30[113]},
      {stage1_30[46]}
   );
   gpc1_1 gpc686 (
      {stage0_30[114]},
      {stage1_30[47]}
   );
   gpc1_1 gpc687 (
      {stage0_30[115]},
      {stage1_30[48]}
   );
   gpc1_1 gpc688 (
      {stage0_30[116]},
      {stage1_30[49]}
   );
   gpc1_1 gpc689 (
      {stage0_30[117]},
      {stage1_30[50]}
   );
   gpc1_1 gpc690 (
      {stage0_30[118]},
      {stage1_30[51]}
   );
   gpc1_1 gpc691 (
      {stage0_30[119]},
      {stage1_30[52]}
   );
   gpc1_1 gpc692 (
      {stage0_30[120]},
      {stage1_30[53]}
   );
   gpc1_1 gpc693 (
      {stage0_30[121]},
      {stage1_30[54]}
   );
   gpc1_1 gpc694 (
      {stage0_30[122]},
      {stage1_30[55]}
   );
   gpc1_1 gpc695 (
      {stage0_30[123]},
      {stage1_30[56]}
   );
   gpc1_1 gpc696 (
      {stage0_30[124]},
      {stage1_30[57]}
   );
   gpc1_1 gpc697 (
      {stage0_30[125]},
      {stage1_30[58]}
   );
   gpc1_1 gpc698 (
      {stage0_30[126]},
      {stage1_30[59]}
   );
   gpc1_1 gpc699 (
      {stage0_30[127]},
      {stage1_30[60]}
   );
   gpc1_1 gpc700 (
      {stage0_31[96]},
      {stage1_31[39]}
   );
   gpc1_1 gpc701 (
      {stage0_31[97]},
      {stage1_31[40]}
   );
   gpc1_1 gpc702 (
      {stage0_31[98]},
      {stage1_31[41]}
   );
   gpc1_1 gpc703 (
      {stage0_31[99]},
      {stage1_31[42]}
   );
   gpc1_1 gpc704 (
      {stage0_31[100]},
      {stage1_31[43]}
   );
   gpc1_1 gpc705 (
      {stage0_31[101]},
      {stage1_31[44]}
   );
   gpc1_1 gpc706 (
      {stage0_31[102]},
      {stage1_31[45]}
   );
   gpc1_1 gpc707 (
      {stage0_31[103]},
      {stage1_31[46]}
   );
   gpc1_1 gpc708 (
      {stage0_31[104]},
      {stage1_31[47]}
   );
   gpc1_1 gpc709 (
      {stage0_31[105]},
      {stage1_31[48]}
   );
   gpc1_1 gpc710 (
      {stage0_31[106]},
      {stage1_31[49]}
   );
   gpc1_1 gpc711 (
      {stage0_31[107]},
      {stage1_31[50]}
   );
   gpc1_1 gpc712 (
      {stage0_31[108]},
      {stage1_31[51]}
   );
   gpc1_1 gpc713 (
      {stage0_31[109]},
      {stage1_31[52]}
   );
   gpc1_1 gpc714 (
      {stage0_31[110]},
      {stage1_31[53]}
   );
   gpc1_1 gpc715 (
      {stage0_31[111]},
      {stage1_31[54]}
   );
   gpc1_1 gpc716 (
      {stage0_31[112]},
      {stage1_31[55]}
   );
   gpc1_1 gpc717 (
      {stage0_31[113]},
      {stage1_31[56]}
   );
   gpc1_1 gpc718 (
      {stage0_31[114]},
      {stage1_31[57]}
   );
   gpc1_1 gpc719 (
      {stage0_31[115]},
      {stage1_31[58]}
   );
   gpc1_1 gpc720 (
      {stage0_31[116]},
      {stage1_31[59]}
   );
   gpc1_1 gpc721 (
      {stage0_31[117]},
      {stage1_31[60]}
   );
   gpc1_1 gpc722 (
      {stage0_31[118]},
      {stage1_31[61]}
   );
   gpc1_1 gpc723 (
      {stage0_31[119]},
      {stage1_31[62]}
   );
   gpc1_1 gpc724 (
      {stage0_31[120]},
      {stage1_31[63]}
   );
   gpc1_1 gpc725 (
      {stage0_31[121]},
      {stage1_31[64]}
   );
   gpc1_1 gpc726 (
      {stage0_31[122]},
      {stage1_31[65]}
   );
   gpc1_1 gpc727 (
      {stage0_31[123]},
      {stage1_31[66]}
   );
   gpc1_1 gpc728 (
      {stage0_31[124]},
      {stage1_31[67]}
   );
   gpc1_1 gpc729 (
      {stage0_31[125]},
      {stage1_31[68]}
   );
   gpc1_1 gpc730 (
      {stage0_31[126]},
      {stage1_31[69]}
   );
   gpc1_1 gpc731 (
      {stage0_31[127]},
      {stage1_31[70]}
   );
   gpc606_5 gpc732 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0]}
   );
   gpc606_5 gpc733 (
      {stage1_1[6], stage1_1[7], stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11]},
      {stage1_3[6], stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11]},
      {stage2_5[1],stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1]}
   );
   gpc606_5 gpc734 (
      {stage1_1[12], stage1_1[13], stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17]},
      {stage1_3[12], stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17]},
      {stage2_5[2],stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2]}
   );
   gpc606_5 gpc735 (
      {stage1_1[18], stage1_1[19], stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23]},
      {stage1_3[18], stage1_3[19], stage1_3[20], stage1_3[21], stage1_3[22], stage1_3[23]},
      {stage2_5[3],stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3]}
   );
   gpc606_5 gpc736 (
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[4],stage2_4[4],stage2_3[4],stage2_2[4]}
   );
   gpc606_5 gpc737 (
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[5],stage2_4[5],stage2_3[5],stage2_2[5]}
   );
   gpc606_5 gpc738 (
      {stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[6],stage2_4[6],stage2_3[6],stage2_2[6]}
   );
   gpc615_5 gpc739 (
      {stage1_2[18], stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22]},
      {stage1_3[24]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[7],stage2_4[7],stage2_3[7],stage2_2[7]}
   );
   gpc615_5 gpc740 (
      {stage1_2[23], stage1_2[24], stage1_2[25], stage1_2[26], stage1_2[27]},
      {stage1_3[25]},
      {stage1_4[24], stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29]},
      {stage2_6[4],stage2_5[8],stage2_4[8],stage2_3[8],stage2_2[8]}
   );
   gpc615_5 gpc741 (
      {stage1_2[28], stage1_2[29], stage1_2[30], stage1_2[31], stage1_2[32]},
      {stage1_3[26]},
      {stage1_4[30], stage1_4[31], stage1_4[32], stage1_4[33], stage1_4[34], stage1_4[35]},
      {stage2_6[5],stage2_5[9],stage2_4[9],stage2_3[9],stage2_2[9]}
   );
   gpc615_5 gpc742 (
      {stage1_2[33], stage1_2[34], stage1_2[35], stage1_2[36], stage1_2[37]},
      {stage1_3[27]},
      {stage1_4[36], stage1_4[37], stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41]},
      {stage2_6[6],stage2_5[10],stage2_4[10],stage2_3[10],stage2_2[10]}
   );
   gpc615_5 gpc743 (
      {stage1_2[38], stage1_2[39], stage1_2[40], stage1_2[41], stage1_2[42]},
      {stage1_3[28]},
      {stage1_4[42], stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage2_6[7],stage2_5[11],stage2_4[11],stage2_3[11],stage2_2[11]}
   );
   gpc615_5 gpc744 (
      {stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33]},
      {stage1_4[48]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[8],stage2_5[12],stage2_4[12],stage2_3[12]}
   );
   gpc615_5 gpc745 (
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38]},
      {stage1_4[49]},
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage2_7[1],stage2_6[9],stage2_5[13],stage2_4[13],stage2_3[13]}
   );
   gpc606_5 gpc746 (
      {stage1_4[50], stage1_4[51], stage1_4[52], stage1_4[53], stage1_4[54], stage1_4[55]},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[2],stage2_6[10],stage2_5[14],stage2_4[14]}
   );
   gpc606_5 gpc747 (
      {stage1_5[12], stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[1],stage2_7[3],stage2_6[11],stage2_5[15]}
   );
   gpc606_5 gpc748 (
      {stage1_5[18], stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23]},
      {stage1_7[6], stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11]},
      {stage2_9[1],stage2_8[2],stage2_7[4],stage2_6[12],stage2_5[16]}
   );
   gpc606_5 gpc749 (
      {stage1_5[24], stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29]},
      {stage1_7[12], stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17]},
      {stage2_9[2],stage2_8[3],stage2_7[5],stage2_6[13],stage2_5[17]}
   );
   gpc606_5 gpc750 (
      {stage1_5[30], stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35]},
      {stage1_7[18], stage1_7[19], stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23]},
      {stage2_9[3],stage2_8[4],stage2_7[6],stage2_6[14],stage2_5[18]}
   );
   gpc606_5 gpc751 (
      {stage1_5[36], stage1_5[37], stage1_5[38], stage1_5[39], stage1_5[40], stage1_5[41]},
      {stage1_7[24], stage1_7[25], stage1_7[26], stage1_7[27], stage1_7[28], stage1_7[29]},
      {stage2_9[4],stage2_8[5],stage2_7[7],stage2_6[15],stage2_5[19]}
   );
   gpc606_5 gpc752 (
      {stage1_5[42], stage1_5[43], stage1_5[44], stage1_5[45], stage1_5[46], stage1_5[47]},
      {stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33], stage1_7[34], stage1_7[35]},
      {stage2_9[5],stage2_8[6],stage2_7[8],stage2_6[16],stage2_5[20]}
   );
   gpc606_5 gpc753 (
      {stage1_5[48], stage1_5[49], stage1_5[50], stage1_5[51], stage1_5[52], stage1_5[53]},
      {stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40], stage1_7[41]},
      {stage2_9[6],stage2_8[7],stage2_7[9],stage2_6[17],stage2_5[21]}
   );
   gpc606_5 gpc754 (
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[7],stage2_8[8],stage2_7[10],stage2_6[18]}
   );
   gpc606_5 gpc755 (
      {stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[8],stage2_8[9],stage2_7[11],stage2_6[19]}
   );
   gpc615_5 gpc756 (
      {stage1_6[18], stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22]},
      {stage1_7[42]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[9],stage2_8[10],stage2_7[12],stage2_6[20]}
   );
   gpc615_5 gpc757 (
      {stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46], stage1_7[47]},
      {stage1_8[18]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage2_11[0],stage2_10[3],stage2_9[10],stage2_8[11],stage2_7[13]}
   );
   gpc615_5 gpc758 (
      {stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52]},
      {stage1_8[19]},
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage2_11[1],stage2_10[4],stage2_9[11],stage2_8[12],stage2_7[14]}
   );
   gpc615_5 gpc759 (
      {stage1_7[53], stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57]},
      {stage1_8[20]},
      {stage1_9[12], stage1_9[13], stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17]},
      {stage2_11[2],stage2_10[5],stage2_9[12],stage2_8[13],stage2_7[15]}
   );
   gpc615_5 gpc760 (
      {stage1_7[58], stage1_7[59], stage1_7[60], stage1_7[61], stage1_7[62]},
      {stage1_8[21]},
      {stage1_9[18], stage1_9[19], stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23]},
      {stage2_11[3],stage2_10[6],stage2_9[13],stage2_8[14],stage2_7[16]}
   );
   gpc615_5 gpc761 (
      {stage1_7[63], stage1_7[64], stage1_7[65], stage1_7[66], stage1_7[67]},
      {stage1_8[22]},
      {stage1_9[24], stage1_9[25], stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29]},
      {stage2_11[4],stage2_10[7],stage2_9[14],stage2_8[15],stage2_7[17]}
   );
   gpc606_5 gpc762 (
      {stage1_8[23], stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28]},
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage2_12[0],stage2_11[5],stage2_10[8],stage2_9[15],stage2_8[16]}
   );
   gpc606_5 gpc763 (
      {stage1_8[29], stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34]},
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage2_12[1],stage2_11[6],stage2_10[9],stage2_9[16],stage2_8[17]}
   );
   gpc606_5 gpc764 (
      {stage1_9[30], stage1_9[31], stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[2],stage2_11[7],stage2_10[10],stage2_9[17]}
   );
   gpc606_5 gpc765 (
      {stage1_9[36], stage1_9[37], stage1_9[38], stage1_9[39], stage1_9[40], stage1_9[41]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[3],stage2_11[8],stage2_10[11],stage2_9[18]}
   );
   gpc606_5 gpc766 (
      {stage1_9[42], stage1_9[43], stage1_9[44], stage1_9[45], stage1_9[46], stage1_9[47]},
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17]},
      {stage2_13[2],stage2_12[4],stage2_11[9],stage2_10[12],stage2_9[19]}
   );
   gpc606_5 gpc767 (
      {stage1_9[48], stage1_9[49], stage1_9[50], stage1_9[51], stage1_9[52], stage1_9[53]},
      {stage1_11[18], stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23]},
      {stage2_13[3],stage2_12[5],stage2_11[10],stage2_10[13],stage2_9[20]}
   );
   gpc606_5 gpc768 (
      {stage1_9[54], stage1_9[55], stage1_9[56], stage1_9[57], stage1_9[58], stage1_9[59]},
      {stage1_11[24], stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29]},
      {stage2_13[4],stage2_12[6],stage2_11[11],stage2_10[14],stage2_9[21]}
   );
   gpc606_5 gpc769 (
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[5],stage2_12[7],stage2_11[12],stage2_10[15]}
   );
   gpc606_5 gpc770 (
      {stage1_10[18], stage1_10[19], stage1_10[20], stage1_10[21], stage1_10[22], stage1_10[23]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[6],stage2_12[8],stage2_11[13],stage2_10[16]}
   );
   gpc606_5 gpc771 (
      {stage1_10[24], stage1_10[25], stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[7],stage2_12[9],stage2_11[14],stage2_10[17]}
   );
   gpc606_5 gpc772 (
      {stage1_10[30], stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[8],stage2_12[10],stage2_11[15],stage2_10[18]}
   );
   gpc606_5 gpc773 (
      {stage1_10[36], stage1_10[37], stage1_10[38], stage1_10[39], stage1_10[40], stage1_10[41]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[9],stage2_12[11],stage2_11[16],stage2_10[19]}
   );
   gpc606_5 gpc774 (
      {stage1_10[42], stage1_10[43], stage1_10[44], stage1_10[45], stage1_10[46], stage1_10[47]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[10],stage2_12[12],stage2_11[17],stage2_10[20]}
   );
   gpc606_5 gpc775 (
      {stage1_10[48], stage1_10[49], stage1_10[50], stage1_10[51], stage1_10[52], stage1_10[53]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[11],stage2_12[13],stage2_11[18],stage2_10[21]}
   );
   gpc615_5 gpc776 (
      {stage1_11[30], stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34]},
      {stage1_12[42]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[7],stage2_13[12],stage2_12[14],stage2_11[19]}
   );
   gpc615_5 gpc777 (
      {stage1_11[35], stage1_11[36], stage1_11[37], stage1_11[38], stage1_11[39]},
      {stage1_12[43]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[8],stage2_13[13],stage2_12[15],stage2_11[20]}
   );
   gpc615_5 gpc778 (
      {stage1_11[40], stage1_11[41], stage1_11[42], stage1_11[43], stage1_11[44]},
      {stage1_12[44]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[9],stage2_13[14],stage2_12[16],stage2_11[21]}
   );
   gpc615_5 gpc779 (
      {stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48], stage1_11[49]},
      {stage1_12[45]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[10],stage2_13[15],stage2_12[17],stage2_11[22]}
   );
   gpc615_5 gpc780 (
      {stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53], stage1_11[54]},
      {stage1_12[46]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[11],stage2_13[16],stage2_12[18],stage2_11[23]}
   );
   gpc606_5 gpc781 (
      {stage1_12[47], stage1_12[48], stage1_12[49], stage1_12[50], stage1_12[51], stage1_12[52]},
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage2_16[0],stage2_15[5],stage2_14[12],stage2_13[17],stage2_12[19]}
   );
   gpc606_5 gpc782 (
      {stage1_12[53], stage1_12[54], stage1_12[55], stage1_12[56], stage1_12[57], 1'b0},
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage2_16[1],stage2_15[6],stage2_14[13],stage2_13[18],stage2_12[20]}
   );
   gpc606_5 gpc783 (
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[2],stage2_15[7],stage2_14[14],stage2_13[19]}
   );
   gpc606_5 gpc784 (
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage2_17[1],stage2_16[3],stage2_15[8],stage2_14[15],stage2_13[20]}
   );
   gpc606_5 gpc785 (
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage2_17[2],stage2_16[4],stage2_15[9],stage2_14[16],stage2_13[21]}
   );
   gpc615_5 gpc786 (
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16]},
      {stage1_15[18]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[3],stage2_16[5],stage2_15[10],stage2_14[17]}
   );
   gpc615_5 gpc787 (
      {stage1_14[17], stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21]},
      {stage1_15[19]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[4],stage2_16[6],stage2_15[11],stage2_14[18]}
   );
   gpc615_5 gpc788 (
      {stage1_14[22], stage1_14[23], stage1_14[24], stage1_14[25], stage1_14[26]},
      {stage1_15[20]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[5],stage2_16[7],stage2_15[12],stage2_14[19]}
   );
   gpc615_5 gpc789 (
      {stage1_14[27], stage1_14[28], stage1_14[29], stage1_14[30], stage1_14[31]},
      {stage1_15[21]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[6],stage2_16[8],stage2_15[13],stage2_14[20]}
   );
   gpc615_5 gpc790 (
      {stage1_14[32], stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36]},
      {stage1_15[22]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[7],stage2_16[9],stage2_15[14],stage2_14[21]}
   );
   gpc615_5 gpc791 (
      {stage1_14[37], stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41]},
      {stage1_15[23]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[8],stage2_16[10],stage2_15[15],stage2_14[22]}
   );
   gpc615_5 gpc792 (
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28]},
      {stage1_16[36]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5]},
      {stage2_19[0],stage2_18[6],stage2_17[9],stage2_16[11],stage2_15[16]}
   );
   gpc615_5 gpc793 (
      {stage1_15[29], stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33]},
      {stage1_16[37]},
      {stage1_17[6], stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11]},
      {stage2_19[1],stage2_18[7],stage2_17[10],stage2_16[12],stage2_15[17]}
   );
   gpc615_5 gpc794 (
      {stage1_15[34], stage1_15[35], stage1_15[36], stage1_15[37], stage1_15[38]},
      {stage1_16[38]},
      {stage1_17[12], stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17]},
      {stage2_19[2],stage2_18[8],stage2_17[11],stage2_16[13],stage2_15[18]}
   );
   gpc615_5 gpc795 (
      {stage1_15[39], stage1_15[40], stage1_15[41], stage1_15[42], stage1_15[43]},
      {stage1_16[39]},
      {stage1_17[18], stage1_17[19], stage1_17[20], stage1_17[21], stage1_17[22], stage1_17[23]},
      {stage2_19[3],stage2_18[9],stage2_17[12],stage2_16[14],stage2_15[19]}
   );
   gpc606_5 gpc796 (
      {stage1_16[40], stage1_16[41], stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[4],stage2_18[10],stage2_17[13],stage2_16[15]}
   );
   gpc606_5 gpc797 (
      {stage1_16[46], stage1_16[47], stage1_16[48], stage1_16[49], stage1_16[50], stage1_16[51]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], stage1_18[11]},
      {stage2_20[1],stage2_19[5],stage2_18[11],stage2_17[14],stage2_16[16]}
   );
   gpc606_5 gpc798 (
      {stage1_16[52], stage1_16[53], stage1_16[54], stage1_16[55], stage1_16[56], stage1_16[57]},
      {stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16], stage1_18[17]},
      {stage2_20[2],stage2_19[6],stage2_18[12],stage2_17[15],stage2_16[17]}
   );
   gpc606_5 gpc799 (
      {stage1_16[58], stage1_16[59], stage1_16[60], stage1_16[61], stage1_16[62], stage1_16[63]},
      {stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22], stage1_18[23]},
      {stage2_20[3],stage2_19[7],stage2_18[13],stage2_17[16],stage2_16[18]}
   );
   gpc606_5 gpc800 (
      {stage1_16[64], stage1_16[65], stage1_16[66], stage1_16[67], stage1_16[68], stage1_16[69]},
      {stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28], stage1_18[29]},
      {stage2_20[4],stage2_19[8],stage2_18[14],stage2_17[17],stage2_16[19]}
   );
   gpc606_5 gpc801 (
      {stage1_16[70], stage1_16[71], stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75]},
      {stage1_18[30], stage1_18[31], stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35]},
      {stage2_20[5],stage2_19[9],stage2_18[15],stage2_17[18],stage2_16[20]}
   );
   gpc606_5 gpc802 (
      {stage1_16[76], stage1_16[77], stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81]},
      {stage1_18[36], stage1_18[37], stage1_18[38], stage1_18[39], stage1_18[40], stage1_18[41]},
      {stage2_20[6],stage2_19[10],stage2_18[16],stage2_17[19],stage2_16[21]}
   );
   gpc615_5 gpc803 (
      {stage1_16[82], stage1_16[83], stage1_16[84], stage1_16[85], stage1_16[86]},
      {stage1_17[24]},
      {stage1_18[42], stage1_18[43], stage1_18[44], stage1_18[45], stage1_18[46], stage1_18[47]},
      {stage2_20[7],stage2_19[11],stage2_18[17],stage2_17[20],stage2_16[22]}
   );
   gpc606_5 gpc804 (
      {stage1_17[25], stage1_17[26], stage1_17[27], stage1_17[28], stage1_17[29], stage1_17[30]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[8],stage2_19[12],stage2_18[18],stage2_17[21]}
   );
   gpc606_5 gpc805 (
      {stage1_17[31], stage1_17[32], stage1_17[33], stage1_17[34], stage1_17[35], stage1_17[36]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[9],stage2_19[13],stage2_18[19],stage2_17[22]}
   );
   gpc615_5 gpc806 (
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16]},
      {stage1_20[0]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[0],stage2_21[2],stage2_20[10],stage2_19[14]}
   );
   gpc615_5 gpc807 (
      {stage1_19[17], stage1_19[18], stage1_19[19], stage1_19[20], stage1_19[21]},
      {stage1_20[1]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[1],stage2_21[3],stage2_20[11],stage2_19[15]}
   );
   gpc615_5 gpc808 (
      {stage1_19[22], stage1_19[23], stage1_19[24], stage1_19[25], stage1_19[26]},
      {stage1_20[2]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[2],stage2_21[4],stage2_20[12],stage2_19[16]}
   );
   gpc615_5 gpc809 (
      {stage1_19[27], stage1_19[28], stage1_19[29], stage1_19[30], stage1_19[31]},
      {stage1_20[3]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[3],stage2_21[5],stage2_20[13],stage2_19[17]}
   );
   gpc615_5 gpc810 (
      {stage1_19[32], stage1_19[33], stage1_19[34], stage1_19[35], stage1_19[36]},
      {stage1_20[4]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[4],stage2_21[6],stage2_20[14],stage2_19[18]}
   );
   gpc615_5 gpc811 (
      {stage1_19[37], stage1_19[38], stage1_19[39], stage1_19[40], stage1_19[41]},
      {stage1_20[5]},
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage2_23[5],stage2_22[5],stage2_21[7],stage2_20[15],stage2_19[19]}
   );
   gpc606_5 gpc812 (
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[6],stage2_22[6],stage2_21[8],stage2_20[16]}
   );
   gpc606_5 gpc813 (
      {stage1_20[12], stage1_20[13], stage1_20[14], stage1_20[15], stage1_20[16], stage1_20[17]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[7],stage2_22[7],stage2_21[9],stage2_20[17]}
   );
   gpc606_5 gpc814 (
      {stage1_20[18], stage1_20[19], stage1_20[20], stage1_20[21], stage1_20[22], stage1_20[23]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[8],stage2_22[8],stage2_21[10],stage2_20[18]}
   );
   gpc606_5 gpc815 (
      {stage1_20[24], stage1_20[25], stage1_20[26], stage1_20[27], stage1_20[28], stage1_20[29]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[9],stage2_22[9],stage2_21[11],stage2_20[19]}
   );
   gpc606_5 gpc816 (
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[4],stage2_23[10],stage2_22[10],stage2_21[12]}
   );
   gpc606_5 gpc817 (
      {stage1_21[42], stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[5],stage2_23[11],stage2_22[11],stage2_21[13]}
   );
   gpc606_5 gpc818 (
      {stage1_21[48], stage1_21[49], stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53]},
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage2_25[2],stage2_24[6],stage2_23[12],stage2_22[12],stage2_21[14]}
   );
   gpc606_5 gpc819 (
      {stage1_21[54], stage1_21[55], stage1_21[56], stage1_21[57], stage1_21[58], stage1_21[59]},
      {stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21], stage1_23[22], stage1_23[23]},
      {stage2_25[3],stage2_24[7],stage2_23[13],stage2_22[13],stage2_21[15]}
   );
   gpc606_5 gpc820 (
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage1_24[0], stage1_24[1], stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5]},
      {stage2_26[0],stage2_25[4],stage2_24[8],stage2_23[14],stage2_22[14]}
   );
   gpc606_5 gpc821 (
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage1_24[6], stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage2_26[1],stage2_25[5],stage2_24[9],stage2_23[15],stage2_22[15]}
   );
   gpc606_5 gpc822 (
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage1_24[12], stage1_24[13], stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17]},
      {stage2_26[2],stage2_25[6],stage2_24[10],stage2_23[16],stage2_22[16]}
   );
   gpc606_5 gpc823 (
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage1_24[18], stage1_24[19], stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23]},
      {stage2_26[3],stage2_25[7],stage2_24[11],stage2_23[17],stage2_22[17]}
   );
   gpc615_5 gpc824 (
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52]},
      {stage1_23[24]},
      {stage1_24[24], stage1_24[25], stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29]},
      {stage2_26[4],stage2_25[8],stage2_24[12],stage2_23[18],stage2_22[18]}
   );
   gpc615_5 gpc825 (
      {stage1_23[25], stage1_23[26], stage1_23[27], stage1_23[28], stage1_23[29]},
      {stage1_24[30]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[5],stage2_25[9],stage2_24[13],stage2_23[19]}
   );
   gpc606_5 gpc826 (
      {stage1_24[31], stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35], stage1_24[36]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[1],stage2_26[6],stage2_25[10],stage2_24[14]}
   );
   gpc606_5 gpc827 (
      {stage1_24[37], stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41], stage1_24[42]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[2],stage2_26[7],stage2_25[11],stage2_24[15]}
   );
   gpc606_5 gpc828 (
      {stage1_24[43], stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47], stage1_24[48]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[3],stage2_26[8],stage2_25[12],stage2_24[16]}
   );
   gpc606_5 gpc829 (
      {stage1_24[49], stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53], stage1_24[54]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[4],stage2_26[9],stage2_25[13],stage2_24[17]}
   );
   gpc606_5 gpc830 (
      {stage1_24[55], stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59], stage1_24[60]},
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage2_28[4],stage2_27[5],stage2_26[10],stage2_25[14],stage2_24[18]}
   );
   gpc606_5 gpc831 (
      {stage1_24[61], stage1_24[62], stage1_24[63], stage1_24[64], stage1_24[65], stage1_24[66]},
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage2_28[5],stage2_27[6],stage2_26[11],stage2_25[15],stage2_24[19]}
   );
   gpc606_5 gpc832 (
      {stage1_24[67], stage1_24[68], stage1_24[69], stage1_24[70], stage1_24[71], stage1_24[72]},
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage2_28[6],stage2_27[7],stage2_26[12],stage2_25[16],stage2_24[20]}
   );
   gpc606_5 gpc833 (
      {stage1_24[73], stage1_24[74], stage1_24[75], stage1_24[76], stage1_24[77], stage1_24[78]},
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage2_28[7],stage2_27[8],stage2_26[13],stage2_25[17],stage2_24[21]}
   );
   gpc606_5 gpc834 (
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[8],stage2_27[9],stage2_26[14],stage2_25[18]}
   );
   gpc606_5 gpc835 (
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], stage1_27[11]},
      {stage2_29[1],stage2_28[9],stage2_27[10],stage2_26[15],stage2_25[19]}
   );
   gpc606_5 gpc836 (
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage1_27[12], stage1_27[13], stage1_27[14], stage1_27[15], stage1_27[16], stage1_27[17]},
      {stage2_29[2],stage2_28[10],stage2_27[11],stage2_26[16],stage2_25[20]}
   );
   gpc606_5 gpc837 (
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage1_27[18], stage1_27[19], stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23]},
      {stage2_29[3],stage2_28[11],stage2_27[12],stage2_26[17],stage2_25[21]}
   );
   gpc606_5 gpc838 (
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage1_27[24], stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28], stage1_27[29]},
      {stage2_29[4],stage2_28[12],stage2_27[13],stage2_26[18],stage2_25[22]}
   );
   gpc606_5 gpc839 (
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33], stage1_27[34], stage1_27[35]},
      {stage2_29[5],stage2_28[13],stage2_27[14],stage2_26[19],stage2_25[23]}
   );
   gpc606_5 gpc840 (
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage1_27[36], stage1_27[37], stage1_27[38], stage1_27[39], stage1_27[40], stage1_27[41]},
      {stage2_29[6],stage2_28[14],stage2_27[15],stage2_26[20],stage2_25[24]}
   );
   gpc606_5 gpc841 (
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[7],stage2_28[15],stage2_27[16],stage2_26[21]}
   );
   gpc606_5 gpc842 (
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[0],stage2_30[1],stage2_29[8],stage2_28[16]}
   );
   gpc606_5 gpc843 (
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage2_32[1],stage2_31[1],stage2_30[2],stage2_29[9],stage2_28[17]}
   );
   gpc606_5 gpc844 (
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16], stage1_30[17]},
      {stage2_32[2],stage2_31[2],stage2_30[3],stage2_29[10],stage2_28[18]}
   );
   gpc606_5 gpc845 (
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21], stage1_30[22], stage1_30[23]},
      {stage2_32[3],stage2_31[3],stage2_30[4],stage2_29[11],stage2_28[19]}
   );
   gpc606_5 gpc846 (
      {stage1_28[30], stage1_28[31], stage1_28[32], stage1_28[33], stage1_28[34], stage1_28[35]},
      {stage1_30[24], stage1_30[25], stage1_30[26], stage1_30[27], stage1_30[28], stage1_30[29]},
      {stage2_32[4],stage2_31[4],stage2_30[5],stage2_29[12],stage2_28[20]}
   );
   gpc606_5 gpc847 (
      {stage1_28[36], stage1_28[37], stage1_28[38], stage1_28[39], stage1_28[40], stage1_28[41]},
      {stage1_30[30], stage1_30[31], stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35]},
      {stage2_32[5],stage2_31[5],stage2_30[6],stage2_29[13],stage2_28[21]}
   );
   gpc606_5 gpc848 (
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[6],stage2_31[6],stage2_30[7],stage2_29[14]}
   );
   gpc606_5 gpc849 (
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[7],stage2_31[7],stage2_30[8],stage2_29[15]}
   );
   gpc606_5 gpc850 (
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[8],stage2_31[8],stage2_30[9],stage2_29[16]}
   );
   gpc606_5 gpc851 (
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage1_31[18], stage1_31[19], stage1_31[20], stage1_31[21], stage1_31[22], stage1_31[23]},
      {stage2_33[3],stage2_32[9],stage2_31[9],stage2_30[10],stage2_29[17]}
   );
   gpc606_5 gpc852 (
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage1_31[24], stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29]},
      {stage2_33[4],stage2_32[10],stage2_31[10],stage2_30[11],stage2_29[18]}
   );
   gpc606_5 gpc853 (
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage1_31[30], stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35]},
      {stage2_33[5],stage2_32[11],stage2_31[11],stage2_30[12],stage2_29[19]}
   );
   gpc606_5 gpc854 (
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage1_31[36], stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41]},
      {stage2_33[6],stage2_32[12],stage2_31[12],stage2_30[13],stage2_29[20]}
   );
   gpc1325_5 gpc855 (
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46]},
      {stage1_30[36], stage1_30[37]},
      {stage1_31[42], stage1_31[43], stage1_31[44]},
      {stage1_32[0]},
      {stage2_33[7],stage2_32[13],stage2_31[13],stage2_30[14],stage2_29[21]}
   );
   gpc606_5 gpc856 (
      {stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41], stage1_30[42], stage1_30[43]},
      {stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5], stage1_32[6]},
      {stage2_34[0],stage2_33[8],stage2_32[14],stage2_31[14],stage2_30[15]}
   );
   gpc606_5 gpc857 (
      {stage1_30[44], stage1_30[45], stage1_30[46], stage1_30[47], stage1_30[48], stage1_30[49]},
      {stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11], stage1_32[12]},
      {stage2_34[1],stage2_33[9],stage2_32[15],stage2_31[15],stage2_30[16]}
   );
   gpc606_5 gpc858 (
      {stage1_30[50], stage1_30[51], stage1_30[52], stage1_30[53], stage1_30[54], stage1_30[55]},
      {stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17], stage1_32[18]},
      {stage2_34[2],stage2_33[10],stage2_32[16],stage2_31[16],stage2_30[17]}
   );
   gpc606_5 gpc859 (
      {stage1_30[56], stage1_30[57], stage1_30[58], stage1_30[59], stage1_30[60], 1'b0},
      {stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23], stage1_32[24]},
      {stage2_34[3],stage2_33[11],stage2_32[17],stage2_31[17],stage2_30[18]}
   );
   gpc606_5 gpc860 (
      {stage1_31[45], stage1_31[46], stage1_31[47], stage1_31[48], stage1_31[49], stage1_31[50]},
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5]},
      {stage2_35[0],stage2_34[4],stage2_33[12],stage2_32[18],stage2_31[18]}
   );
   gpc606_5 gpc861 (
      {stage1_31[51], stage1_31[52], stage1_31[53], stage1_31[54], stage1_31[55], stage1_31[56]},
      {stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11]},
      {stage2_35[1],stage2_34[5],stage2_33[13],stage2_32[19],stage2_31[19]}
   );
   gpc1_1 gpc862 (
      {stage1_0[0]},
      {stage2_0[0]}
   );
   gpc1_1 gpc863 (
      {stage1_0[1]},
      {stage2_0[1]}
   );
   gpc1_1 gpc864 (
      {stage1_0[2]},
      {stage2_0[2]}
   );
   gpc1_1 gpc865 (
      {stage1_0[3]},
      {stage2_0[3]}
   );
   gpc1_1 gpc866 (
      {stage1_0[4]},
      {stage2_0[4]}
   );
   gpc1_1 gpc867 (
      {stage1_0[5]},
      {stage2_0[5]}
   );
   gpc1_1 gpc868 (
      {stage1_0[6]},
      {stage2_0[6]}
   );
   gpc1_1 gpc869 (
      {stage1_0[7]},
      {stage2_0[7]}
   );
   gpc1_1 gpc870 (
      {stage1_0[8]},
      {stage2_0[8]}
   );
   gpc1_1 gpc871 (
      {stage1_0[9]},
      {stage2_0[9]}
   );
   gpc1_1 gpc872 (
      {stage1_0[10]},
      {stage2_0[10]}
   );
   gpc1_1 gpc873 (
      {stage1_0[11]},
      {stage2_0[11]}
   );
   gpc1_1 gpc874 (
      {stage1_0[12]},
      {stage2_0[12]}
   );
   gpc1_1 gpc875 (
      {stage1_0[13]},
      {stage2_0[13]}
   );
   gpc1_1 gpc876 (
      {stage1_0[14]},
      {stage2_0[14]}
   );
   gpc1_1 gpc877 (
      {stage1_0[15]},
      {stage2_0[15]}
   );
   gpc1_1 gpc878 (
      {stage1_0[16]},
      {stage2_0[16]}
   );
   gpc1_1 gpc879 (
      {stage1_0[17]},
      {stage2_0[17]}
   );
   gpc1_1 gpc880 (
      {stage1_0[18]},
      {stage2_0[18]}
   );
   gpc1_1 gpc881 (
      {stage1_0[19]},
      {stage2_0[19]}
   );
   gpc1_1 gpc882 (
      {stage1_0[20]},
      {stage2_0[20]}
   );
   gpc1_1 gpc883 (
      {stage1_0[21]},
      {stage2_0[21]}
   );
   gpc1_1 gpc884 (
      {stage1_0[22]},
      {stage2_0[22]}
   );
   gpc1_1 gpc885 (
      {stage1_0[23]},
      {stage2_0[23]}
   );
   gpc1_1 gpc886 (
      {stage1_0[24]},
      {stage2_0[24]}
   );
   gpc1_1 gpc887 (
      {stage1_0[25]},
      {stage2_0[25]}
   );
   gpc1_1 gpc888 (
      {stage1_0[26]},
      {stage2_0[26]}
   );
   gpc1_1 gpc889 (
      {stage1_0[27]},
      {stage2_0[27]}
   );
   gpc1_1 gpc890 (
      {stage1_0[28]},
      {stage2_0[28]}
   );
   gpc1_1 gpc891 (
      {stage1_0[29]},
      {stage2_0[29]}
   );
   gpc1_1 gpc892 (
      {stage1_0[30]},
      {stage2_0[30]}
   );
   gpc1_1 gpc893 (
      {stage1_0[31]},
      {stage2_0[31]}
   );
   gpc1_1 gpc894 (
      {stage1_0[32]},
      {stage2_0[32]}
   );
   gpc1_1 gpc895 (
      {stage1_0[33]},
      {stage2_0[33]}
   );
   gpc1_1 gpc896 (
      {stage1_0[34]},
      {stage2_0[34]}
   );
   gpc1_1 gpc897 (
      {stage1_0[35]},
      {stage2_0[35]}
   );
   gpc1_1 gpc898 (
      {stage1_1[24]},
      {stage2_1[4]}
   );
   gpc1_1 gpc899 (
      {stage1_1[25]},
      {stage2_1[5]}
   );
   gpc1_1 gpc900 (
      {stage1_1[26]},
      {stage2_1[6]}
   );
   gpc1_1 gpc901 (
      {stage1_1[27]},
      {stage2_1[7]}
   );
   gpc1_1 gpc902 (
      {stage1_1[28]},
      {stage2_1[8]}
   );
   gpc1_1 gpc903 (
      {stage1_1[29]},
      {stage2_1[9]}
   );
   gpc1_1 gpc904 (
      {stage1_1[30]},
      {stage2_1[10]}
   );
   gpc1_1 gpc905 (
      {stage1_1[31]},
      {stage2_1[11]}
   );
   gpc1_1 gpc906 (
      {stage1_1[32]},
      {stage2_1[12]}
   );
   gpc1_1 gpc907 (
      {stage1_1[33]},
      {stage2_1[13]}
   );
   gpc1_1 gpc908 (
      {stage1_1[34]},
      {stage2_1[14]}
   );
   gpc1_1 gpc909 (
      {stage1_1[35]},
      {stage2_1[15]}
   );
   gpc1_1 gpc910 (
      {stage1_1[36]},
      {stage2_1[16]}
   );
   gpc1_1 gpc911 (
      {stage1_1[37]},
      {stage2_1[17]}
   );
   gpc1_1 gpc912 (
      {stage1_1[38]},
      {stage2_1[18]}
   );
   gpc1_1 gpc913 (
      {stage1_1[39]},
      {stage2_1[19]}
   );
   gpc1_1 gpc914 (
      {stage1_2[43]},
      {stage2_2[12]}
   );
   gpc1_1 gpc915 (
      {stage1_2[44]},
      {stage2_2[13]}
   );
   gpc1_1 gpc916 (
      {stage1_2[45]},
      {stage2_2[14]}
   );
   gpc1_1 gpc917 (
      {stage1_2[46]},
      {stage2_2[15]}
   );
   gpc1_1 gpc918 (
      {stage1_2[47]},
      {stage2_2[16]}
   );
   gpc1_1 gpc919 (
      {stage1_2[48]},
      {stage2_2[17]}
   );
   gpc1_1 gpc920 (
      {stage1_2[49]},
      {stage2_2[18]}
   );
   gpc1_1 gpc921 (
      {stage1_2[50]},
      {stage2_2[19]}
   );
   gpc1_1 gpc922 (
      {stage1_2[51]},
      {stage2_2[20]}
   );
   gpc1_1 gpc923 (
      {stage1_2[52]},
      {stage2_2[21]}
   );
   gpc1_1 gpc924 (
      {stage1_2[53]},
      {stage2_2[22]}
   );
   gpc1_1 gpc925 (
      {stage1_2[54]},
      {stage2_2[23]}
   );
   gpc1_1 gpc926 (
      {stage1_2[55]},
      {stage2_2[24]}
   );
   gpc1_1 gpc927 (
      {stage1_2[56]},
      {stage2_2[25]}
   );
   gpc1_1 gpc928 (
      {stage1_2[57]},
      {stage2_2[26]}
   );
   gpc1_1 gpc929 (
      {stage1_3[39]},
      {stage2_3[14]}
   );
   gpc1_1 gpc930 (
      {stage1_3[40]},
      {stage2_3[15]}
   );
   gpc1_1 gpc931 (
      {stage1_3[41]},
      {stage2_3[16]}
   );
   gpc1_1 gpc932 (
      {stage1_3[42]},
      {stage2_3[17]}
   );
   gpc1_1 gpc933 (
      {stage1_3[43]},
      {stage2_3[18]}
   );
   gpc1_1 gpc934 (
      {stage1_3[44]},
      {stage2_3[19]}
   );
   gpc1_1 gpc935 (
      {stage1_3[45]},
      {stage2_3[20]}
   );
   gpc1_1 gpc936 (
      {stage1_3[46]},
      {stage2_3[21]}
   );
   gpc1_1 gpc937 (
      {stage1_3[47]},
      {stage2_3[22]}
   );
   gpc1_1 gpc938 (
      {stage1_3[48]},
      {stage2_3[23]}
   );
   gpc1_1 gpc939 (
      {stage1_3[49]},
      {stage2_3[24]}
   );
   gpc1_1 gpc940 (
      {stage1_3[50]},
      {stage2_3[25]}
   );
   gpc1_1 gpc941 (
      {stage1_3[51]},
      {stage2_3[26]}
   );
   gpc1_1 gpc942 (
      {stage1_3[52]},
      {stage2_3[27]}
   );
   gpc1_1 gpc943 (
      {stage1_3[53]},
      {stage2_3[28]}
   );
   gpc1_1 gpc944 (
      {stage1_3[54]},
      {stage2_3[29]}
   );
   gpc1_1 gpc945 (
      {stage1_3[55]},
      {stage2_3[30]}
   );
   gpc1_1 gpc946 (
      {stage1_3[56]},
      {stage2_3[31]}
   );
   gpc1_1 gpc947 (
      {stage1_3[57]},
      {stage2_3[32]}
   );
   gpc1_1 gpc948 (
      {stage1_3[58]},
      {stage2_3[33]}
   );
   gpc1_1 gpc949 (
      {stage1_4[56]},
      {stage2_4[15]}
   );
   gpc1_1 gpc950 (
      {stage1_4[57]},
      {stage2_4[16]}
   );
   gpc1_1 gpc951 (
      {stage1_4[58]},
      {stage2_4[17]}
   );
   gpc1_1 gpc952 (
      {stage1_4[59]},
      {stage2_4[18]}
   );
   gpc1_1 gpc953 (
      {stage1_4[60]},
      {stage2_4[19]}
   );
   gpc1_1 gpc954 (
      {stage1_4[61]},
      {stage2_4[20]}
   );
   gpc1_1 gpc955 (
      {stage1_4[62]},
      {stage2_4[21]}
   );
   gpc1_1 gpc956 (
      {stage1_4[63]},
      {stage2_4[22]}
   );
   gpc1_1 gpc957 (
      {stage1_4[64]},
      {stage2_4[23]}
   );
   gpc1_1 gpc958 (
      {stage1_4[65]},
      {stage2_4[24]}
   );
   gpc1_1 gpc959 (
      {stage1_4[66]},
      {stage2_4[25]}
   );
   gpc1_1 gpc960 (
      {stage1_5[54]},
      {stage2_5[22]}
   );
   gpc1_1 gpc961 (
      {stage1_5[55]},
      {stage2_5[23]}
   );
   gpc1_1 gpc962 (
      {stage1_5[56]},
      {stage2_5[24]}
   );
   gpc1_1 gpc963 (
      {stage1_5[57]},
      {stage2_5[25]}
   );
   gpc1_1 gpc964 (
      {stage1_5[58]},
      {stage2_5[26]}
   );
   gpc1_1 gpc965 (
      {stage1_5[59]},
      {stage2_5[27]}
   );
   gpc1_1 gpc966 (
      {stage1_5[60]},
      {stage2_5[28]}
   );
   gpc1_1 gpc967 (
      {stage1_5[61]},
      {stage2_5[29]}
   );
   gpc1_1 gpc968 (
      {stage1_5[62]},
      {stage2_5[30]}
   );
   gpc1_1 gpc969 (
      {stage1_6[23]},
      {stage2_6[21]}
   );
   gpc1_1 gpc970 (
      {stage1_6[24]},
      {stage2_6[22]}
   );
   gpc1_1 gpc971 (
      {stage1_6[25]},
      {stage2_6[23]}
   );
   gpc1_1 gpc972 (
      {stage1_6[26]},
      {stage2_6[24]}
   );
   gpc1_1 gpc973 (
      {stage1_6[27]},
      {stage2_6[25]}
   );
   gpc1_1 gpc974 (
      {stage1_6[28]},
      {stage2_6[26]}
   );
   gpc1_1 gpc975 (
      {stage1_6[29]},
      {stage2_6[27]}
   );
   gpc1_1 gpc976 (
      {stage1_6[30]},
      {stage2_6[28]}
   );
   gpc1_1 gpc977 (
      {stage1_6[31]},
      {stage2_6[29]}
   );
   gpc1_1 gpc978 (
      {stage1_6[32]},
      {stage2_6[30]}
   );
   gpc1_1 gpc979 (
      {stage1_6[33]},
      {stage2_6[31]}
   );
   gpc1_1 gpc980 (
      {stage1_6[34]},
      {stage2_6[32]}
   );
   gpc1_1 gpc981 (
      {stage1_6[35]},
      {stage2_6[33]}
   );
   gpc1_1 gpc982 (
      {stage1_6[36]},
      {stage2_6[34]}
   );
   gpc1_1 gpc983 (
      {stage1_6[37]},
      {stage2_6[35]}
   );
   gpc1_1 gpc984 (
      {stage1_6[38]},
      {stage2_6[36]}
   );
   gpc1_1 gpc985 (
      {stage1_6[39]},
      {stage2_6[37]}
   );
   gpc1_1 gpc986 (
      {stage1_6[40]},
      {stage2_6[38]}
   );
   gpc1_1 gpc987 (
      {stage1_6[41]},
      {stage2_6[39]}
   );
   gpc1_1 gpc988 (
      {stage1_6[42]},
      {stage2_6[40]}
   );
   gpc1_1 gpc989 (
      {stage1_6[43]},
      {stage2_6[41]}
   );
   gpc1_1 gpc990 (
      {stage1_6[44]},
      {stage2_6[42]}
   );
   gpc1_1 gpc991 (
      {stage1_6[45]},
      {stage2_6[43]}
   );
   gpc1_1 gpc992 (
      {stage1_6[46]},
      {stage2_6[44]}
   );
   gpc1_1 gpc993 (
      {stage1_6[47]},
      {stage2_6[45]}
   );
   gpc1_1 gpc994 (
      {stage1_6[48]},
      {stage2_6[46]}
   );
   gpc1_1 gpc995 (
      {stage1_6[49]},
      {stage2_6[47]}
   );
   gpc1_1 gpc996 (
      {stage1_7[68]},
      {stage2_7[18]}
   );
   gpc1_1 gpc997 (
      {stage1_7[69]},
      {stage2_7[19]}
   );
   gpc1_1 gpc998 (
      {stage1_8[35]},
      {stage2_8[18]}
   );
   gpc1_1 gpc999 (
      {stage1_8[36]},
      {stage2_8[19]}
   );
   gpc1_1 gpc1000 (
      {stage1_8[37]},
      {stage2_8[20]}
   );
   gpc1_1 gpc1001 (
      {stage1_8[38]},
      {stage2_8[21]}
   );
   gpc1_1 gpc1002 (
      {stage1_8[39]},
      {stage2_8[22]}
   );
   gpc1_1 gpc1003 (
      {stage1_8[40]},
      {stage2_8[23]}
   );
   gpc1_1 gpc1004 (
      {stage1_8[41]},
      {stage2_8[24]}
   );
   gpc1_1 gpc1005 (
      {stage1_8[42]},
      {stage2_8[25]}
   );
   gpc1_1 gpc1006 (
      {stage1_8[43]},
      {stage2_8[26]}
   );
   gpc1_1 gpc1007 (
      {stage1_8[44]},
      {stage2_8[27]}
   );
   gpc1_1 gpc1008 (
      {stage1_8[45]},
      {stage2_8[28]}
   );
   gpc1_1 gpc1009 (
      {stage1_8[46]},
      {stage2_8[29]}
   );
   gpc1_1 gpc1010 (
      {stage1_8[47]},
      {stage2_8[30]}
   );
   gpc1_1 gpc1011 (
      {stage1_8[48]},
      {stage2_8[31]}
   );
   gpc1_1 gpc1012 (
      {stage1_8[49]},
      {stage2_8[32]}
   );
   gpc1_1 gpc1013 (
      {stage1_8[50]},
      {stage2_8[33]}
   );
   gpc1_1 gpc1014 (
      {stage1_8[51]},
      {stage2_8[34]}
   );
   gpc1_1 gpc1015 (
      {stage1_8[52]},
      {stage2_8[35]}
   );
   gpc1_1 gpc1016 (
      {stage1_8[53]},
      {stage2_8[36]}
   );
   gpc1_1 gpc1017 (
      {stage1_8[54]},
      {stage2_8[37]}
   );
   gpc1_1 gpc1018 (
      {stage1_8[55]},
      {stage2_8[38]}
   );
   gpc1_1 gpc1019 (
      {stage1_9[60]},
      {stage2_9[22]}
   );
   gpc1_1 gpc1020 (
      {stage1_11[55]},
      {stage2_11[24]}
   );
   gpc1_1 gpc1021 (
      {stage1_11[56]},
      {stage2_11[25]}
   );
   gpc1_1 gpc1022 (
      {stage1_11[57]},
      {stage2_11[26]}
   );
   gpc1_1 gpc1023 (
      {stage1_13[48]},
      {stage2_13[22]}
   );
   gpc1_1 gpc1024 (
      {stage1_13[49]},
      {stage2_13[23]}
   );
   gpc1_1 gpc1025 (
      {stage1_13[50]},
      {stage2_13[24]}
   );
   gpc1_1 gpc1026 (
      {stage1_13[51]},
      {stage2_13[25]}
   );
   gpc1_1 gpc1027 (
      {stage1_13[52]},
      {stage2_13[26]}
   );
   gpc1_1 gpc1028 (
      {stage1_13[53]},
      {stage2_13[27]}
   );
   gpc1_1 gpc1029 (
      {stage1_13[54]},
      {stage2_13[28]}
   );
   gpc1_1 gpc1030 (
      {stage1_13[55]},
      {stage2_13[29]}
   );
   gpc1_1 gpc1031 (
      {stage1_13[56]},
      {stage2_13[30]}
   );
   gpc1_1 gpc1032 (
      {stage1_13[57]},
      {stage2_13[31]}
   );
   gpc1_1 gpc1033 (
      {stage1_13[58]},
      {stage2_13[32]}
   );
   gpc1_1 gpc1034 (
      {stage1_13[59]},
      {stage2_13[33]}
   );
   gpc1_1 gpc1035 (
      {stage1_13[60]},
      {stage2_13[34]}
   );
   gpc1_1 gpc1036 (
      {stage1_14[42]},
      {stage2_14[23]}
   );
   gpc1_1 gpc1037 (
      {stage1_14[43]},
      {stage2_14[24]}
   );
   gpc1_1 gpc1038 (
      {stage1_14[44]},
      {stage2_14[25]}
   );
   gpc1_1 gpc1039 (
      {stage1_14[45]},
      {stage2_14[26]}
   );
   gpc1_1 gpc1040 (
      {stage1_15[44]},
      {stage2_15[20]}
   );
   gpc1_1 gpc1041 (
      {stage1_15[45]},
      {stage2_15[21]}
   );
   gpc1_1 gpc1042 (
      {stage1_15[46]},
      {stage2_15[22]}
   );
   gpc1_1 gpc1043 (
      {stage1_17[37]},
      {stage2_17[23]}
   );
   gpc1_1 gpc1044 (
      {stage1_17[38]},
      {stage2_17[24]}
   );
   gpc1_1 gpc1045 (
      {stage1_17[39]},
      {stage2_17[25]}
   );
   gpc1_1 gpc1046 (
      {stage1_17[40]},
      {stage2_17[26]}
   );
   gpc1_1 gpc1047 (
      {stage1_17[41]},
      {stage2_17[27]}
   );
   gpc1_1 gpc1048 (
      {stage1_17[42]},
      {stage2_17[28]}
   );
   gpc1_1 gpc1049 (
      {stage1_17[43]},
      {stage2_17[29]}
   );
   gpc1_1 gpc1050 (
      {stage1_17[44]},
      {stage2_17[30]}
   );
   gpc1_1 gpc1051 (
      {stage1_17[45]},
      {stage2_17[31]}
   );
   gpc1_1 gpc1052 (
      {stage1_17[46]},
      {stage2_17[32]}
   );
   gpc1_1 gpc1053 (
      {stage1_17[47]},
      {stage2_17[33]}
   );
   gpc1_1 gpc1054 (
      {stage1_17[48]},
      {stage2_17[34]}
   );
   gpc1_1 gpc1055 (
      {stage1_17[49]},
      {stage2_17[35]}
   );
   gpc1_1 gpc1056 (
      {stage1_17[50]},
      {stage2_17[36]}
   );
   gpc1_1 gpc1057 (
      {stage1_17[51]},
      {stage2_17[37]}
   );
   gpc1_1 gpc1058 (
      {stage1_17[52]},
      {stage2_17[38]}
   );
   gpc1_1 gpc1059 (
      {stage1_17[53]},
      {stage2_17[39]}
   );
   gpc1_1 gpc1060 (
      {stage1_17[54]},
      {stage2_17[40]}
   );
   gpc1_1 gpc1061 (
      {stage1_17[55]},
      {stage2_17[41]}
   );
   gpc1_1 gpc1062 (
      {stage1_17[56]},
      {stage2_17[42]}
   );
   gpc1_1 gpc1063 (
      {stage1_17[57]},
      {stage2_17[43]}
   );
   gpc1_1 gpc1064 (
      {stage1_17[58]},
      {stage2_17[44]}
   );
   gpc1_1 gpc1065 (
      {stage1_17[59]},
      {stage2_17[45]}
   );
   gpc1_1 gpc1066 (
      {stage1_17[60]},
      {stage2_17[46]}
   );
   gpc1_1 gpc1067 (
      {stage1_17[61]},
      {stage2_17[47]}
   );
   gpc1_1 gpc1068 (
      {stage1_17[62]},
      {stage2_17[48]}
   );
   gpc1_1 gpc1069 (
      {stage1_18[48]},
      {stage2_18[20]}
   );
   gpc1_1 gpc1070 (
      {stage1_18[49]},
      {stage2_18[21]}
   );
   gpc1_1 gpc1071 (
      {stage1_18[50]},
      {stage2_18[22]}
   );
   gpc1_1 gpc1072 (
      {stage1_18[51]},
      {stage2_18[23]}
   );
   gpc1_1 gpc1073 (
      {stage1_18[52]},
      {stage2_18[24]}
   );
   gpc1_1 gpc1074 (
      {stage1_18[53]},
      {stage2_18[25]}
   );
   gpc1_1 gpc1075 (
      {stage1_18[54]},
      {stage2_18[26]}
   );
   gpc1_1 gpc1076 (
      {stage1_18[55]},
      {stage2_18[27]}
   );
   gpc1_1 gpc1077 (
      {stage1_18[56]},
      {stage2_18[28]}
   );
   gpc1_1 gpc1078 (
      {stage1_18[57]},
      {stage2_18[29]}
   );
   gpc1_1 gpc1079 (
      {stage1_18[58]},
      {stage2_18[30]}
   );
   gpc1_1 gpc1080 (
      {stage1_18[59]},
      {stage2_18[31]}
   );
   gpc1_1 gpc1081 (
      {stage1_18[60]},
      {stage2_18[32]}
   );
   gpc1_1 gpc1082 (
      {stage1_18[61]},
      {stage2_18[33]}
   );
   gpc1_1 gpc1083 (
      {stage1_18[62]},
      {stage2_18[34]}
   );
   gpc1_1 gpc1084 (
      {stage1_18[63]},
      {stage2_18[35]}
   );
   gpc1_1 gpc1085 (
      {stage1_18[64]},
      {stage2_18[36]}
   );
   gpc1_1 gpc1086 (
      {stage1_18[65]},
      {stage2_18[37]}
   );
   gpc1_1 gpc1087 (
      {stage1_19[42]},
      {stage2_19[20]}
   );
   gpc1_1 gpc1088 (
      {stage1_20[30]},
      {stage2_20[20]}
   );
   gpc1_1 gpc1089 (
      {stage1_20[31]},
      {stage2_20[21]}
   );
   gpc1_1 gpc1090 (
      {stage1_20[32]},
      {stage2_20[22]}
   );
   gpc1_1 gpc1091 (
      {stage1_20[33]},
      {stage2_20[23]}
   );
   gpc1_1 gpc1092 (
      {stage1_20[34]},
      {stage2_20[24]}
   );
   gpc1_1 gpc1093 (
      {stage1_20[35]},
      {stage2_20[25]}
   );
   gpc1_1 gpc1094 (
      {stage1_20[36]},
      {stage2_20[26]}
   );
   gpc1_1 gpc1095 (
      {stage1_20[37]},
      {stage2_20[27]}
   );
   gpc1_1 gpc1096 (
      {stage1_20[38]},
      {stage2_20[28]}
   );
   gpc1_1 gpc1097 (
      {stage1_20[39]},
      {stage2_20[29]}
   );
   gpc1_1 gpc1098 (
      {stage1_20[40]},
      {stage2_20[30]}
   );
   gpc1_1 gpc1099 (
      {stage1_20[41]},
      {stage2_20[31]}
   );
   gpc1_1 gpc1100 (
      {stage1_20[42]},
      {stage2_20[32]}
   );
   gpc1_1 gpc1101 (
      {stage1_20[43]},
      {stage2_20[33]}
   );
   gpc1_1 gpc1102 (
      {stage1_20[44]},
      {stage2_20[34]}
   );
   gpc1_1 gpc1103 (
      {stage1_20[45]},
      {stage2_20[35]}
   );
   gpc1_1 gpc1104 (
      {stage1_20[46]},
      {stage2_20[36]}
   );
   gpc1_1 gpc1105 (
      {stage1_20[47]},
      {stage2_20[37]}
   );
   gpc1_1 gpc1106 (
      {stage1_20[48]},
      {stage2_20[38]}
   );
   gpc1_1 gpc1107 (
      {stage1_20[49]},
      {stage2_20[39]}
   );
   gpc1_1 gpc1108 (
      {stage1_20[50]},
      {stage2_20[40]}
   );
   gpc1_1 gpc1109 (
      {stage1_20[51]},
      {stage2_20[41]}
   );
   gpc1_1 gpc1110 (
      {stage1_20[52]},
      {stage2_20[42]}
   );
   gpc1_1 gpc1111 (
      {stage1_20[53]},
      {stage2_20[43]}
   );
   gpc1_1 gpc1112 (
      {stage1_20[54]},
      {stage2_20[44]}
   );
   gpc1_1 gpc1113 (
      {stage1_20[55]},
      {stage2_20[45]}
   );
   gpc1_1 gpc1114 (
      {stage1_20[56]},
      {stage2_20[46]}
   );
   gpc1_1 gpc1115 (
      {stage1_20[57]},
      {stage2_20[47]}
   );
   gpc1_1 gpc1116 (
      {stage1_20[58]},
      {stage2_20[48]}
   );
   gpc1_1 gpc1117 (
      {stage1_20[59]},
      {stage2_20[49]}
   );
   gpc1_1 gpc1118 (
      {stage1_20[60]},
      {stage2_20[50]}
   );
   gpc1_1 gpc1119 (
      {stage1_20[61]},
      {stage2_20[51]}
   );
   gpc1_1 gpc1120 (
      {stage1_20[62]},
      {stage2_20[52]}
   );
   gpc1_1 gpc1121 (
      {stage1_20[63]},
      {stage2_20[53]}
   );
   gpc1_1 gpc1122 (
      {stage1_20[64]},
      {stage2_20[54]}
   );
   gpc1_1 gpc1123 (
      {stage1_20[65]},
      {stage2_20[55]}
   );
   gpc1_1 gpc1124 (
      {stage1_21[60]},
      {stage2_21[16]}
   );
   gpc1_1 gpc1125 (
      {stage1_21[61]},
      {stage2_21[17]}
   );
   gpc1_1 gpc1126 (
      {stage1_21[62]},
      {stage2_21[18]}
   );
   gpc1_1 gpc1127 (
      {stage1_21[63]},
      {stage2_21[19]}
   );
   gpc1_1 gpc1128 (
      {stage1_21[64]},
      {stage2_21[20]}
   );
   gpc1_1 gpc1129 (
      {stage1_22[53]},
      {stage2_22[19]}
   );
   gpc1_1 gpc1130 (
      {stage1_22[54]},
      {stage2_22[20]}
   );
   gpc1_1 gpc1131 (
      {stage1_22[55]},
      {stage2_22[21]}
   );
   gpc1_1 gpc1132 (
      {stage1_22[56]},
      {stage2_22[22]}
   );
   gpc1_1 gpc1133 (
      {stage1_22[57]},
      {stage2_22[23]}
   );
   gpc1_1 gpc1134 (
      {stage1_22[58]},
      {stage2_22[24]}
   );
   gpc1_1 gpc1135 (
      {stage1_22[59]},
      {stage2_22[25]}
   );
   gpc1_1 gpc1136 (
      {stage1_22[60]},
      {stage2_22[26]}
   );
   gpc1_1 gpc1137 (
      {stage1_23[30]},
      {stage2_23[20]}
   );
   gpc1_1 gpc1138 (
      {stage1_23[31]},
      {stage2_23[21]}
   );
   gpc1_1 gpc1139 (
      {stage1_23[32]},
      {stage2_23[22]}
   );
   gpc1_1 gpc1140 (
      {stage1_23[33]},
      {stage2_23[23]}
   );
   gpc1_1 gpc1141 (
      {stage1_23[34]},
      {stage2_23[24]}
   );
   gpc1_1 gpc1142 (
      {stage1_23[35]},
      {stage2_23[25]}
   );
   gpc1_1 gpc1143 (
      {stage1_23[36]},
      {stage2_23[26]}
   );
   gpc1_1 gpc1144 (
      {stage1_23[37]},
      {stage2_23[27]}
   );
   gpc1_1 gpc1145 (
      {stage1_23[38]},
      {stage2_23[28]}
   );
   gpc1_1 gpc1146 (
      {stage1_23[39]},
      {stage2_23[29]}
   );
   gpc1_1 gpc1147 (
      {stage1_23[40]},
      {stage2_23[30]}
   );
   gpc1_1 gpc1148 (
      {stage1_23[41]},
      {stage2_23[31]}
   );
   gpc1_1 gpc1149 (
      {stage1_23[42]},
      {stage2_23[32]}
   );
   gpc1_1 gpc1150 (
      {stage1_23[43]},
      {stage2_23[33]}
   );
   gpc1_1 gpc1151 (
      {stage1_24[79]},
      {stage2_24[22]}
   );
   gpc1_1 gpc1152 (
      {stage1_24[80]},
      {stage2_24[23]}
   );
   gpc1_1 gpc1153 (
      {stage1_24[81]},
      {stage2_24[24]}
   );
   gpc1_1 gpc1154 (
      {stage1_24[82]},
      {stage2_24[25]}
   );
   gpc1_1 gpc1155 (
      {stage1_24[83]},
      {stage2_24[26]}
   );
   gpc1_1 gpc1156 (
      {stage1_24[84]},
      {stage2_24[27]}
   );
   gpc1_1 gpc1157 (
      {stage1_24[85]},
      {stage2_24[28]}
   );
   gpc1_1 gpc1158 (
      {stage1_24[86]},
      {stage2_24[29]}
   );
   gpc1_1 gpc1159 (
      {stage1_24[87]},
      {stage2_24[30]}
   );
   gpc1_1 gpc1160 (
      {stage1_24[88]},
      {stage2_24[31]}
   );
   gpc1_1 gpc1161 (
      {stage1_24[89]},
      {stage2_24[32]}
   );
   gpc1_1 gpc1162 (
      {stage1_25[48]},
      {stage2_25[25]}
   );
   gpc1_1 gpc1163 (
      {stage1_25[49]},
      {stage2_25[26]}
   );
   gpc1_1 gpc1164 (
      {stage1_25[50]},
      {stage2_25[27]}
   );
   gpc1_1 gpc1165 (
      {stage1_25[51]},
      {stage2_25[28]}
   );
   gpc1_1 gpc1166 (
      {stage1_25[52]},
      {stage2_25[29]}
   );
   gpc1_1 gpc1167 (
      {stage1_25[53]},
      {stage2_25[30]}
   );
   gpc1_1 gpc1168 (
      {stage1_25[54]},
      {stage2_25[31]}
   );
   gpc1_1 gpc1169 (
      {stage1_25[55]},
      {stage2_25[32]}
   );
   gpc1_1 gpc1170 (
      {stage1_25[56]},
      {stage2_25[33]}
   );
   gpc1_1 gpc1171 (
      {stage1_25[57]},
      {stage2_25[34]}
   );
   gpc1_1 gpc1172 (
      {stage1_25[58]},
      {stage2_25[35]}
   );
   gpc1_1 gpc1173 (
      {stage1_25[59]},
      {stage2_25[36]}
   );
   gpc1_1 gpc1174 (
      {stage1_25[60]},
      {stage2_25[37]}
   );
   gpc1_1 gpc1175 (
      {stage1_25[61]},
      {stage2_25[38]}
   );
   gpc1_1 gpc1176 (
      {stage1_25[62]},
      {stage2_25[39]}
   );
   gpc1_1 gpc1177 (
      {stage1_25[63]},
      {stage2_25[40]}
   );
   gpc1_1 gpc1178 (
      {stage1_25[64]},
      {stage2_25[41]}
   );
   gpc1_1 gpc1179 (
      {stage1_25[65]},
      {stage2_25[42]}
   );
   gpc1_1 gpc1180 (
      {stage1_25[66]},
      {stage2_25[43]}
   );
   gpc1_1 gpc1181 (
      {stage1_25[67]},
      {stage2_25[44]}
   );
   gpc1_1 gpc1182 (
      {stage1_25[68]},
      {stage2_25[45]}
   );
   gpc1_1 gpc1183 (
      {stage1_25[69]},
      {stage2_25[46]}
   );
   gpc1_1 gpc1184 (
      {stage1_26[54]},
      {stage2_26[22]}
   );
   gpc1_1 gpc1185 (
      {stage1_26[55]},
      {stage2_26[23]}
   );
   gpc1_1 gpc1186 (
      {stage1_26[56]},
      {stage2_26[24]}
   );
   gpc1_1 gpc1187 (
      {stage1_26[57]},
      {stage2_26[25]}
   );
   gpc1_1 gpc1188 (
      {stage1_26[58]},
      {stage2_26[26]}
   );
   gpc1_1 gpc1189 (
      {stage1_26[59]},
      {stage2_26[27]}
   );
   gpc1_1 gpc1190 (
      {stage1_26[60]},
      {stage2_26[28]}
   );
   gpc1_1 gpc1191 (
      {stage1_26[61]},
      {stage2_26[29]}
   );
   gpc1_1 gpc1192 (
      {stage1_26[62]},
      {stage2_26[30]}
   );
   gpc1_1 gpc1193 (
      {stage1_26[63]},
      {stage2_26[31]}
   );
   gpc1_1 gpc1194 (
      {stage1_26[64]},
      {stage2_26[32]}
   );
   gpc1_1 gpc1195 (
      {stage1_26[65]},
      {stage2_26[33]}
   );
   gpc1_1 gpc1196 (
      {stage1_26[66]},
      {stage2_26[34]}
   );
   gpc1_1 gpc1197 (
      {stage1_26[67]},
      {stage2_26[35]}
   );
   gpc1_1 gpc1198 (
      {stage1_26[68]},
      {stage2_26[36]}
   );
   gpc1_1 gpc1199 (
      {stage1_27[42]},
      {stage2_27[17]}
   );
   gpc1_1 gpc1200 (
      {stage1_27[43]},
      {stage2_27[18]}
   );
   gpc1_1 gpc1201 (
      {stage1_27[44]},
      {stage2_27[19]}
   );
   gpc1_1 gpc1202 (
      {stage1_27[45]},
      {stage2_27[20]}
   );
   gpc1_1 gpc1203 (
      {stage1_27[46]},
      {stage2_27[21]}
   );
   gpc1_1 gpc1204 (
      {stage1_27[47]},
      {stage2_27[22]}
   );
   gpc1_1 gpc1205 (
      {stage1_27[48]},
      {stage2_27[23]}
   );
   gpc1_1 gpc1206 (
      {stage1_27[49]},
      {stage2_27[24]}
   );
   gpc1_1 gpc1207 (
      {stage1_27[50]},
      {stage2_27[25]}
   );
   gpc1_1 gpc1208 (
      {stage1_27[51]},
      {stage2_27[26]}
   );
   gpc1_1 gpc1209 (
      {stage1_27[52]},
      {stage2_27[27]}
   );
   gpc1_1 gpc1210 (
      {stage1_27[53]},
      {stage2_27[28]}
   );
   gpc1_1 gpc1211 (
      {stage1_27[54]},
      {stage2_27[29]}
   );
   gpc1_1 gpc1212 (
      {stage1_27[55]},
      {stage2_27[30]}
   );
   gpc1_1 gpc1213 (
      {stage1_28[42]},
      {stage2_28[22]}
   );
   gpc1_1 gpc1214 (
      {stage1_28[43]},
      {stage2_28[23]}
   );
   gpc1_1 gpc1215 (
      {stage1_28[44]},
      {stage2_28[24]}
   );
   gpc1_1 gpc1216 (
      {stage1_28[45]},
      {stage2_28[25]}
   );
   gpc1_1 gpc1217 (
      {stage1_28[46]},
      {stage2_28[26]}
   );
   gpc1_1 gpc1218 (
      {stage1_28[47]},
      {stage2_28[27]}
   );
   gpc1_1 gpc1219 (
      {stage1_28[48]},
      {stage2_28[28]}
   );
   gpc1_1 gpc1220 (
      {stage1_28[49]},
      {stage2_28[29]}
   );
   gpc1_1 gpc1221 (
      {stage1_28[50]},
      {stage2_28[30]}
   );
   gpc1_1 gpc1222 (
      {stage1_28[51]},
      {stage2_28[31]}
   );
   gpc1_1 gpc1223 (
      {stage1_28[52]},
      {stage2_28[32]}
   );
   gpc1_1 gpc1224 (
      {stage1_28[53]},
      {stage2_28[33]}
   );
   gpc1_1 gpc1225 (
      {stage1_28[54]},
      {stage2_28[34]}
   );
   gpc1_1 gpc1226 (
      {stage1_28[55]},
      {stage2_28[35]}
   );
   gpc1_1 gpc1227 (
      {stage1_29[47]},
      {stage2_29[22]}
   );
   gpc1_1 gpc1228 (
      {stage1_29[48]},
      {stage2_29[23]}
   );
   gpc1_1 gpc1229 (
      {stage1_29[49]},
      {stage2_29[24]}
   );
   gpc1_1 gpc1230 (
      {stage1_29[50]},
      {stage2_29[25]}
   );
   gpc1_1 gpc1231 (
      {stage1_29[51]},
      {stage2_29[26]}
   );
   gpc1_1 gpc1232 (
      {stage1_29[52]},
      {stage2_29[27]}
   );
   gpc1_1 gpc1233 (
      {stage1_29[53]},
      {stage2_29[28]}
   );
   gpc1_1 gpc1234 (
      {stage1_29[54]},
      {stage2_29[29]}
   );
   gpc1_1 gpc1235 (
      {stage1_29[55]},
      {stage2_29[30]}
   );
   gpc1_1 gpc1236 (
      {stage1_29[56]},
      {stage2_29[31]}
   );
   gpc1_1 gpc1237 (
      {stage1_31[57]},
      {stage2_31[20]}
   );
   gpc1_1 gpc1238 (
      {stage1_31[58]},
      {stage2_31[21]}
   );
   gpc1_1 gpc1239 (
      {stage1_31[59]},
      {stage2_31[22]}
   );
   gpc1_1 gpc1240 (
      {stage1_31[60]},
      {stage2_31[23]}
   );
   gpc1_1 gpc1241 (
      {stage1_31[61]},
      {stage2_31[24]}
   );
   gpc1_1 gpc1242 (
      {stage1_31[62]},
      {stage2_31[25]}
   );
   gpc1_1 gpc1243 (
      {stage1_31[63]},
      {stage2_31[26]}
   );
   gpc1_1 gpc1244 (
      {stage1_31[64]},
      {stage2_31[27]}
   );
   gpc1_1 gpc1245 (
      {stage1_31[65]},
      {stage2_31[28]}
   );
   gpc1_1 gpc1246 (
      {stage1_31[66]},
      {stage2_31[29]}
   );
   gpc1_1 gpc1247 (
      {stage1_31[67]},
      {stage2_31[30]}
   );
   gpc1_1 gpc1248 (
      {stage1_31[68]},
      {stage2_31[31]}
   );
   gpc1_1 gpc1249 (
      {stage1_31[69]},
      {stage2_31[32]}
   );
   gpc1_1 gpc1250 (
      {stage1_31[70]},
      {stage2_31[33]}
   );
   gpc1_1 gpc1251 (
      {stage1_32[25]},
      {stage2_32[20]}
   );
   gpc1_1 gpc1252 (
      {stage1_32[26]},
      {stage2_32[21]}
   );
   gpc1_1 gpc1253 (
      {stage1_32[27]},
      {stage2_32[22]}
   );
   gpc1_1 gpc1254 (
      {stage1_32[28]},
      {stage2_32[23]}
   );
   gpc1_1 gpc1255 (
      {stage1_32[29]},
      {stage2_32[24]}
   );
   gpc1_1 gpc1256 (
      {stage1_32[30]},
      {stage2_32[25]}
   );
   gpc1_1 gpc1257 (
      {stage1_32[31]},
      {stage2_32[26]}
   );
   gpc1_1 gpc1258 (
      {stage1_32[32]},
      {stage2_32[27]}
   );
   gpc1_1 gpc1259 (
      {stage1_32[33]},
      {stage2_32[28]}
   );
   gpc1_1 gpc1260 (
      {stage1_33[12]},
      {stage2_33[14]}
   );
   gpc1_1 gpc1261 (
      {stage1_33[13]},
      {stage2_33[15]}
   );
   gpc1_1 gpc1262 (
      {stage1_33[14]},
      {stage2_33[16]}
   );
   gpc1_1 gpc1263 (
      {stage1_33[15]},
      {stage2_33[17]}
   );
   gpc2135_5 gpc1264 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[0]},
      {stage2_3[0], stage2_3[1]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc2135_5 gpc1265 (
      {stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8], stage2_0[9]},
      {stage2_1[3], stage2_1[4], stage2_1[5]},
      {stage2_2[1]},
      {stage2_3[2], stage2_3[3]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc2135_5 gpc1266 (
      {stage2_0[10], stage2_0[11], stage2_0[12], stage2_0[13], stage2_0[14]},
      {stage2_1[6], stage2_1[7], stage2_1[8]},
      {stage2_2[2]},
      {stage2_3[4], stage2_3[5]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc2135_5 gpc1267 (
      {stage2_0[15], stage2_0[16], stage2_0[17], stage2_0[18], stage2_0[19]},
      {stage2_1[9], stage2_1[10], stage2_1[11]},
      {stage2_2[3]},
      {stage2_3[6], stage2_3[7]},
      {stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3],stage3_0[3]}
   );
   gpc606_5 gpc1268 (
      {stage2_0[20], stage2_0[21], stage2_0[22], stage2_0[23], stage2_0[24], stage2_0[25]},
      {stage2_2[4], stage2_2[5], stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9]},
      {stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4],stage3_0[4]}
   );
   gpc615_5 gpc1269 (
      {stage2_0[26], stage2_0[27], stage2_0[28], stage2_0[29], stage2_0[30]},
      {stage2_1[12]},
      {stage2_2[10], stage2_2[11], stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15]},
      {stage3_4[5],stage3_3[5],stage3_2[5],stage3_1[5],stage3_0[5]}
   );
   gpc615_5 gpc1270 (
      {stage2_0[31], stage2_0[32], stage2_0[33], stage2_0[34], stage2_0[35]},
      {stage2_1[13]},
      {stage2_2[16], stage2_2[17], stage2_2[18], stage2_2[19], stage2_2[20], stage2_2[21]},
      {stage3_4[6],stage3_3[6],stage3_2[6],stage3_1[6],stage3_0[6]}
   );
   gpc615_5 gpc1271 (
      {stage2_2[22], stage2_2[23], stage2_2[24], stage2_2[25], stage2_2[26]},
      {stage2_3[8]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[0],stage3_4[7],stage3_3[7],stage3_2[7]}
   );
   gpc615_5 gpc1272 (
      {stage2_3[9], stage2_3[10], stage2_3[11], stage2_3[12], stage2_3[13]},
      {stage2_4[6]},
      {stage2_5[0], stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5]},
      {stage3_7[0],stage3_6[1],stage3_5[1],stage3_4[8],stage3_3[8]}
   );
   gpc615_5 gpc1273 (
      {stage2_3[14], stage2_3[15], stage2_3[16], stage2_3[17], stage2_3[18]},
      {stage2_4[7]},
      {stage2_5[6], stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11]},
      {stage3_7[1],stage3_6[2],stage3_5[2],stage3_4[9],stage3_3[9]}
   );
   gpc615_5 gpc1274 (
      {stage2_3[19], stage2_3[20], stage2_3[21], stage2_3[22], stage2_3[23]},
      {stage2_4[8]},
      {stage2_5[12], stage2_5[13], stage2_5[14], stage2_5[15], stage2_5[16], stage2_5[17]},
      {stage3_7[2],stage3_6[3],stage3_5[3],stage3_4[10],stage3_3[10]}
   );
   gpc615_5 gpc1275 (
      {stage2_3[24], stage2_3[25], stage2_3[26], stage2_3[27], stage2_3[28]},
      {stage2_4[9]},
      {stage2_5[18], stage2_5[19], stage2_5[20], stage2_5[21], stage2_5[22], stage2_5[23]},
      {stage3_7[3],stage3_6[4],stage3_5[4],stage3_4[11],stage3_3[11]}
   );
   gpc615_5 gpc1276 (
      {stage2_3[29], stage2_3[30], stage2_3[31], stage2_3[32], stage2_3[33]},
      {stage2_4[10]},
      {stage2_5[24], stage2_5[25], stage2_5[26], stage2_5[27], stage2_5[28], stage2_5[29]},
      {stage3_7[4],stage3_6[5],stage3_5[5],stage3_4[12],stage3_3[12]}
   );
   gpc606_5 gpc1277 (
      {stage2_4[11], stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[5],stage3_6[6],stage3_5[6],stage3_4[13]}
   );
   gpc606_5 gpc1278 (
      {stage2_4[17], stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[6],stage3_6[7],stage3_5[7],stage3_4[14]}
   );
   gpc606_5 gpc1279 (
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[0],stage3_8[2],stage3_7[7],stage3_6[8]}
   );
   gpc606_5 gpc1280 (
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22], stage2_6[23]},
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10], stage2_8[11]},
      {stage3_10[1],stage3_9[1],stage3_8[3],stage3_7[8],stage3_6[9]}
   );
   gpc606_5 gpc1281 (
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[2],stage3_9[2],stage3_8[4],stage3_7[9]}
   );
   gpc615_5 gpc1282 (
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10]},
      {stage2_8[12]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[3],stage3_9[3],stage3_8[5],stage3_7[10]}
   );
   gpc615_5 gpc1283 (
      {stage2_7[11], stage2_7[12], stage2_7[13], stage2_7[14], stage2_7[15]},
      {stage2_8[13]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[4],stage3_9[4],stage3_8[6],stage3_7[11]}
   );
   gpc615_5 gpc1284 (
      {stage2_7[16], stage2_7[17], stage2_7[18], stage2_7[19], 1'b0},
      {stage2_8[14]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], 1'b0},
      {stage3_11[3],stage3_10[5],stage3_9[5],stage3_8[7],stage3_7[12]}
   );
   gpc606_5 gpc1285 (
      {stage2_8[15], stage2_8[16], stage2_8[17], stage2_8[18], stage2_8[19], stage2_8[20]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[4],stage3_10[6],stage3_9[6],stage3_8[8]}
   );
   gpc606_5 gpc1286 (
      {stage2_8[21], stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25], stage2_8[26]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[5],stage3_10[7],stage3_9[7],stage3_8[9]}
   );
   gpc606_5 gpc1287 (
      {stage2_8[27], stage2_8[28], stage2_8[29], stage2_8[30], stage2_8[31], stage2_8[32]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[6],stage3_10[8],stage3_9[8],stage3_8[10]}
   );
   gpc615_5 gpc1288 (
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4]},
      {stage2_12[0]},
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5]},
      {stage3_15[0],stage3_14[0],stage3_13[0],stage3_12[3],stage3_11[7]}
   );
   gpc615_5 gpc1289 (
      {stage2_11[5], stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9]},
      {stage2_12[1]},
      {stage2_13[6], stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11]},
      {stage3_15[1],stage3_14[1],stage3_13[1],stage3_12[4],stage3_11[8]}
   );
   gpc615_5 gpc1290 (
      {stage2_11[10], stage2_11[11], stage2_11[12], stage2_11[13], stage2_11[14]},
      {stage2_12[2]},
      {stage2_13[12], stage2_13[13], stage2_13[14], stage2_13[15], stage2_13[16], stage2_13[17]},
      {stage3_15[2],stage3_14[2],stage3_13[2],stage3_12[5],stage3_11[9]}
   );
   gpc615_5 gpc1291 (
      {stage2_11[15], stage2_11[16], stage2_11[17], stage2_11[18], stage2_11[19]},
      {stage2_12[3]},
      {stage2_13[18], stage2_13[19], stage2_13[20], stage2_13[21], stage2_13[22], stage2_13[23]},
      {stage3_15[3],stage3_14[3],stage3_13[3],stage3_12[6],stage3_11[10]}
   );
   gpc615_5 gpc1292 (
      {stage2_11[20], stage2_11[21], stage2_11[22], stage2_11[23], stage2_11[24]},
      {stage2_12[4]},
      {stage2_13[24], stage2_13[25], stage2_13[26], stage2_13[27], stage2_13[28], stage2_13[29]},
      {stage3_15[4],stage3_14[4],stage3_13[4],stage3_12[7],stage3_11[11]}
   );
   gpc606_5 gpc1293 (
      {stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8], stage2_12[9], stage2_12[10]},
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage3_16[0],stage3_15[5],stage3_14[5],stage3_13[5],stage3_12[8]}
   );
   gpc606_5 gpc1294 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[1],stage3_15[6],stage3_14[6]}
   );
   gpc615_5 gpc1295 (
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4]},
      {stage2_16[6]},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[1],stage3_17[1],stage3_16[2],stage3_15[7]}
   );
   gpc615_5 gpc1296 (
      {stage2_15[5], stage2_15[6], stage2_15[7], stage2_15[8], stage2_15[9]},
      {stage2_16[7]},
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage3_19[1],stage3_18[2],stage3_17[2],stage3_16[3],stage3_15[8]}
   );
   gpc615_5 gpc1297 (
      {stage2_15[10], stage2_15[11], stage2_15[12], stage2_15[13], stage2_15[14]},
      {stage2_16[8]},
      {stage2_17[12], stage2_17[13], stage2_17[14], stage2_17[15], stage2_17[16], stage2_17[17]},
      {stage3_19[2],stage3_18[3],stage3_17[3],stage3_16[4],stage3_15[9]}
   );
   gpc615_5 gpc1298 (
      {stage2_15[15], stage2_15[16], stage2_15[17], stage2_15[18], stage2_15[19]},
      {stage2_16[9]},
      {stage2_17[18], stage2_17[19], stage2_17[20], stage2_17[21], stage2_17[22], stage2_17[23]},
      {stage3_19[3],stage3_18[4],stage3_17[4],stage3_16[5],stage3_15[10]}
   );
   gpc615_5 gpc1299 (
      {stage2_15[20], stage2_15[21], stage2_15[22], 1'b0, 1'b0},
      {stage2_16[10]},
      {stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27], stage2_17[28], stage2_17[29]},
      {stage3_19[4],stage3_18[5],stage3_17[5],stage3_16[6],stage3_15[11]}
   );
   gpc117_4 gpc1300 (
      {stage2_16[11], stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage2_17[30]},
      {stage2_18[0]},
      {stage3_19[5],stage3_18[6],stage3_17[6],stage3_16[7]}
   );
   gpc606_5 gpc1301 (
      {stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5], stage2_18[6]},
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage3_22[0],stage3_21[0],stage3_20[0],stage3_19[6],stage3_18[7]}
   );
   gpc606_5 gpc1302 (
      {stage2_18[7], stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11], stage2_18[12]},
      {stage2_20[6], stage2_20[7], stage2_20[8], stage2_20[9], stage2_20[10], stage2_20[11]},
      {stage3_22[1],stage3_21[1],stage3_20[1],stage3_19[7],stage3_18[8]}
   );
   gpc606_5 gpc1303 (
      {stage2_18[13], stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17], stage2_18[18]},
      {stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15], stage2_20[16], stage2_20[17]},
      {stage3_22[2],stage3_21[2],stage3_20[2],stage3_19[8],stage3_18[9]}
   );
   gpc615_5 gpc1304 (
      {stage2_18[19], stage2_18[20], stage2_18[21], stage2_18[22], stage2_18[23]},
      {stage2_19[0]},
      {stage2_20[18], stage2_20[19], stage2_20[20], stage2_20[21], stage2_20[22], stage2_20[23]},
      {stage3_22[3],stage3_21[3],stage3_20[3],stage3_19[9],stage3_18[10]}
   );
   gpc615_5 gpc1305 (
      {stage2_18[24], stage2_18[25], stage2_18[26], stage2_18[27], stage2_18[28]},
      {stage2_19[1]},
      {stage2_20[24], stage2_20[25], stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29]},
      {stage3_22[4],stage3_21[4],stage3_20[4],stage3_19[10],stage3_18[11]}
   );
   gpc615_5 gpc1306 (
      {stage2_18[29], stage2_18[30], stage2_18[31], stage2_18[32], stage2_18[33]},
      {stage2_19[2]},
      {stage2_20[30], stage2_20[31], stage2_20[32], stage2_20[33], stage2_20[34], stage2_20[35]},
      {stage3_22[5],stage3_21[5],stage3_20[5],stage3_19[11],stage3_18[12]}
   );
   gpc615_5 gpc1307 (
      {stage2_18[34], stage2_18[35], stage2_18[36], stage2_18[37], 1'b0},
      {stage2_19[3]},
      {stage2_20[36], stage2_20[37], stage2_20[38], stage2_20[39], stage2_20[40], stage2_20[41]},
      {stage3_22[6],stage3_21[6],stage3_20[6],stage3_19[12],stage3_18[13]}
   );
   gpc615_5 gpc1308 (
      {stage2_19[4], stage2_19[5], stage2_19[6], stage2_19[7], stage2_19[8]},
      {stage2_20[42]},
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5]},
      {stage3_23[0],stage3_22[7],stage3_21[7],stage3_20[7],stage3_19[13]}
   );
   gpc606_5 gpc1309 (
      {stage2_20[43], stage2_20[44], stage2_20[45], stage2_20[46], stage2_20[47], stage2_20[48]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[1],stage3_22[8],stage3_21[8],stage3_20[8]}
   );
   gpc606_5 gpc1310 (
      {stage2_21[6], stage2_21[7], stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage2_23[0], stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage3_25[0],stage3_24[1],stage3_23[2],stage3_22[9],stage3_21[9]}
   );
   gpc606_5 gpc1311 (
      {stage2_21[12], stage2_21[13], stage2_21[14], stage2_21[15], stage2_21[16], stage2_21[17]},
      {stage2_23[6], stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage3_25[1],stage3_24[2],stage3_23[3],stage3_22[10],stage3_21[10]}
   );
   gpc615_5 gpc1312 (
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10]},
      {stage2_23[12]},
      {stage2_24[0], stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage3_26[0],stage3_25[2],stage3_24[3],stage3_23[4],stage3_22[11]}
   );
   gpc615_5 gpc1313 (
      {stage2_22[11], stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15]},
      {stage2_23[13]},
      {stage2_24[6], stage2_24[7], stage2_24[8], stage2_24[9], stage2_24[10], stage2_24[11]},
      {stage3_26[1],stage3_25[3],stage3_24[4],stage3_23[5],stage3_22[12]}
   );
   gpc615_5 gpc1314 (
      {stage2_22[16], stage2_22[17], stage2_22[18], stage2_22[19], stage2_22[20]},
      {stage2_23[14]},
      {stage2_24[12], stage2_24[13], stage2_24[14], stage2_24[15], stage2_24[16], stage2_24[17]},
      {stage3_26[2],stage3_25[4],stage3_24[5],stage3_23[6],stage3_22[13]}
   );
   gpc615_5 gpc1315 (
      {stage2_22[21], stage2_22[22], stage2_22[23], stage2_22[24], stage2_22[25]},
      {stage2_23[15]},
      {stage2_24[18], stage2_24[19], stage2_24[20], stage2_24[21], stage2_24[22], stage2_24[23]},
      {stage3_26[3],stage3_25[5],stage3_24[6],stage3_23[7],stage3_22[14]}
   );
   gpc606_5 gpc1316 (
      {stage2_23[16], stage2_23[17], stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[4],stage3_25[6],stage3_24[7],stage3_23[8]}
   );
   gpc606_5 gpc1317 (
      {stage2_23[22], stage2_23[23], stage2_23[24], stage2_23[25], stage2_23[26], stage2_23[27]},
      {stage2_25[6], stage2_25[7], stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11]},
      {stage3_27[1],stage3_26[5],stage3_25[7],stage3_24[8],stage3_23[9]}
   );
   gpc606_5 gpc1318 (
      {stage2_23[28], stage2_23[29], stage2_23[30], stage2_23[31], stage2_23[32], stage2_23[33]},
      {stage2_25[12], stage2_25[13], stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17]},
      {stage3_27[2],stage3_26[6],stage3_25[8],stage3_24[9],stage3_23[10]}
   );
   gpc606_5 gpc1319 (
      {stage2_25[18], stage2_25[19], stage2_25[20], stage2_25[21], stage2_25[22], stage2_25[23]},
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4], stage2_27[5]},
      {stage3_29[0],stage3_28[0],stage3_27[3],stage3_26[7],stage3_25[9]}
   );
   gpc606_5 gpc1320 (
      {stage2_25[24], stage2_25[25], stage2_25[26], stage2_25[27], stage2_25[28], stage2_25[29]},
      {stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9], stage2_27[10], stage2_27[11]},
      {stage3_29[1],stage3_28[1],stage3_27[4],stage3_26[8],stage3_25[10]}
   );
   gpc606_5 gpc1321 (
      {stage2_25[30], stage2_25[31], stage2_25[32], stage2_25[33], stage2_25[34], stage2_25[35]},
      {stage2_27[12], stage2_27[13], stage2_27[14], stage2_27[15], stage2_27[16], stage2_27[17]},
      {stage3_29[2],stage3_28[2],stage3_27[5],stage3_26[9],stage3_25[11]}
   );
   gpc606_5 gpc1322 (
      {stage2_25[36], stage2_25[37], stage2_25[38], stage2_25[39], stage2_25[40], stage2_25[41]},
      {stage2_27[18], stage2_27[19], stage2_27[20], stage2_27[21], stage2_27[22], stage2_27[23]},
      {stage3_29[3],stage3_28[3],stage3_27[6],stage3_26[10],stage3_25[12]}
   );
   gpc615_5 gpc1323 (
      {stage2_25[42], stage2_25[43], stage2_25[44], stage2_25[45], stage2_25[46]},
      {stage2_26[0]},
      {stage2_27[24], stage2_27[25], stage2_27[26], stage2_27[27], stage2_27[28], stage2_27[29]},
      {stage3_29[4],stage3_28[4],stage3_27[7],stage3_26[11],stage3_25[13]}
   );
   gpc606_5 gpc1324 (
      {stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5], stage2_26[6]},
      {stage2_28[0], stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5]},
      {stage3_30[0],stage3_29[5],stage3_28[5],stage3_27[8],stage3_26[12]}
   );
   gpc606_5 gpc1325 (
      {stage2_26[7], stage2_26[8], stage2_26[9], stage2_26[10], stage2_26[11], stage2_26[12]},
      {stage2_28[6], stage2_28[7], stage2_28[8], stage2_28[9], stage2_28[10], stage2_28[11]},
      {stage3_30[1],stage3_29[6],stage3_28[6],stage3_27[9],stage3_26[13]}
   );
   gpc606_5 gpc1326 (
      {stage2_26[13], stage2_26[14], stage2_26[15], stage2_26[16], stage2_26[17], stage2_26[18]},
      {stage2_28[12], stage2_28[13], stage2_28[14], stage2_28[15], stage2_28[16], stage2_28[17]},
      {stage3_30[2],stage3_29[7],stage3_28[7],stage3_27[10],stage3_26[14]}
   );
   gpc606_5 gpc1327 (
      {stage2_26[19], stage2_26[20], stage2_26[21], stage2_26[22], stage2_26[23], stage2_26[24]},
      {stage2_28[18], stage2_28[19], stage2_28[20], stage2_28[21], stage2_28[22], stage2_28[23]},
      {stage3_30[3],stage3_29[8],stage3_28[8],stage3_27[11],stage3_26[15]}
   );
   gpc606_5 gpc1328 (
      {stage2_26[25], stage2_26[26], stage2_26[27], stage2_26[28], stage2_26[29], stage2_26[30]},
      {stage2_28[24], stage2_28[25], stage2_28[26], stage2_28[27], stage2_28[28], stage2_28[29]},
      {stage3_30[4],stage3_29[9],stage3_28[9],stage3_27[12],stage3_26[16]}
   );
   gpc615_5 gpc1329 (
      {stage2_26[31], stage2_26[32], stage2_26[33], stage2_26[34], stage2_26[35]},
      {stage2_27[30]},
      {stage2_28[30], stage2_28[31], stage2_28[32], stage2_28[33], stage2_28[34], stage2_28[35]},
      {stage3_30[5],stage3_29[10],stage3_28[10],stage3_27[13],stage3_26[17]}
   );
   gpc606_5 gpc1330 (
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage3_33[0],stage3_32[0],stage3_31[0],stage3_30[6],stage3_29[11]}
   );
   gpc606_5 gpc1331 (
      {stage2_29[6], stage2_29[7], stage2_29[8], stage2_29[9], stage2_29[10], stage2_29[11]},
      {stage2_31[6], stage2_31[7], stage2_31[8], stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage3_33[1],stage3_32[1],stage3_31[1],stage3_30[7],stage3_29[12]}
   );
   gpc606_5 gpc1332 (
      {stage2_29[12], stage2_29[13], stage2_29[14], stage2_29[15], stage2_29[16], stage2_29[17]},
      {stage2_31[12], stage2_31[13], stage2_31[14], stage2_31[15], stage2_31[16], stage2_31[17]},
      {stage3_33[2],stage3_32[2],stage3_31[2],stage3_30[8],stage3_29[13]}
   );
   gpc606_5 gpc1333 (
      {stage2_29[18], stage2_29[19], stage2_29[20], stage2_29[21], stage2_29[22], stage2_29[23]},
      {stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage3_33[3],stage3_32[3],stage3_31[3],stage3_30[9],stage3_29[14]}
   );
   gpc606_5 gpc1334 (
      {stage2_29[24], stage2_29[25], stage2_29[26], stage2_29[27], stage2_29[28], stage2_29[29]},
      {stage2_31[24], stage2_31[25], stage2_31[26], stage2_31[27], stage2_31[28], stage2_31[29]},
      {stage3_33[4],stage3_32[4],stage3_31[4],stage3_30[10],stage3_29[15]}
   );
   gpc606_5 gpc1335 (
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage2_32[0], stage2_32[1], stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5]},
      {stage3_34[0],stage3_33[5],stage3_32[5],stage3_31[5],stage3_30[11]}
   );
   gpc606_5 gpc1336 (
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10], stage2_32[11]},
      {stage3_34[1],stage3_33[6],stage3_32[6],stage3_31[6],stage3_30[12]}
   );
   gpc606_5 gpc1337 (
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16], stage2_32[17]},
      {stage3_34[2],stage3_33[7],stage3_32[7],stage3_31[7],stage3_30[13]}
   );
   gpc1415_5 gpc1338 (
      {stage2_31[30], stage2_31[31], stage2_31[32], stage2_31[33], 1'b0},
      {stage2_32[18]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3]},
      {stage2_34[0]},
      {stage3_35[0],stage3_34[3],stage3_33[8],stage3_32[8],stage3_31[8]}
   );
   gpc2135_5 gpc1339 (
      {stage2_32[19], stage2_32[20], stage2_32[21], stage2_32[22], stage2_32[23]},
      {stage2_33[4], stage2_33[5], stage2_33[6]},
      {stage2_34[1]},
      {stage2_35[0], stage2_35[1]},
      {stage3_36[0],stage3_35[1],stage3_34[4],stage3_33[9],stage3_32[9]}
   );
   gpc1_1 gpc1340 (
      {stage2_1[14]},
      {stage3_1[7]}
   );
   gpc1_1 gpc1341 (
      {stage2_1[15]},
      {stage3_1[8]}
   );
   gpc1_1 gpc1342 (
      {stage2_1[16]},
      {stage3_1[9]}
   );
   gpc1_1 gpc1343 (
      {stage2_1[17]},
      {stage3_1[10]}
   );
   gpc1_1 gpc1344 (
      {stage2_1[18]},
      {stage3_1[11]}
   );
   gpc1_1 gpc1345 (
      {stage2_1[19]},
      {stage3_1[12]}
   );
   gpc1_1 gpc1346 (
      {stage2_4[23]},
      {stage3_4[15]}
   );
   gpc1_1 gpc1347 (
      {stage2_4[24]},
      {stage3_4[16]}
   );
   gpc1_1 gpc1348 (
      {stage2_4[25]},
      {stage3_4[17]}
   );
   gpc1_1 gpc1349 (
      {stage2_5[30]},
      {stage3_5[8]}
   );
   gpc1_1 gpc1350 (
      {stage2_6[24]},
      {stage3_6[10]}
   );
   gpc1_1 gpc1351 (
      {stage2_6[25]},
      {stage3_6[11]}
   );
   gpc1_1 gpc1352 (
      {stage2_6[26]},
      {stage3_6[12]}
   );
   gpc1_1 gpc1353 (
      {stage2_6[27]},
      {stage3_6[13]}
   );
   gpc1_1 gpc1354 (
      {stage2_6[28]},
      {stage3_6[14]}
   );
   gpc1_1 gpc1355 (
      {stage2_6[29]},
      {stage3_6[15]}
   );
   gpc1_1 gpc1356 (
      {stage2_6[30]},
      {stage3_6[16]}
   );
   gpc1_1 gpc1357 (
      {stage2_6[31]},
      {stage3_6[17]}
   );
   gpc1_1 gpc1358 (
      {stage2_6[32]},
      {stage3_6[18]}
   );
   gpc1_1 gpc1359 (
      {stage2_6[33]},
      {stage3_6[19]}
   );
   gpc1_1 gpc1360 (
      {stage2_6[34]},
      {stage3_6[20]}
   );
   gpc1_1 gpc1361 (
      {stage2_6[35]},
      {stage3_6[21]}
   );
   gpc1_1 gpc1362 (
      {stage2_6[36]},
      {stage3_6[22]}
   );
   gpc1_1 gpc1363 (
      {stage2_6[37]},
      {stage3_6[23]}
   );
   gpc1_1 gpc1364 (
      {stage2_6[38]},
      {stage3_6[24]}
   );
   gpc1_1 gpc1365 (
      {stage2_6[39]},
      {stage3_6[25]}
   );
   gpc1_1 gpc1366 (
      {stage2_6[40]},
      {stage3_6[26]}
   );
   gpc1_1 gpc1367 (
      {stage2_6[41]},
      {stage3_6[27]}
   );
   gpc1_1 gpc1368 (
      {stage2_6[42]},
      {stage3_6[28]}
   );
   gpc1_1 gpc1369 (
      {stage2_6[43]},
      {stage3_6[29]}
   );
   gpc1_1 gpc1370 (
      {stage2_6[44]},
      {stage3_6[30]}
   );
   gpc1_1 gpc1371 (
      {stage2_6[45]},
      {stage3_6[31]}
   );
   gpc1_1 gpc1372 (
      {stage2_6[46]},
      {stage3_6[32]}
   );
   gpc1_1 gpc1373 (
      {stage2_6[47]},
      {stage3_6[33]}
   );
   gpc1_1 gpc1374 (
      {stage2_8[33]},
      {stage3_8[11]}
   );
   gpc1_1 gpc1375 (
      {stage2_8[34]},
      {stage3_8[12]}
   );
   gpc1_1 gpc1376 (
      {stage2_8[35]},
      {stage3_8[13]}
   );
   gpc1_1 gpc1377 (
      {stage2_8[36]},
      {stage3_8[14]}
   );
   gpc1_1 gpc1378 (
      {stage2_8[37]},
      {stage3_8[15]}
   );
   gpc1_1 gpc1379 (
      {stage2_8[38]},
      {stage3_8[16]}
   );
   gpc1_1 gpc1380 (
      {stage2_10[18]},
      {stage3_10[9]}
   );
   gpc1_1 gpc1381 (
      {stage2_10[19]},
      {stage3_10[10]}
   );
   gpc1_1 gpc1382 (
      {stage2_10[20]},
      {stage3_10[11]}
   );
   gpc1_1 gpc1383 (
      {stage2_10[21]},
      {stage3_10[12]}
   );
   gpc1_1 gpc1384 (
      {stage2_11[25]},
      {stage3_11[12]}
   );
   gpc1_1 gpc1385 (
      {stage2_11[26]},
      {stage3_11[13]}
   );
   gpc1_1 gpc1386 (
      {stage2_12[11]},
      {stage3_12[9]}
   );
   gpc1_1 gpc1387 (
      {stage2_12[12]},
      {stage3_12[10]}
   );
   gpc1_1 gpc1388 (
      {stage2_12[13]},
      {stage3_12[11]}
   );
   gpc1_1 gpc1389 (
      {stage2_12[14]},
      {stage3_12[12]}
   );
   gpc1_1 gpc1390 (
      {stage2_12[15]},
      {stage3_12[13]}
   );
   gpc1_1 gpc1391 (
      {stage2_12[16]},
      {stage3_12[14]}
   );
   gpc1_1 gpc1392 (
      {stage2_12[17]},
      {stage3_12[15]}
   );
   gpc1_1 gpc1393 (
      {stage2_12[18]},
      {stage3_12[16]}
   );
   gpc1_1 gpc1394 (
      {stage2_12[19]},
      {stage3_12[17]}
   );
   gpc1_1 gpc1395 (
      {stage2_12[20]},
      {stage3_12[18]}
   );
   gpc1_1 gpc1396 (
      {stage2_13[30]},
      {stage3_13[6]}
   );
   gpc1_1 gpc1397 (
      {stage2_13[31]},
      {stage3_13[7]}
   );
   gpc1_1 gpc1398 (
      {stage2_13[32]},
      {stage3_13[8]}
   );
   gpc1_1 gpc1399 (
      {stage2_13[33]},
      {stage3_13[9]}
   );
   gpc1_1 gpc1400 (
      {stage2_13[34]},
      {stage3_13[10]}
   );
   gpc1_1 gpc1401 (
      {stage2_14[12]},
      {stage3_14[7]}
   );
   gpc1_1 gpc1402 (
      {stage2_14[13]},
      {stage3_14[8]}
   );
   gpc1_1 gpc1403 (
      {stage2_14[14]},
      {stage3_14[9]}
   );
   gpc1_1 gpc1404 (
      {stage2_14[15]},
      {stage3_14[10]}
   );
   gpc1_1 gpc1405 (
      {stage2_14[16]},
      {stage3_14[11]}
   );
   gpc1_1 gpc1406 (
      {stage2_14[17]},
      {stage3_14[12]}
   );
   gpc1_1 gpc1407 (
      {stage2_14[18]},
      {stage3_14[13]}
   );
   gpc1_1 gpc1408 (
      {stage2_14[19]},
      {stage3_14[14]}
   );
   gpc1_1 gpc1409 (
      {stage2_14[20]},
      {stage3_14[15]}
   );
   gpc1_1 gpc1410 (
      {stage2_14[21]},
      {stage3_14[16]}
   );
   gpc1_1 gpc1411 (
      {stage2_14[22]},
      {stage3_14[17]}
   );
   gpc1_1 gpc1412 (
      {stage2_14[23]},
      {stage3_14[18]}
   );
   gpc1_1 gpc1413 (
      {stage2_14[24]},
      {stage3_14[19]}
   );
   gpc1_1 gpc1414 (
      {stage2_14[25]},
      {stage3_14[20]}
   );
   gpc1_1 gpc1415 (
      {stage2_14[26]},
      {stage3_14[21]}
   );
   gpc1_1 gpc1416 (
      {stage2_16[18]},
      {stage3_16[8]}
   );
   gpc1_1 gpc1417 (
      {stage2_16[19]},
      {stage3_16[9]}
   );
   gpc1_1 gpc1418 (
      {stage2_16[20]},
      {stage3_16[10]}
   );
   gpc1_1 gpc1419 (
      {stage2_16[21]},
      {stage3_16[11]}
   );
   gpc1_1 gpc1420 (
      {stage2_16[22]},
      {stage3_16[12]}
   );
   gpc1_1 gpc1421 (
      {stage2_17[31]},
      {stage3_17[7]}
   );
   gpc1_1 gpc1422 (
      {stage2_17[32]},
      {stage3_17[8]}
   );
   gpc1_1 gpc1423 (
      {stage2_17[33]},
      {stage3_17[9]}
   );
   gpc1_1 gpc1424 (
      {stage2_17[34]},
      {stage3_17[10]}
   );
   gpc1_1 gpc1425 (
      {stage2_17[35]},
      {stage3_17[11]}
   );
   gpc1_1 gpc1426 (
      {stage2_17[36]},
      {stage3_17[12]}
   );
   gpc1_1 gpc1427 (
      {stage2_17[37]},
      {stage3_17[13]}
   );
   gpc1_1 gpc1428 (
      {stage2_17[38]},
      {stage3_17[14]}
   );
   gpc1_1 gpc1429 (
      {stage2_17[39]},
      {stage3_17[15]}
   );
   gpc1_1 gpc1430 (
      {stage2_17[40]},
      {stage3_17[16]}
   );
   gpc1_1 gpc1431 (
      {stage2_17[41]},
      {stage3_17[17]}
   );
   gpc1_1 gpc1432 (
      {stage2_17[42]},
      {stage3_17[18]}
   );
   gpc1_1 gpc1433 (
      {stage2_17[43]},
      {stage3_17[19]}
   );
   gpc1_1 gpc1434 (
      {stage2_17[44]},
      {stage3_17[20]}
   );
   gpc1_1 gpc1435 (
      {stage2_17[45]},
      {stage3_17[21]}
   );
   gpc1_1 gpc1436 (
      {stage2_17[46]},
      {stage3_17[22]}
   );
   gpc1_1 gpc1437 (
      {stage2_17[47]},
      {stage3_17[23]}
   );
   gpc1_1 gpc1438 (
      {stage2_17[48]},
      {stage3_17[24]}
   );
   gpc1_1 gpc1439 (
      {stage2_19[9]},
      {stage3_19[14]}
   );
   gpc1_1 gpc1440 (
      {stage2_19[10]},
      {stage3_19[15]}
   );
   gpc1_1 gpc1441 (
      {stage2_19[11]},
      {stage3_19[16]}
   );
   gpc1_1 gpc1442 (
      {stage2_19[12]},
      {stage3_19[17]}
   );
   gpc1_1 gpc1443 (
      {stage2_19[13]},
      {stage3_19[18]}
   );
   gpc1_1 gpc1444 (
      {stage2_19[14]},
      {stage3_19[19]}
   );
   gpc1_1 gpc1445 (
      {stage2_19[15]},
      {stage3_19[20]}
   );
   gpc1_1 gpc1446 (
      {stage2_19[16]},
      {stage3_19[21]}
   );
   gpc1_1 gpc1447 (
      {stage2_19[17]},
      {stage3_19[22]}
   );
   gpc1_1 gpc1448 (
      {stage2_19[18]},
      {stage3_19[23]}
   );
   gpc1_1 gpc1449 (
      {stage2_19[19]},
      {stage3_19[24]}
   );
   gpc1_1 gpc1450 (
      {stage2_19[20]},
      {stage3_19[25]}
   );
   gpc1_1 gpc1451 (
      {stage2_20[49]},
      {stage3_20[9]}
   );
   gpc1_1 gpc1452 (
      {stage2_20[50]},
      {stage3_20[10]}
   );
   gpc1_1 gpc1453 (
      {stage2_20[51]},
      {stage3_20[11]}
   );
   gpc1_1 gpc1454 (
      {stage2_20[52]},
      {stage3_20[12]}
   );
   gpc1_1 gpc1455 (
      {stage2_20[53]},
      {stage3_20[13]}
   );
   gpc1_1 gpc1456 (
      {stage2_20[54]},
      {stage3_20[14]}
   );
   gpc1_1 gpc1457 (
      {stage2_20[55]},
      {stage3_20[15]}
   );
   gpc1_1 gpc1458 (
      {stage2_21[18]},
      {stage3_21[11]}
   );
   gpc1_1 gpc1459 (
      {stage2_21[19]},
      {stage3_21[12]}
   );
   gpc1_1 gpc1460 (
      {stage2_21[20]},
      {stage3_21[13]}
   );
   gpc1_1 gpc1461 (
      {stage2_22[26]},
      {stage3_22[15]}
   );
   gpc1_1 gpc1462 (
      {stage2_24[24]},
      {stage3_24[10]}
   );
   gpc1_1 gpc1463 (
      {stage2_24[25]},
      {stage3_24[11]}
   );
   gpc1_1 gpc1464 (
      {stage2_24[26]},
      {stage3_24[12]}
   );
   gpc1_1 gpc1465 (
      {stage2_24[27]},
      {stage3_24[13]}
   );
   gpc1_1 gpc1466 (
      {stage2_24[28]},
      {stage3_24[14]}
   );
   gpc1_1 gpc1467 (
      {stage2_24[29]},
      {stage3_24[15]}
   );
   gpc1_1 gpc1468 (
      {stage2_24[30]},
      {stage3_24[16]}
   );
   gpc1_1 gpc1469 (
      {stage2_24[31]},
      {stage3_24[17]}
   );
   gpc1_1 gpc1470 (
      {stage2_24[32]},
      {stage3_24[18]}
   );
   gpc1_1 gpc1471 (
      {stage2_26[36]},
      {stage3_26[18]}
   );
   gpc1_1 gpc1472 (
      {stage2_29[30]},
      {stage3_29[16]}
   );
   gpc1_1 gpc1473 (
      {stage2_29[31]},
      {stage3_29[17]}
   );
   gpc1_1 gpc1474 (
      {stage2_30[18]},
      {stage3_30[14]}
   );
   gpc1_1 gpc1475 (
      {stage2_32[24]},
      {stage3_32[10]}
   );
   gpc1_1 gpc1476 (
      {stage2_32[25]},
      {stage3_32[11]}
   );
   gpc1_1 gpc1477 (
      {stage2_32[26]},
      {stage3_32[12]}
   );
   gpc1_1 gpc1478 (
      {stage2_32[27]},
      {stage3_32[13]}
   );
   gpc1_1 gpc1479 (
      {stage2_32[28]},
      {stage3_32[14]}
   );
   gpc1_1 gpc1480 (
      {stage2_33[7]},
      {stage3_33[10]}
   );
   gpc1_1 gpc1481 (
      {stage2_33[8]},
      {stage3_33[11]}
   );
   gpc1_1 gpc1482 (
      {stage2_33[9]},
      {stage3_33[12]}
   );
   gpc1_1 gpc1483 (
      {stage2_33[10]},
      {stage3_33[13]}
   );
   gpc1_1 gpc1484 (
      {stage2_33[11]},
      {stage3_33[14]}
   );
   gpc1_1 gpc1485 (
      {stage2_33[12]},
      {stage3_33[15]}
   );
   gpc1_1 gpc1486 (
      {stage2_33[13]},
      {stage3_33[16]}
   );
   gpc1_1 gpc1487 (
      {stage2_33[14]},
      {stage3_33[17]}
   );
   gpc1_1 gpc1488 (
      {stage2_33[15]},
      {stage3_33[18]}
   );
   gpc1_1 gpc1489 (
      {stage2_33[16]},
      {stage3_33[19]}
   );
   gpc1_1 gpc1490 (
      {stage2_33[17]},
      {stage3_33[20]}
   );
   gpc1_1 gpc1491 (
      {stage2_34[2]},
      {stage3_34[5]}
   );
   gpc1_1 gpc1492 (
      {stage2_34[3]},
      {stage3_34[6]}
   );
   gpc1_1 gpc1493 (
      {stage2_34[4]},
      {stage3_34[7]}
   );
   gpc1_1 gpc1494 (
      {stage2_34[5]},
      {stage3_34[8]}
   );
   gpc606_5 gpc1495 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4], stage3_0[5]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc207_4 gpc1496 (
      {stage3_1[0], stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5], stage3_1[6]},
      {stage3_3[0], stage3_3[1]},
      {stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc117_4 gpc1497 (
      {stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5], stage3_3[6], stage3_3[7], stage3_3[8]},
      {stage3_4[0]},
      {stage3_5[0]},
      {stage4_6[0],stage4_5[0],stage4_4[2],stage4_3[2]}
   );
   gpc615_5 gpc1498 (
      {stage3_4[1], stage3_4[2], stage3_4[3], stage3_4[4], stage3_4[5]},
      {stage3_5[1]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[1],stage4_4[3]}
   );
   gpc615_5 gpc1499 (
      {stage3_4[6], stage3_4[7], stage3_4[8], stage3_4[9], stage3_4[10]},
      {stage3_5[2]},
      {stage3_6[6], stage3_6[7], stage3_6[8], stage3_6[9], stage3_6[10], stage3_6[11]},
      {stage4_8[1],stage4_7[1],stage4_6[2],stage4_5[2],stage4_4[4]}
   );
   gpc615_5 gpc1500 (
      {stage3_4[11], stage3_4[12], stage3_4[13], stage3_4[14], stage3_4[15]},
      {stage3_5[3]},
      {stage3_6[12], stage3_6[13], stage3_6[14], stage3_6[15], stage3_6[16], stage3_6[17]},
      {stage4_8[2],stage4_7[2],stage4_6[3],stage4_5[3],stage4_4[5]}
   );
   gpc1343_5 gpc1501 (
      {stage3_6[18], stage3_6[19], stage3_6[20]},
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3]},
      {stage3_8[0], stage3_8[1], stage3_8[2]},
      {stage3_9[0]},
      {stage4_10[0],stage4_9[0],stage4_8[3],stage4_7[3],stage4_6[4]}
   );
   gpc1343_5 gpc1502 (
      {stage3_6[21], stage3_6[22], stage3_6[23]},
      {stage3_7[4], stage3_7[5], stage3_7[6], stage3_7[7]},
      {stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage3_9[1]},
      {stage4_10[1],stage4_9[1],stage4_8[4],stage4_7[4],stage4_6[5]}
   );
   gpc606_5 gpc1503 (
      {stage3_6[24], stage3_6[25], stage3_6[26], stage3_6[27], stage3_6[28], stage3_6[29]},
      {stage3_8[6], stage3_8[7], stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11]},
      {stage4_10[2],stage4_9[2],stage4_8[5],stage4_7[5],stage4_6[6]}
   );
   gpc1343_5 gpc1504 (
      {stage3_9[2], stage3_9[3], stage3_9[4]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3]},
      {stage3_11[0], stage3_11[1], stage3_11[2]},
      {stage3_12[0]},
      {stage4_13[0],stage4_12[0],stage4_11[0],stage4_10[3],stage4_9[3]}
   );
   gpc1343_5 gpc1505 (
      {stage3_9[5], stage3_9[6], stage3_9[7]},
      {stage3_10[4], stage3_10[5], stage3_10[6], stage3_10[7]},
      {stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage3_12[1]},
      {stage4_13[1],stage4_12[1],stage4_11[1],stage4_10[4],stage4_9[4]}
   );
   gpc1343_5 gpc1506 (
      {stage3_9[8], 1'b0, 1'b0},
      {stage3_10[8], stage3_10[9], stage3_10[10], stage3_10[11]},
      {stage3_11[6], stage3_11[7], stage3_11[8]},
      {stage3_12[2]},
      {stage4_13[2],stage4_12[2],stage4_11[2],stage4_10[5],stage4_9[5]}
   );
   gpc615_5 gpc1507 (
      {stage3_11[9], stage3_11[10], stage3_11[11], stage3_11[12], stage3_11[13]},
      {stage3_12[3]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[0],stage4_13[3],stage4_12[3],stage4_11[3]}
   );
   gpc606_5 gpc1508 (
      {stage3_12[4], stage3_12[5], stage3_12[6], stage3_12[7], stage3_12[8], stage3_12[9]},
      {stage3_14[0], stage3_14[1], stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5]},
      {stage4_16[0],stage4_15[1],stage4_14[1],stage4_13[4],stage4_12[4]}
   );
   gpc606_5 gpc1509 (
      {stage3_12[10], stage3_12[11], stage3_12[12], stage3_12[13], stage3_12[14], stage3_12[15]},
      {stage3_14[6], stage3_14[7], stage3_14[8], stage3_14[9], stage3_14[10], stage3_14[11]},
      {stage4_16[1],stage4_15[2],stage4_14[2],stage4_13[5],stage4_12[5]}
   );
   gpc207_4 gpc1510 (
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], 1'b0, 1'b0},
      {stage3_15[0], stage3_15[1]},
      {stage4_16[2],stage4_15[3],stage4_14[3],stage4_13[6]}
   );
   gpc615_5 gpc1511 (
      {stage3_14[12], stage3_14[13], stage3_14[14], stage3_14[15], stage3_14[16]},
      {stage3_15[2]},
      {stage3_16[0], stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5]},
      {stage4_18[0],stage4_17[0],stage4_16[3],stage4_15[4],stage4_14[4]}
   );
   gpc615_5 gpc1512 (
      {stage3_14[17], stage3_14[18], stage3_14[19], stage3_14[20], stage3_14[21]},
      {stage3_15[3]},
      {stage3_16[6], stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11]},
      {stage4_18[1],stage4_17[1],stage4_16[4],stage4_15[5],stage4_14[5]}
   );
   gpc606_5 gpc1513 (
      {stage3_15[4], stage3_15[5], stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9]},
      {stage3_17[0], stage3_17[1], stage3_17[2], stage3_17[3], stage3_17[4], stage3_17[5]},
      {stage4_19[0],stage4_18[2],stage4_17[2],stage4_16[5],stage4_15[6]}
   );
   gpc606_5 gpc1514 (
      {stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9], stage3_17[10], stage3_17[11]},
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4], stage3_19[5]},
      {stage4_21[0],stage4_20[0],stage4_19[1],stage4_18[3],stage4_17[3]}
   );
   gpc606_5 gpc1515 (
      {stage3_17[12], stage3_17[13], stage3_17[14], stage3_17[15], stage3_17[16], stage3_17[17]},
      {stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9], stage3_19[10], stage3_19[11]},
      {stage4_21[1],stage4_20[1],stage4_19[2],stage4_18[4],stage4_17[4]}
   );
   gpc606_5 gpc1516 (
      {stage3_17[18], stage3_17[19], stage3_17[20], stage3_17[21], stage3_17[22], stage3_17[23]},
      {stage3_19[12], stage3_19[13], stage3_19[14], stage3_19[15], stage3_19[16], stage3_19[17]},
      {stage4_21[2],stage4_20[2],stage4_19[3],stage4_18[5],stage4_17[5]}
   );
   gpc615_5 gpc1517 (
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4]},
      {stage3_19[18]},
      {stage3_20[0], stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4], stage3_20[5]},
      {stage4_22[0],stage4_21[3],stage4_20[3],stage4_19[4],stage4_18[6]}
   );
   gpc615_5 gpc1518 (
      {stage3_18[5], stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9]},
      {stage3_19[19]},
      {stage3_20[6], stage3_20[7], stage3_20[8], stage3_20[9], stage3_20[10], stage3_20[11]},
      {stage4_22[1],stage4_21[4],stage4_20[4],stage4_19[5],stage4_18[7]}
   );
   gpc615_5 gpc1519 (
      {stage3_19[20], stage3_19[21], stage3_19[22], stage3_19[23], stage3_19[24]},
      {stage3_20[12]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[2],stage4_21[5],stage4_20[5],stage4_19[6]}
   );
   gpc606_5 gpc1520 (
      {stage3_20[13], stage3_20[14], stage3_20[15], 1'b0, 1'b0, 1'b0},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[1],stage4_22[3],stage4_21[6],stage4_20[6]}
   );
   gpc606_5 gpc1521 (
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage4_25[0],stage4_24[1],stage4_23[2],stage4_22[4],stage4_21[7]}
   );
   gpc615_5 gpc1522 (
      {stage3_22[6], stage3_22[7], stage3_22[8], stage3_22[9], stage3_22[10]},
      {stage3_23[6]},
      {stage3_24[0], stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5]},
      {stage4_26[0],stage4_25[1],stage4_24[2],stage4_23[3],stage4_22[5]}
   );
   gpc615_5 gpc1523 (
      {stage3_22[11], stage3_22[12], stage3_22[13], stage3_22[14], stage3_22[15]},
      {stage3_23[7]},
      {stage3_24[6], stage3_24[7], stage3_24[8], stage3_24[9], stage3_24[10], stage3_24[11]},
      {stage4_26[1],stage4_25[2],stage4_24[3],stage4_23[4],stage4_22[6]}
   );
   gpc615_5 gpc1524 (
      {stage3_25[0], stage3_25[1], stage3_25[2], stage3_25[3], stage3_25[4]},
      {stage3_26[0]},
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5]},
      {stage4_29[0],stage4_28[0],stage4_27[0],stage4_26[2],stage4_25[3]}
   );
   gpc1325_5 gpc1525 (
      {stage3_25[5], stage3_25[6], stage3_25[7], stage3_25[8], stage3_25[9]},
      {stage3_26[1], stage3_26[2]},
      {stage3_27[6], stage3_27[7], stage3_27[8]},
      {stage3_28[0]},
      {stage4_29[1],stage4_28[1],stage4_27[1],stage4_26[3],stage4_25[4]}
   );
   gpc1325_5 gpc1526 (
      {stage3_25[10], stage3_25[11], stage3_25[12], stage3_25[13], 1'b0},
      {stage3_26[3], stage3_26[4]},
      {stage3_27[9], stage3_27[10], stage3_27[11]},
      {stage3_28[1]},
      {stage4_29[2],stage4_28[2],stage4_27[2],stage4_26[4],stage4_25[5]}
   );
   gpc7_3 gpc1527 (
      {stage3_26[5], stage3_26[6], stage3_26[7], stage3_26[8], stage3_26[9], stage3_26[10], stage3_26[11]},
      {stage4_28[3],stage4_27[3],stage4_26[5]}
   );
   gpc1163_5 gpc1528 (
      {stage3_28[2], stage3_28[3], stage3_28[4]},
      {stage3_29[0], stage3_29[1], stage3_29[2], stage3_29[3], stage3_29[4], stage3_29[5]},
      {stage3_30[0]},
      {stage3_31[0]},
      {stage4_32[0],stage4_31[0],stage4_30[0],stage4_29[3],stage4_28[4]}
   );
   gpc1163_5 gpc1529 (
      {stage3_28[5], stage3_28[6], stage3_28[7]},
      {stage3_29[6], stage3_29[7], stage3_29[8], stage3_29[9], stage3_29[10], stage3_29[11]},
      {stage3_30[1]},
      {stage3_31[1]},
      {stage4_32[1],stage4_31[1],stage4_30[1],stage4_29[4],stage4_28[5]}
   );
   gpc1163_5 gpc1530 (
      {stage3_28[8], stage3_28[9], stage3_28[10]},
      {stage3_29[12], stage3_29[13], stage3_29[14], stage3_29[15], stage3_29[16], stage3_29[17]},
      {stage3_30[2]},
      {stage3_31[2]},
      {stage4_32[2],stage4_31[2],stage4_30[2],stage4_29[5],stage4_28[6]}
   );
   gpc606_5 gpc1531 (
      {stage3_30[3], stage3_30[4], stage3_30[5], stage3_30[6], stage3_30[7], stage3_30[8]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5]},
      {stage4_34[0],stage4_33[0],stage4_32[3],stage4_31[3],stage4_30[3]}
   );
   gpc606_5 gpc1532 (
      {stage3_30[9], stage3_30[10], stage3_30[11], stage3_30[12], stage3_30[13], stage3_30[14]},
      {stage3_32[6], stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage4_34[1],stage4_33[1],stage4_32[4],stage4_31[4],stage4_30[4]}
   );
   gpc606_5 gpc1533 (
      {stage3_31[3], stage3_31[4], stage3_31[5], stage3_31[6], stage3_31[7], stage3_31[8]},
      {stage3_33[0], stage3_33[1], stage3_33[2], stage3_33[3], stage3_33[4], stage3_33[5]},
      {stage4_35[0],stage4_34[2],stage4_33[2],stage4_32[5],stage4_31[5]}
   );
   gpc1163_5 gpc1534 (
      {stage3_32[12], stage3_32[13], stage3_32[14]},
      {stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9], stage3_33[10], stage3_33[11]},
      {stage3_34[0]},
      {stage3_35[0]},
      {stage4_36[0],stage4_35[1],stage4_34[3],stage4_33[3],stage4_32[6]}
   );
   gpc1_1 gpc1535 (
      {stage3_0[6]},
      {stage4_0[1]}
   );
   gpc1_1 gpc1536 (
      {stage3_1[7]},
      {stage4_1[2]}
   );
   gpc1_1 gpc1537 (
      {stage3_1[8]},
      {stage4_1[3]}
   );
   gpc1_1 gpc1538 (
      {stage3_1[9]},
      {stage4_1[4]}
   );
   gpc1_1 gpc1539 (
      {stage3_1[10]},
      {stage4_1[5]}
   );
   gpc1_1 gpc1540 (
      {stage3_1[11]},
      {stage4_1[6]}
   );
   gpc1_1 gpc1541 (
      {stage3_1[12]},
      {stage4_1[7]}
   );
   gpc1_1 gpc1542 (
      {stage3_2[6]},
      {stage4_2[2]}
   );
   gpc1_1 gpc1543 (
      {stage3_2[7]},
      {stage4_2[3]}
   );
   gpc1_1 gpc1544 (
      {stage3_3[9]},
      {stage4_3[3]}
   );
   gpc1_1 gpc1545 (
      {stage3_3[10]},
      {stage4_3[4]}
   );
   gpc1_1 gpc1546 (
      {stage3_3[11]},
      {stage4_3[5]}
   );
   gpc1_1 gpc1547 (
      {stage3_3[12]},
      {stage4_3[6]}
   );
   gpc1_1 gpc1548 (
      {stage3_4[16]},
      {stage4_4[6]}
   );
   gpc1_1 gpc1549 (
      {stage3_4[17]},
      {stage4_4[7]}
   );
   gpc1_1 gpc1550 (
      {stage3_5[4]},
      {stage4_5[4]}
   );
   gpc1_1 gpc1551 (
      {stage3_5[5]},
      {stage4_5[5]}
   );
   gpc1_1 gpc1552 (
      {stage3_5[6]},
      {stage4_5[6]}
   );
   gpc1_1 gpc1553 (
      {stage3_5[7]},
      {stage4_5[7]}
   );
   gpc1_1 gpc1554 (
      {stage3_5[8]},
      {stage4_5[8]}
   );
   gpc1_1 gpc1555 (
      {stage3_6[30]},
      {stage4_6[7]}
   );
   gpc1_1 gpc1556 (
      {stage3_6[31]},
      {stage4_6[8]}
   );
   gpc1_1 gpc1557 (
      {stage3_6[32]},
      {stage4_6[9]}
   );
   gpc1_1 gpc1558 (
      {stage3_6[33]},
      {stage4_6[10]}
   );
   gpc1_1 gpc1559 (
      {stage3_7[8]},
      {stage4_7[6]}
   );
   gpc1_1 gpc1560 (
      {stage3_7[9]},
      {stage4_7[7]}
   );
   gpc1_1 gpc1561 (
      {stage3_7[10]},
      {stage4_7[8]}
   );
   gpc1_1 gpc1562 (
      {stage3_7[11]},
      {stage4_7[9]}
   );
   gpc1_1 gpc1563 (
      {stage3_7[12]},
      {stage4_7[10]}
   );
   gpc1_1 gpc1564 (
      {stage3_8[12]},
      {stage4_8[6]}
   );
   gpc1_1 gpc1565 (
      {stage3_8[13]},
      {stage4_8[7]}
   );
   gpc1_1 gpc1566 (
      {stage3_8[14]},
      {stage4_8[8]}
   );
   gpc1_1 gpc1567 (
      {stage3_8[15]},
      {stage4_8[9]}
   );
   gpc1_1 gpc1568 (
      {stage3_8[16]},
      {stage4_8[10]}
   );
   gpc1_1 gpc1569 (
      {stage3_10[12]},
      {stage4_10[6]}
   );
   gpc1_1 gpc1570 (
      {stage3_12[16]},
      {stage4_12[6]}
   );
   gpc1_1 gpc1571 (
      {stage3_12[17]},
      {stage4_12[7]}
   );
   gpc1_1 gpc1572 (
      {stage3_12[18]},
      {stage4_12[8]}
   );
   gpc1_1 gpc1573 (
      {stage3_15[10]},
      {stage4_15[7]}
   );
   gpc1_1 gpc1574 (
      {stage3_15[11]},
      {stage4_15[8]}
   );
   gpc1_1 gpc1575 (
      {stage3_16[12]},
      {stage4_16[6]}
   );
   gpc1_1 gpc1576 (
      {stage3_17[24]},
      {stage4_17[6]}
   );
   gpc1_1 gpc1577 (
      {stage3_18[10]},
      {stage4_18[8]}
   );
   gpc1_1 gpc1578 (
      {stage3_18[11]},
      {stage4_18[9]}
   );
   gpc1_1 gpc1579 (
      {stage3_18[12]},
      {stage4_18[10]}
   );
   gpc1_1 gpc1580 (
      {stage3_18[13]},
      {stage4_18[11]}
   );
   gpc1_1 gpc1581 (
      {stage3_19[25]},
      {stage4_19[7]}
   );
   gpc1_1 gpc1582 (
      {stage3_21[12]},
      {stage4_21[8]}
   );
   gpc1_1 gpc1583 (
      {stage3_21[13]},
      {stage4_21[9]}
   );
   gpc1_1 gpc1584 (
      {stage3_23[8]},
      {stage4_23[5]}
   );
   gpc1_1 gpc1585 (
      {stage3_23[9]},
      {stage4_23[6]}
   );
   gpc1_1 gpc1586 (
      {stage3_23[10]},
      {stage4_23[7]}
   );
   gpc1_1 gpc1587 (
      {stage3_24[12]},
      {stage4_24[4]}
   );
   gpc1_1 gpc1588 (
      {stage3_24[13]},
      {stage4_24[5]}
   );
   gpc1_1 gpc1589 (
      {stage3_24[14]},
      {stage4_24[6]}
   );
   gpc1_1 gpc1590 (
      {stage3_24[15]},
      {stage4_24[7]}
   );
   gpc1_1 gpc1591 (
      {stage3_24[16]},
      {stage4_24[8]}
   );
   gpc1_1 gpc1592 (
      {stage3_24[17]},
      {stage4_24[9]}
   );
   gpc1_1 gpc1593 (
      {stage3_24[18]},
      {stage4_24[10]}
   );
   gpc1_1 gpc1594 (
      {stage3_26[12]},
      {stage4_26[6]}
   );
   gpc1_1 gpc1595 (
      {stage3_26[13]},
      {stage4_26[7]}
   );
   gpc1_1 gpc1596 (
      {stage3_26[14]},
      {stage4_26[8]}
   );
   gpc1_1 gpc1597 (
      {stage3_26[15]},
      {stage4_26[9]}
   );
   gpc1_1 gpc1598 (
      {stage3_26[16]},
      {stage4_26[10]}
   );
   gpc1_1 gpc1599 (
      {stage3_26[17]},
      {stage4_26[11]}
   );
   gpc1_1 gpc1600 (
      {stage3_26[18]},
      {stage4_26[12]}
   );
   gpc1_1 gpc1601 (
      {stage3_27[12]},
      {stage4_27[4]}
   );
   gpc1_1 gpc1602 (
      {stage3_27[13]},
      {stage4_27[5]}
   );
   gpc1_1 gpc1603 (
      {stage3_33[12]},
      {stage4_33[4]}
   );
   gpc1_1 gpc1604 (
      {stage3_33[13]},
      {stage4_33[5]}
   );
   gpc1_1 gpc1605 (
      {stage3_33[14]},
      {stage4_33[6]}
   );
   gpc1_1 gpc1606 (
      {stage3_33[15]},
      {stage4_33[7]}
   );
   gpc1_1 gpc1607 (
      {stage3_33[16]},
      {stage4_33[8]}
   );
   gpc1_1 gpc1608 (
      {stage3_33[17]},
      {stage4_33[9]}
   );
   gpc1_1 gpc1609 (
      {stage3_33[18]},
      {stage4_33[10]}
   );
   gpc1_1 gpc1610 (
      {stage3_33[19]},
      {stage4_33[11]}
   );
   gpc1_1 gpc1611 (
      {stage3_33[20]},
      {stage4_33[12]}
   );
   gpc1_1 gpc1612 (
      {stage3_34[1]},
      {stage4_34[4]}
   );
   gpc1_1 gpc1613 (
      {stage3_34[2]},
      {stage4_34[5]}
   );
   gpc1_1 gpc1614 (
      {stage3_34[3]},
      {stage4_34[6]}
   );
   gpc1_1 gpc1615 (
      {stage3_34[4]},
      {stage4_34[7]}
   );
   gpc1_1 gpc1616 (
      {stage3_34[5]},
      {stage4_34[8]}
   );
   gpc1_1 gpc1617 (
      {stage3_34[6]},
      {stage4_34[9]}
   );
   gpc1_1 gpc1618 (
      {stage3_34[7]},
      {stage4_34[10]}
   );
   gpc1_1 gpc1619 (
      {stage3_34[8]},
      {stage4_34[11]}
   );
   gpc1_1 gpc1620 (
      {stage3_35[1]},
      {stage4_35[2]}
   );
   gpc1_1 gpc1621 (
      {stage3_36[0]},
      {stage4_36[1]}
   );
   gpc207_4 gpc1622 (
      {stage4_1[0], stage4_1[1], stage4_1[2], stage4_1[3], stage4_1[4], stage4_1[5], stage4_1[6]},
      {stage4_3[0], stage4_3[1]},
      {stage5_4[0],stage5_3[0],stage5_2[0],stage5_1[0]}
   );
   gpc1325_5 gpc1623 (
      {stage4_2[0], stage4_2[1], stage4_2[2], stage4_2[3], 1'b0},
      {stage4_3[2], stage4_3[3]},
      {stage4_4[0], stage4_4[1], stage4_4[2]},
      {stage4_5[0]},
      {stage5_6[0],stage5_5[0],stage5_4[1],stage5_3[1],stage5_2[1]}
   );
   gpc615_5 gpc1624 (
      {stage4_4[3], stage4_4[4], stage4_4[5], stage4_4[6], stage4_4[7]},
      {stage4_5[1]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[0],stage5_6[1],stage5_5[1],stage5_4[2]}
   );
   gpc606_5 gpc1625 (
      {stage4_5[2], stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6], stage4_5[7]},
      {stage4_7[0], stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5]},
      {stage5_9[0],stage5_8[1],stage5_7[1],stage5_6[2],stage5_5[2]}
   );
   gpc606_5 gpc1626 (
      {stage4_6[6], stage4_6[7], stage4_6[8], stage4_6[9], stage4_6[10], 1'b0},
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage5_10[0],stage5_9[1],stage5_8[2],stage5_7[2],stage5_6[3]}
   );
   gpc615_5 gpc1627 (
      {stage4_7[6], stage4_7[7], stage4_7[8], stage4_7[9], stage4_7[10]},
      {stage4_8[6]},
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5]},
      {stage5_11[0],stage5_10[1],stage5_9[2],stage5_8[3],stage5_7[3]}
   );
   gpc207_4 gpc1628 (
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5], stage4_10[6]},
      {stage4_12[0], stage4_12[1]},
      {stage5_13[0],stage5_12[0],stage5_11[1],stage5_10[2]}
   );
   gpc606_5 gpc1629 (
      {stage4_12[2], stage4_12[3], stage4_12[4], stage4_12[5], stage4_12[6], stage4_12[7]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[1],stage5_12[1]}
   );
   gpc7_3 gpc1630 (
      {stage4_13[0], stage4_13[1], stage4_13[2], stage4_13[3], stage4_13[4], stage4_13[5], stage4_13[6]},
      {stage5_15[1],stage5_14[1],stage5_13[2]}
   );
   gpc615_5 gpc1631 (
      {stage4_15[0], stage4_15[1], stage4_15[2], stage4_15[3], stage4_15[4]},
      {stage4_16[0]},
      {stage4_17[0], stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5]},
      {stage5_19[0],stage5_18[0],stage5_17[0],stage5_16[1],stage5_15[2]}
   );
   gpc606_5 gpc1632 (
      {stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4], stage4_16[5], stage4_16[6]},
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage5_20[0],stage5_19[1],stage5_18[1],stage5_17[1],stage5_16[2]}
   );
   gpc615_5 gpc1633 (
      {stage4_18[6], stage4_18[7], stage4_18[8], stage4_18[9], stage4_18[10]},
      {stage4_19[0]},
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4], stage4_20[5]},
      {stage5_22[0],stage5_21[0],stage5_20[1],stage5_19[2],stage5_18[2]}
   );
   gpc615_5 gpc1634 (
      {stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage4_20[6]},
      {stage4_21[0], stage4_21[1], stage4_21[2], stage4_21[3], stage4_21[4], stage4_21[5]},
      {stage5_23[0],stage5_22[1],stage5_21[1],stage5_20[2],stage5_19[3]}
   );
   gpc207_4 gpc1635 (
      {stage4_22[0], stage4_22[1], stage4_22[2], stage4_22[3], stage4_22[4], stage4_22[5], stage4_22[6]},
      {stage4_24[0], stage4_24[1]},
      {stage5_25[0],stage5_24[0],stage5_23[1],stage5_22[2]}
   );
   gpc615_5 gpc1636 (
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4]},
      {stage4_24[2]},
      {stage4_25[0], stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5]},
      {stage5_27[0],stage5_26[0],stage5_25[1],stage5_24[1],stage5_23[2]}
   );
   gpc606_5 gpc1637 (
      {stage4_24[3], stage4_24[4], stage4_24[5], stage4_24[6], stage4_24[7], stage4_24[8]},
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5]},
      {stage5_28[0],stage5_27[1],stage5_26[1],stage5_25[2],stage5_24[2]}
   );
   gpc606_5 gpc1638 (
      {stage4_26[6], stage4_26[7], stage4_26[8], stage4_26[9], stage4_26[10], stage4_26[11]},
      {stage4_28[0], stage4_28[1], stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5]},
      {stage5_30[0],stage5_29[0],stage5_28[1],stage5_27[2],stage5_26[2]}
   );
   gpc606_5 gpc1639 (
      {stage4_27[0], stage4_27[1], stage4_27[2], stage4_27[3], stage4_27[4], stage4_27[5]},
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage5_31[0],stage5_30[1],stage5_29[1],stage5_28[2],stage5_27[3]}
   );
   gpc606_5 gpc1640 (
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage5_35[0],stage5_34[0],stage5_33[0],stage5_32[0],stage5_31[1]}
   );
   gpc606_5 gpc1641 (
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5]},
      {stage4_34[0], stage4_34[1], stage4_34[2], stage4_34[3], stage4_34[4], stage4_34[5]},
      {stage5_36[0],stage5_35[1],stage5_34[1],stage5_33[1],stage5_32[1]}
   );
   gpc606_5 gpc1642 (
      {stage4_33[6], stage4_33[7], stage4_33[8], stage4_33[9], stage4_33[10], stage4_33[11]},
      {stage4_35[0], stage4_35[1], stage4_35[2], 1'b0, 1'b0, 1'b0},
      {stage5_37[0],stage5_36[1],stage5_35[2],stage5_34[2],stage5_33[2]}
   );
   gpc1406_5 gpc1643 (
      {stage4_34[6], stage4_34[7], stage4_34[8], stage4_34[9], stage4_34[10], stage4_34[11]},
      {stage4_36[0], stage4_36[1], 1'b0, 1'b0},
      {1'b0},
      {stage5_38[0],stage5_37[1],stage5_36[2],stage5_35[3],stage5_34[3]}
   );
   gpc1_1 gpc1644 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc1645 (
      {stage4_0[1]},
      {stage5_0[1]}
   );
   gpc1_1 gpc1646 (
      {stage4_1[7]},
      {stage5_1[1]}
   );
   gpc1_1 gpc1647 (
      {stage4_3[4]},
      {stage5_3[2]}
   );
   gpc1_1 gpc1648 (
      {stage4_3[5]},
      {stage5_3[3]}
   );
   gpc1_1 gpc1649 (
      {stage4_3[6]},
      {stage5_3[4]}
   );
   gpc1_1 gpc1650 (
      {stage4_5[8]},
      {stage5_5[3]}
   );
   gpc1_1 gpc1651 (
      {stage4_8[7]},
      {stage5_8[4]}
   );
   gpc1_1 gpc1652 (
      {stage4_8[8]},
      {stage5_8[5]}
   );
   gpc1_1 gpc1653 (
      {stage4_8[9]},
      {stage5_8[6]}
   );
   gpc1_1 gpc1654 (
      {stage4_8[10]},
      {stage5_8[7]}
   );
   gpc1_1 gpc1655 (
      {stage4_11[0]},
      {stage5_11[2]}
   );
   gpc1_1 gpc1656 (
      {stage4_11[1]},
      {stage5_11[3]}
   );
   gpc1_1 gpc1657 (
      {stage4_11[2]},
      {stage5_11[4]}
   );
   gpc1_1 gpc1658 (
      {stage4_11[3]},
      {stage5_11[5]}
   );
   gpc1_1 gpc1659 (
      {stage4_12[8]},
      {stage5_12[2]}
   );
   gpc1_1 gpc1660 (
      {stage4_15[5]},
      {stage5_15[3]}
   );
   gpc1_1 gpc1661 (
      {stage4_15[6]},
      {stage5_15[4]}
   );
   gpc1_1 gpc1662 (
      {stage4_15[7]},
      {stage5_15[5]}
   );
   gpc1_1 gpc1663 (
      {stage4_15[8]},
      {stage5_15[6]}
   );
   gpc1_1 gpc1664 (
      {stage4_17[6]},
      {stage5_17[2]}
   );
   gpc1_1 gpc1665 (
      {stage4_18[11]},
      {stage5_18[3]}
   );
   gpc1_1 gpc1666 (
      {stage4_19[6]},
      {stage5_19[4]}
   );
   gpc1_1 gpc1667 (
      {stage4_19[7]},
      {stage5_19[5]}
   );
   gpc1_1 gpc1668 (
      {stage4_21[6]},
      {stage5_21[2]}
   );
   gpc1_1 gpc1669 (
      {stage4_21[7]},
      {stage5_21[3]}
   );
   gpc1_1 gpc1670 (
      {stage4_21[8]},
      {stage5_21[4]}
   );
   gpc1_1 gpc1671 (
      {stage4_21[9]},
      {stage5_21[5]}
   );
   gpc1_1 gpc1672 (
      {stage4_23[5]},
      {stage5_23[3]}
   );
   gpc1_1 gpc1673 (
      {stage4_23[6]},
      {stage5_23[4]}
   );
   gpc1_1 gpc1674 (
      {stage4_23[7]},
      {stage5_23[5]}
   );
   gpc1_1 gpc1675 (
      {stage4_24[9]},
      {stage5_24[3]}
   );
   gpc1_1 gpc1676 (
      {stage4_24[10]},
      {stage5_24[4]}
   );
   gpc1_1 gpc1677 (
      {stage4_26[12]},
      {stage5_26[3]}
   );
   gpc1_1 gpc1678 (
      {stage4_28[6]},
      {stage5_28[3]}
   );
   gpc1_1 gpc1679 (
      {stage4_30[0]},
      {stage5_30[2]}
   );
   gpc1_1 gpc1680 (
      {stage4_30[1]},
      {stage5_30[3]}
   );
   gpc1_1 gpc1681 (
      {stage4_30[2]},
      {stage5_30[4]}
   );
   gpc1_1 gpc1682 (
      {stage4_30[3]},
      {stage5_30[5]}
   );
   gpc1_1 gpc1683 (
      {stage4_30[4]},
      {stage5_30[6]}
   );
   gpc1_1 gpc1684 (
      {stage4_32[6]},
      {stage5_32[2]}
   );
   gpc1_1 gpc1685 (
      {stage4_33[12]},
      {stage5_33[3]}
   );
   gpc1325_5 gpc1686 (
      {stage5_3[0], stage5_3[1], stage5_3[2], stage5_3[3], stage5_3[4]},
      {stage5_4[0], stage5_4[1]},
      {stage5_5[0], stage5_5[1], stage5_5[2]},
      {stage5_6[0]},
      {stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0]}
   );
   gpc1343_5 gpc1687 (
      {stage5_6[1], stage5_6[2], stage5_6[3]},
      {stage5_7[0], stage5_7[1], stage5_7[2], stage5_7[3]},
      {stage5_8[0], stage5_8[1], stage5_8[2]},
      {stage5_9[0]},
      {stage6_10[0],stage6_9[0],stage6_8[0],stage6_7[1],stage6_6[1]}
   );
   gpc1325_5 gpc1688 (
      {stage5_8[3], stage5_8[4], stage5_8[5], stage5_8[6], stage5_8[7]},
      {stage5_9[1], stage5_9[2]},
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[0],stage6_10[1],stage6_9[1],stage6_8[1]}
   );
   gpc135_4 gpc1689 (
      {stage5_11[1], stage5_11[2], stage5_11[3], stage5_11[4], stage5_11[5]},
      {stage5_12[0], stage5_12[1], stage5_12[2]},
      {stage5_13[0]},
      {stage6_14[0],stage6_13[0],stage6_12[1],stage6_11[1]}
   );
   gpc623_5 gpc1690 (
      {stage5_13[1], stage5_13[2], 1'b0},
      {stage5_14[0], stage5_14[1]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5]},
      {stage6_17[0],stage6_16[0],stage6_15[0],stage6_14[1],stage6_13[1]}
   );
   gpc1343_5 gpc1691 (
      {stage5_16[0], stage5_16[1], stage5_16[2]},
      {stage5_17[0], stage5_17[1], stage5_17[2], 1'b0},
      {stage5_18[0], stage5_18[1], stage5_18[2]},
      {stage5_19[0]},
      {stage6_20[0],stage6_19[0],stage6_18[0],stage6_17[1],stage6_16[1]}
   );
   gpc2135_5 gpc1692 (
      {stage5_19[1], stage5_19[2], stage5_19[3], stage5_19[4], stage5_19[5]},
      {stage5_20[0], stage5_20[1], stage5_20[2]},
      {stage5_21[0]},
      {stage5_22[0], stage5_22[1]},
      {stage6_23[0],stage6_22[0],stage6_21[0],stage6_20[1],stage6_19[1]}
   );
   gpc615_5 gpc1693 (
      {stage5_21[1], stage5_21[2], stage5_21[3], stage5_21[4], stage5_21[5]},
      {stage5_22[2]},
      {stage5_23[0], stage5_23[1], stage5_23[2], stage5_23[3], stage5_23[4], stage5_23[5]},
      {stage6_25[0],stage6_24[0],stage6_23[1],stage6_22[1],stage6_21[1]}
   );
   gpc135_4 gpc1694 (
      {stage5_24[0], stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4]},
      {stage5_25[0], stage5_25[1], stage5_25[2]},
      {stage5_26[0]},
      {stage6_27[0],stage6_26[0],stage6_25[1],stage6_24[1]}
   );
   gpc1343_5 gpc1695 (
      {stage5_26[1], stage5_26[2], stage5_26[3]},
      {stage5_27[0], stage5_27[1], stage5_27[2], stage5_27[3]},
      {stage5_28[0], stage5_28[1], stage5_28[2]},
      {stage5_29[0]},
      {stage6_30[0],stage6_29[0],stage6_28[0],stage6_27[1],stage6_26[1]}
   );
   gpc7_3 gpc1696 (
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], stage5_30[4], stage5_30[5], stage5_30[6]},
      {stage6_32[0],stage6_31[0],stage6_30[1]}
   );
   gpc1343_5 gpc1697 (
      {stage5_31[0], stage5_31[1], 1'b0},
      {stage5_32[0], stage5_32[1], stage5_32[2], 1'b0},
      {stage5_33[0], stage5_33[1], stage5_33[2]},
      {stage5_34[0]},
      {stage6_35[0],stage6_34[0],stage6_33[0],stage6_32[1],stage6_31[1]}
   );
   gpc1343_5 gpc1698 (
      {stage5_34[1], stage5_34[2], stage5_34[3]},
      {stage5_35[0], stage5_35[1], stage5_35[2], stage5_35[3]},
      {stage5_36[0], stage5_36[1], stage5_36[2]},
      {stage5_37[0]},
      {stage6_38[0],stage6_37[0],stage6_36[0],stage6_35[1],stage6_34[1]}
   );
   gpc1_1 gpc1699 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc1700 (
      {stage5_0[1]},
      {stage6_0[1]}
   );
   gpc1_1 gpc1701 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc1702 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc1703 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc1704 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc1705 (
      {stage5_4[2]},
      {stage6_4[1]}
   );
   gpc1_1 gpc1706 (
      {stage5_5[3]},
      {stage6_5[1]}
   );
   gpc1_1 gpc1707 (
      {stage5_15[6]},
      {stage6_15[1]}
   );
   gpc1_1 gpc1708 (
      {stage5_18[3]},
      {stage6_18[1]}
   );
   gpc1_1 gpc1709 (
      {stage5_28[3]},
      {stage6_28[1]}
   );
   gpc1_1 gpc1710 (
      {stage5_29[1]},
      {stage6_29[1]}
   );
   gpc1_1 gpc1711 (
      {stage5_33[3]},
      {stage6_33[1]}
   );
   gpc1_1 gpc1712 (
      {stage5_37[1]},
      {stage6_37[1]}
   );
   gpc1_1 gpc1713 (
      {stage5_38[0]},
      {stage6_38[1]}
   );
endmodule

module testbench();
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    reg [127:0] src12;
    reg [127:0] src13;
    reg [127:0] src14;
    reg [127:0] src15;
    reg [127:0] src16;
    reg [127:0] src17;
    reg [127:0] src18;
    reg [127:0] src19;
    reg [127:0] src20;
    reg [127:0] src21;
    reg [127:0] src22;
    reg [127:0] src23;
    reg [127:0] src24;
    reg [127:0] src25;
    reg [127:0] src26;
    reg [127:0] src27;
    reg [127:0] src28;
    reg [127:0] src29;
    reg [127:0] src30;
    reg [127:0] src31;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [38:0] srcsum;
    wire [38:0] dstsum;
    wire test;
    compressor_CLA128_32 compressor_CLA128_32(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127])<<31);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd2dc89aba3829bc2ec7be051f293a7c33a201d7b85bca897f20fad9f1554b8f0a253326ea1a7882d0459fddc1dec28bd19c146d932c08dfb40c205939d4a303e999e6240ac4edb14a920f518b364de91f548c8d327c09d3b3d10e9c5b5d859177fc70a842c79784b0d5decd7e097b4e3630dd9bdf9f990fce77c63a69b559e6076793ea1d5df5f7abb247ec1de9659e7346b08b6d70cf300c9b79ada6dd9e26c39fd882a8b2602920a4be4840dcbc505082f6e2c9046bc321f75d4633ec5ea22efa0c127e69b65d84786d9b1ce507d877cdc7451b83b83d79fb6fd56d54332b27da4872c6fc53dcb400e1f275f56efc83b9adfcbdabf07abba475ae285ddac0f75c972a41abd82db205dacbf453f3cc907ac31c96b6387886d16f167e148cc68790e898bd67f33b75683c20e6d47a925df74711c298139ee79d9ce751ea3975f4c4b379030c21e54b368b14edc3e781017f46fb552828ae1b3c4d35f4f48005a029ed2063181bb598513c03faa88fc33236154b7ee2e78df1c29082a953f91f9e6c5c779473dd522653bd0bfb6d1aa4eaa23423b610206e9885e8b78090dc7e045ce2fc65e6340a93d352e74db12a5f31b9611531da1be43737672a9120ede3ef74ba370cf03aafb2f42e333a65a623a4fb7e2fdf0cfaa81d65744723b845acb77c23780af46c4e1328fd8a4cfebe983915c13184b96470615e3f85e4169fa4f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hdf659c10325a350ac17455a3814d545483c978b31539ecf93105d99957798e3a1b2a2099d758ce3fff25853d34b5aa6b28977ce25a36fe11be0a56b53699b665341909403d97fd91c82e33e8ae6bb2a1176c52a9f0602ae9dee194d9e147a186d8b23923be759ddbf791d080d355de6d415f7de0451dd907b998aee27c06596131e7e7bc9b34eb9da721e606dd5762fee97f3cfbf2f175eb901cc548a70cc95b732e50c0c56bd202b202deaab4e66a9e990edf0144382ad1ed18ed59c521c2568723fab4284b7ab1aea4ff4fe8ec133b4f95f5be4fd310306eb8f131ed9d981362f79fa1305c314e7c2a401654fa0223fef89e723dc7b71af32c43e349e25a758bbd1a8664b59f12484048edea313fffa28e28956b4e52319775b9dce1cef24762b4dc028efad5221edf219c3f0981f5c436d1a20ab12c44c083f4530026f5fc16b2f655d697caebf8b4e593b32da1db3b4292317d681adc9a0ef5d5e2a020a783a014485fe4f1a18b141e246abcd15cb62bff87af7da34d6ef7d41f3283f11c2bba77ec75a2c35e31c195d7e935c7389cac117d378b31a6a0cec9edb8ea887f585223bff2c6cffc70bda86fa51a1c585e8e133d045fdc57966c403408a1300fa6ca99cb8902020d933da49f7847030b29db3fdb123e25825a4b3a11fc885b0f2781414f3421cad8fc658a448efbff7edbfa2c21a0f106b157f74028c1942ce3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h891919ff848c3e5336124b1a10fd394cfae638b261f9c7df87285f0735c7585ff070795dcbab0d59af7992d4cf4b0f0b7d56a3cc2f131ef70eaac8e6314d91a81197dbeee0bb1803d35f4647c54aab6c31f33edb85583bab973e972b09ae17ce0af5455697d386b8c51fbf611d9606aa9e84027830df7d2edf7118adc5bef7c81e4a0eb6bd7177bdc79a010fd332c09829a8895aa9a0ec8730343e439cc126d4fccd1d405049470d8b7db4b6aa461d77a381790b08f722e121cbd150496cb9d6adabd792b3b5b05873c6b0b2d4503a0ffe77130ec048a25328be8856fe4e60792f94ac355dabd964da01e36a06313e3828eba5c1638a78d5cf1e8af752367fa8cfdda82e098d370f330eae8e932822f16e0ea7a4bbe83cb8829356d78537a998152dd90b3e2936f6d1977a4f25ad3a96de6bdd49bc401d9998d46a7cb3fe7684d7944c3f2bdebd0e7fed9a2ee2a37455ba000f1b3948652352a150ddfe65cd227d7706bf33544cfc63a7540846b652fed0865a10f1c5217fbb778af56fc128209f47d5d776b9171a6757c01b46bebd2923673c5d8a3280569689ef1f5201a1b7012cd4c9a89be4e4cb416e529a701dd0af41d635dfa7bee90734549a7fc72224ed6180398276e7fa8a2760a93c96c68509ca158f874c1cda04086bb6bf55d51f93a17dc84740e47e990a1d38cee3d08de87d7fdd03bbc90c176e608fde1e6bb6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf018a510693fdbb67c31128c0656bb3938d6226870e5b5854def2f115e58c5f6e8ca76d6fb62c6a1478c3e840b53422f1aba4347acf67da7d9c02cd5596740e1f87cd7c79d7b73e7bd1e592dc6288a433e142b68bc7946bfabe7f678a2579b789226f198c038f244e758684a23f20e270568104fb90079f687a94be289e92bc02ab8882f618da1da499a73801c8454518572285cd85cfc07d6c53c490c634075ff210e483bf12298f676a70a6a1c4a0ef13f25f5af32e4b65ad547d2ec45b24c20ad8d428bb2ee99af8fd808dcd2b37bf1cd330548730455a722a5f2e57184823b2f72a9b9f367722a5976dc2d64f2c8e5af2e692a10a283b21003b7ed5eadccf7ab2de0ac6df0adb754d8a24b6097522e48aeb594b485aa9be146ccb03ae3060a318ef3c93770f42659ea61f48d25e6ea7cf463b0f712e9ed52ef60ccc448e30d266a5230093a505ab380a767e9d232d1a64448c0c2452ae3c165f287f0ef761c64e41a52c71c6b9e98f1f4ecdf1e1e8fb4b89af3e579ff383c9884617a965e8cd999ef61d10b5719221dfa6a0134e61451ef114837d92583256d6fd69146c7be4c7a6d6458998243c20d7a58fb10ed8e5a4c5b8dde7fd07a68cff3101646eae65269db9ae6cf91e934cb2cac097b7f0eeafeaa090d282f02a7dcdf915b8d8777b8146ec6050cff0d2ded930124d74c7d8a41603e0887548d92fa51400f569b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hfc187d23e7f2fa70e8b1ab1be2e61189bad50350c7693b15055f6b2849225c8165177d5fd8e8f8210c62330aa1376d802b3678b80e4c46b656c66b38419e5870962880ed74640f35bee1cf4ee0ad7a608c3ec5685208c5362d59824a8cfaf06743b7e8e92dd2fd583ae46d15311e5f3ee71ccbf417b6818c4c9798c6c6ce735e40fa50db9bc7f87836ca32c8fe7924b29731d33cf42b0ee6356423a9c97c89c76f2b868ea509a29fc59ebe9b293905069daba8601ba7579511746ce78d8b8cc553e847f220933215d8ba700dc6f51ec4123347ea46ff6922418a719feeee287da5f34a3ee3d25ce53130b1fe4db13d60b8f57790eaada84754299dd522af5e24efa70cf288b212167b13566dcb6a0ba32c40cc0e1eb2dc96ef9205fc01ba3b9b2fb92c3e7d6393b174c821542e280489323efb514a5b7e25f813e3896a8dd4ce1e091f1bfe29d098e3467619edc92b7ec51db78045eea4266a675fc26842f1af97460723979b18134280ce906fd5adcb92cf3ac7a63ac4e27828834b24378eb0c47f99497d29b9a88624413bf99aeb56f71fea660904811e211a7fb83ea0b8df7837e910419fa705996688aed4af93179d5829abedc82057d0399e59137196e9f29688299d43866784c5e31c7c16be724c113926272fb028779b224f7d38aba13f7a9c4c187d3c2b5d7ec375f31c1f5bfdbebf4b52e6d74319fcd4a3ea309b1c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1822245acc0c80956703e9f2df18a46d67e056b182408e005afedd36fab25c77ecf0d5fc7c6c83afe64a6e1048f32feb7d1235bbdb9fc012884c80e91adb64ed09e11fdeed9660da4e4a485b5249acaba9af47c75b9ccd5df9e88ba3724fbf11a675e21c8b9706ba487a9f4f87e09665e686a50550b2f4afb3a51ee0dd2b8dec42949a736c3f89589bbb1c5a8b9479e8d0d3c9533615586bf5912334f237773b7dfbb8564596a7c3dfe232ba5b24ac12f7a3d781789535e1c1493db5cedc1e6400597c98b81722471ead7a13e50b5e2b96a62941d5286ded6e3e22f87a4b60fb753379ee09748c0f88a183fbf64474e87d7caf66f98e0ebbe978530e7439443cf58edefff9ff682a213a46128d91a8ef7cd4e928819a936573b7b86efa8df2b6d5c9ba783569205cfd2c70217d00942e47c01d5f5796ecce30006adea0223833bfbede2fc61086652b0a85a6d9d58e2f4216a4ee98fa67933454036866f9f1ad5455da655f52fbd8b947ebf6053e12b899d4d163678ed0fa12755549b98c30905b81abea488678ffaa89e183ddaa945f95607077e9dd429488cf3373e0e0632ca3ab72a35d47faa05ea56cb704795f5a198e116e9135433c55990f7bf0fa6321913fa8c6821b62a77b5b75131cdbecaed0e2f3c5d55132552279d97d1af1ec9b86e4c3c169d5cfca34208f513067f2dc734ad7febdef83acec6816857fd261f6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5b7d6509dec8422b2a41fa85ffba38b529f03f673c1bc442ffb4867ea0f666cf0a592c52e6db1f6fb0a8443e537fbf5a60a547b754c8d971c8468dca383a3c062fabbc071d3a42456905e2753d46ce3fc3da35a7605065e7a71017fef3de55f4bb0a4a5b44484ec802293d81d21df4c7dd559c7f6059c26d2fff48157990c974206fa5e40e7bfb5d020b5306b8420c386eaa15773b40e3f3be8db4cfc089276dd0bfd98125e3e1872c1c45fc48309ce98d25886c59fb3d0807be9279e94cee9134ed52d9de63158a500c3b82484c67663159bdaff14c885b0fae91b2b4e090e993614ece4bb204f8862d3672cb04a1fa2f75a209612f4b5ebdf140188e01ec57203b9e0c83f437833310f7b5c2c92836f008de9d46e65beecf85e7c4335dcae994160fed3206f09a2f98de95a2021cee764fd33bf90c28dff851e24b6fc2adff35e599edb616532ed5e2d1000a48343772a91f6e8b76d9e494fbbe7dfd1d09171f1564af75d08283e2e42de62be602d711dffec884195b14afc886824f8889e553545d9d27e1093adfc481bf0e1bbbbb50397d670709a3fabce74481b1f984072d5db93203a97c2161ecd261811c7cdd58e99488553e5a4e49dfcd5b820b5dbfaf19bb7dadb99f72c464116ea721994589b0dcb4097800056c20399b93fee75c6cfc47930e5c865d1241b3a5bbf9485705c3234f5db79e14c37ce01d724ed18f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha440d108557431dfcc47fa417681b4743e2fd40cf815596087859279ec0ae823332ff908e4a032b39f657705cfe63e99e9928e29bcbf44b6fdb4b84b0bb216f86b7c4a6f860a097b5d4b5ef795f2a3c036c70eb42d4b44b013e7a20253c4c74b4089514cc6486d49ef0255a806c6e6879d82a643f396f6a72067bff4f1bf1f3b8a532423bf67e631399d1abe75e363695b5d08b04ee34ad2bf262036e29b468f90f89dc8ea52b9d83d650614d97fa2c286b58a96148d882e4d3c5f6f74f36ca14bacf540285dd4023a2d902fae202e2157bdbe5a29a864a074a116831b9fc3d8faaf0390f33448d2a749f58403e44c1abfb645b0ae72fea710b71491302b50e06dca585a70ed3d716d5d96e2230c8291d8d94016fe3f7f4996e08d56bf2bee70d92bfe08329663148e5705c8fb2b30a8ee7d255c04422a05408489b689301525e2dd2f05e75d485e0504bb8a8ff86d3d6917d7a54b9bf885e372df90448fbc4439977150403a1590b05594927839857165ab5287dcd2d02495fb2e0d7a7e5a7ce4bcb3f93e7d003e256c4b9fe2eb0809d13b93bce8a8f797fdc5d35d536aa96ad015ec48580b489208daf72985c417e86c2b68e4af777cf26f2888eb18737702ad9367be6ba6fa395e457f1e6e4258cbc3ff8cef458639ffb73997ec3e9b4856d84184a4f40baa7b1737273c6c2ed61b8a493184e6f955a733a76e0d5a2ad8d1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h61a943d30c222268c2274d40f9d1ee7ae51c7666a31e425839f17cee64424ef9ce75365afae144f9c65df9026406ad0045d7f7bdf9eaed2442c2e50da50926856043aab4ab12a10419d86a09bd121e776ac755f332edba41ba06e726dbe041e5c95bfe20ad07809f7240ea1b26e857fa1aba2c4edd3e1b05ebecedc841283a8321a569a56fc5c6b3d53ac5ee8e12cdc8885d5c55aae0ca43435cb40b0618b9fd0d860084b864299a69f390588a7df354407d97ad6b5577541e56f51958e0ad96b228c16282224a22f4ad2e89662b32a8d49f8ed776628a94f744e28d9a97b11d7af81463713c418c77daaa04445ced6a8eac9501febbfa0a6ff2d7727a265be98e02bc23ad85bf79be29ea5b19b045f1c6b436a48e6423e5b4764dfdf096d3f142ec14dbbc6fc3fb19683f328e5072cae2a5d791de1c28ad5d8cae1fe1aa99c6ad064a3c234ebbbc929ffd054c7a514cbabf06ecdab23afe590f69050d99eb110cc8565e4b5fb22176ea0f16b885e873790da14a4597c51be258d6dc0ecf5df6fdcbb40f0584184b8539d50a3d6da6db265f37c4860195b35ea6a75126bbf608db90856f3363ccc534fcfb7769f5a2fa98352a9db3b17ef82c843952fb013dd023503e542ada0e34a22866f769a8d4d185930ee57b5208e30690e2a01a8341575a69df000e14e12f3651e02ccba6f280ee373265ed10a9bfe086718ca7c1c929;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3ba66af9a84e2cce7dab92d65d3ec9e7e63132b52a8b7190de56ae2727e8d5de97c2672fceac6d5b36476a432660011c32b6bba516fd95d45ffddfe9d2e7fc6b99ebf8134f1c4eebc61220e149eba255a682f5ef6dda480411f78a7ca056542fac05c9546f5d7c5fc74bc142e89576e0dd2f22a09cc9aebed4dc146f9f08e83f1fbdbbe15f5e34aeb036422cec6a50fefead5f277cad62b3c0d063852549d1e0e5ffaeac4d39b5858ef4777ed007d8f1ca42fb3add64c7b93c14f9f55d199f4fb0965d9889d1a559efbcf7c4b569c2f038c0ef35a75c24da60b334e357fd90346bed2f09ffa887602b82371a1511db9105d5a249042b416d129cda5c17b2a1cf36f3f0518597cb82643e4e1ea520f0cca6fb321cfa07b29a4b9e9189e51825a03361ed094dcbd3c2213b9456d6c3b5e7d9f043a1dfe39f62c8697be9e9601d361ef996bfab2d07d8ee7710d1204ab5bfd213d39fe5bb70c7b77506b88e513c25259ddf3e54a5263b5cb78d0984c5d3310d077e5be934afd773d6787d81681128b8331c7af0e9b31326ecd587419db2eda0f6f403ab61fc85e48c31ae73e53554173871c245e61fb0d051fbbad68a176b708bf4e7db3020c307e6728f8671f2e7b12f42a702f46960ac8b408f00fdcabd910e04214757816ba398b07a33dc960b82c89026b5e47e051c5bbb7495d964a8344e267bdcec3ee0bde6ac5a966025ad;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h51271903fe19fd686786b92142ed8db9221475faada406bbecbfb1d3435354a4013d40d2762e2ce2e659ccc602dfe0e8dd07578fb6039ed89fdadbddc46d51736d38be0988323dfe54521dfd6a171453fae4a636d6c4975ba4c2e04a2c07d3eef2d97ea6fb8988a6fc09dccb7e13e58dc2c3b1135f2cd70c95a452ab57bf7e9d6cf9a15bae3273996d80f1b09549f2d4ae4911dcba6680706bcaee6fbe001949565b71079de02a71f7e04e0e91f4b4c4e02a9fbf7b7250d32a66229422989d886da312784db1b7cb44ca385d1e2b187b046803e7e950c68ea530e4cb160bfbdffae06bcd71850d4b324ccbd11102d29e7071a7ecbe4de66daff8bc4e6e5bf6f4a63b27463615ce716d9cc63499fa5dc8f94b3de6e6a92b9cdd5deea3e80b14e2950fbc12e4339ed2fb9e1815652a2bacace51e3963062e03fa03fba588242c4be1c1b3664ef7021ea2995c9fa24ff0bf1b4ab2b8b605bded77eee09d46e14f4d00411a6995e62161f88442825280a81cdc199b42e019e79bd66858b08ab40be01e189c1d4951cf5603f3c86bba37ab0857fc4b8284a1fe1f677c5d9b252387c067957fb76638ec3611e6c34328c744a922745bedd7e0a1ca01ead872d6647b3834f6afd8c6ab8118eeaef563cf1e83e8d5f30740eab0034192cebcd9c936139563080d76e76cfb4d7f5147724dcfaafeba9d5779510cf40e95322d12182d2ec8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h12c67e86df12cf465bfe168f0ebf0d45e4530b148d66148e07846b0a1d36d96b048f4d6b7498043e00b582d73084ba07380cd872e10cfdff395f67c8baaa3efb80ef9ff3ce0af8b6706e914082a48e47d93a78382b78d917e5471aed857920aff31bcfbe24d2f7ed2d939b66c308f4df6258e5d8c8e27de9813719e6228ca555ee3d0e19d46b93d773b4489440868ca6cdb4f540ec0168525e3ef425459270c5e4b7145eedd111d1712dcc447406da2f02f695c200fc329e134b65c7c73ca16100343854fff332ad12351164a10e838b74992b1c447ed9dced085c4de44fa046a7693d5b9ba6e3eef6dcaf771c93429daca163b20638e37decbcd1c50307f7110eeeafa06e15b8c5a1f4b5232d7542f2a7e8f563ea6d8731c4e115ee3b61b2f0d0faa61eccf7ca20d4c504b7618e664a14960d268fe8260e057ee941ed57904d38c26a263e14439a42b71a70cb5905c48d779fbdbd2dd306a6943f2480fe1e294808093f7ef1701b4eaf3b268b5bdda3721e8dfedbf3e8dcf571d2801d2ef8351250fbdc1e69de7de509460e19f3e6db5046dc28cded34b05c0ae96e77ea608c01142e2f3e6662c2e0a236867978d303f488a43b3952ed94a8b3b55a88be323f23fc897e1193d2fd1be6e94ffebdf374059d3848bf4c95e549c9d6bfcc408592500c4efc871ad7b7ec5caafc9a862cf10935676b5762c394496f73a32a7b05c2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h876d94d4baece83ab831514e09fa407c4de817a7c6b7781e4b308686e15f3047f7e83903306896c123ea2624791a2078c806a1ed8c76c0534056f1329f1391e4b302012400d781855f292d065fb9874ab7964037bc8d0665377f728f75be20e8c9045878dd4a9a07114c0c43a639dc4d7252b4f96dcdc51e5f4020b8f3b230165172433d803cc6b34f199f2c0b08784d4349a85d96ed742aab6221f750bd106f928bd8ed3708971d1a447351f4dd7bb94979b04190a1e7bd2de67ca162a1d60aa7008ea5972c0995d39cdb4bdd79242f7878bc0ec493e3a762fa90e78f25c083c241bbfe320aa0abcc64a35c20c1d5fc9aa6d5e78555af9466c95e1deb2299019538b3c031551f32893948543fdface0cbc761739fb191ce6d4abec467e83bae780f539a19b79b3c0b18f0d7d886d3149f53d315207a2e71748e1ab44fbe8b2fe7cada148a64511576df547241d0266822bf1e038a38d2b7c8c1fbcb1f414cd249f2232c43e3ae28bce273d707c250297361a3d961a248a6f21b4878583ce71736d4666bb4107ba748120eef76d4ecce39518aa74468a9edc88d99bcec670666af21985815e1a7afc0be3f22818b72bf51d9fd6202485c3124d599726ac03fe9ddd1fd9ab2727e9fff70f4cd9c813e1f118ccd6e399a3e02e0f3f0b2d3fb73ef4c4a919f56fa1aff559fd42fa2f5474fb7a364ccbf4ac7b5847ea916db3c6e84;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb14066be32655d13fa5229b7c42fe5f8b185a8ee4f02b3c46e3f898fad3cdefc975f8e440a681110ae3d526450c51c27486d33f911e693b3bb2aa0ef22260a10f4146b92e6a8e9fa55b4484f835bd45400189960bf0635b6df7c1edc18c1b887d40d6ea85b6d8397f4ae8bff8dbae4136094d29ced0d834a9c4a71e34a55ca9111831ddde73d291be7ee5ed5e61f3b481d78b0521d766be167e0853b7a92317c3ffb157c8b3fe58ddb0a5a83ebced13286366bfe109e0dfe86b466cbae96ebf4b1d5b346632fa2879c9f56fc85c3ab83d6f14dc2cde7389b21f64e09e0fc9e10d79d524cf5962039a919cde8070cec47065b62638367da130d7e4cce394b0d7d4be5f4a0afe99846c545a483282a6c76e5c8829381880de5364e7e21c793571dfaa80142b2b7dc044441d37bd1a5830ee41613f0039317dc5d5e419582424a5cbc6a3863a4d9861a1de475c1be577508950a39a88d5ef5d5068e213a1a665f6b919531090c407710695a731f7c03eac8359c40df5feda7235c2d3362a21c60bec3f876d23f02b328be70a105d86071b2bc3d8f4cd99f8d1aa64077b4884d9c88a3a67818b1a3175cc632abb75195cb32dee7b7d1085cf13f95a88a67c42206688cba050eb5946b6f31b043e02e4acebd76f59e8f8c80bca15a8199c62c1f579e3a8a6bca4f5dcc6e698c03619f7f1daeae6ca8f9ca2df2126252357dafaea06f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha663b3ff607eeccd8922cfae6b57f71190cdb8e74a5213ee5eaa2b527117223800c1201628ff0845d6994e47036ec50e21bc4e634a20d53319556709f8803505a1056c79efbfe78d4bdc92e9a5d8ac7ba730b956dd1e4d7a8f6b0f4b43baea2d3406b4fd8f3b49375a4e785a9d122ac468dbfeef6a4263881c2efea579dc2cc90fc5d01ab716f6cfb9a68245d99497e2a525b9f87695afb3246838fbd72791cb53ed9e1783409111910e1a01a56cb9a0bf069e869259d9d6a1fbda2b2eb1101728104715b82d9c5520ccf261bd7ec3bf8e8251138650c616a358e3883266c0d862c77f2b8b9023007de59952ac83d22104d700654333b6d5cd02549a840afbfb15d200d6f1456fc9d9912d6e8b14979b8569763a8b002717b961951410b2d61fa0d2b75781757a058c66a6d3ad33066e3c4b62674bb36eb079d9eff737055e5d151f778f762a29f95fd2f4157b90029fef379ab7b66020c84ea209145b7f7669c0b21714cd8198f06ee8633e6a83943e76264f908ec9bbe7d098834beae85752ef24143aa08a804e2b37a110c09c719cac86ebaff43ddeeebb0bed772ed209cb6dc9879e536f1666d139f1aababcf7903f91cc6c7ee7db246591b843c69e670a2bac7cdc77914d5157bbe763d41f4aa3f768ef80779d631357c7b09a5fa8921b44062ff81e565ea2b19621b43955b3159c415d6460f56d19f43b515859af06e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hedcbc5e1c9d247e5dc9e4dbe3658164ba9c4c8a63cd13aaded258746c73f2d65810c45425446f5441db51a671dcb5bb5cf20fe12e35244f188ca6ff85706806ecef896a62b9cc9c65baf0f7468637cfac5a85bd9fb641e616d819aff5031a4dd514b631f7c70b408e2d7d52113b5da36a9a827181c67596a754cd8099cc295ac24c332c935bfd3f0205d34c269ca15c71382ebe35446a378063f345c912e2ee2e731be30c49227aa70bde04ee22a7001f0ec7553aefcaea9e6c1c82988b3d17edb769716e08c8f7ee55bf5a78bf1cb5802e4deeea0c6e4af237d479245360c0e3676106bcaf66aa991f865cf196c109357e56e1b93b2afeb60cf624e2d2f4a00c0e171a71ee6c24323c4723f303b98ceedb57babe4231c28cd50393913013823863b6885226eea105df2e9958c58b9699d9cc67d0b30d3c5594a58ce978689098b81408f3c74776dac17b190a3be6bb44147abb69348a2f5cb3e371a461a9d77c0f35cd54a6c5a7ed1e9aabaac7b2e2701c13bb6efc5423ecc9771965ce7e796b7504829bbc7ea4328a87f17c8a58bb67a65606113d89396c39acf9b9e8569cf78a76ae4461a3bff9db6fdfbb9591366168738ccd29e2c365cc4715b9f5310049694c456d5c35d2bc1b5762f13bcd285a396d88c174332d7440837b21ec8db0be918968d77549f89979b9d76c7e032b118b20859746cba5490b9a4fc6a46fb0d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h15d5d33bc71b22a0f2e41430a95867f1385a2bd767495c811bfa763d62dd8057d675b025146f44cf74fefd89ea4c5aa935b0e65cd29ec78ee96451161a2302ed1d4932313218d42d0adabcc1ce2529b676655f183aebb5aab2f02c4730ba479e452279002fdae1d527f916baad5adb14dd023c1fe71254c00aa577e04d8784b7c721752562b3e3be3716fe69cbe7eb4b20ff53f4aa9a93a5bc401d31686c033230515f1980d8e7fd0c339fb15a7cebbecc29ee278be5bda8a4e58ccae1f0d38b38c976305c40c538e3a8e25dfa14a872136ac6130a986e3bd0c09036837f3fb1ddc933384b396ffd9ab737b9842be26f20dd08e5fabb98187852d4009aacae738fb8fb11632801bf36171bc91cfc6dd9ec45f74bf44789e3c52d4df2a99ab4f56821e0abff9a1a3ecf0ddaf7c27251cc890d4c26ceceb8fdcf053b86f2a5138563d6e0b64cd6c806c4fee168ee0afd79d6cf9aa50a09a59862e8c2950c9faa0f4100f63d52707b134c82005896d5dc1df171e20282b2f5ed62493e2d912a95c137ae11e494f028c8e80873b14ff094a6d7640b18e645e2d334a84635e87ced8276b8ea79d36e623c9c278b83cefb996550dbd1339000efacf34d438df92eb36d54c4fcec4b01d7f81a5e0f10e8a56da2c7d1c8ee493e1fc61c6074b64be8186757521e3d4ab9c73b0f8a33730cb9981639f651a043ff89c14688d5357a917e8a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1501fafa5e0212c6858edc8f50274ec20ee6e4930ccbdbde2a540f076371dbaf4a5eea2962f99bb716a9a7d1737c2c91b44537a09d7dd44e19d5dce8e42d885415bbdc03ddb1fdbd190a087136810d42ab1571ef7ad2a5bfde3715fb03fc6e105ec43f31f90dfabc5aa6e962e9281714577a53f7dfe4244490aadf23919c0b7880aee070e9016e4f70d6e6f59ba4d6efb379d2a13a7910a4501b640f73228a5ed5e5a63e7109fa51591d9b48467d9c6d80a29a0788997dc3619142eb490d33416cdf11227b5b3282c3d0664c5e5b78deb17c63e1259db232deb685087c839c879df3a7e2b4fb8c9dc6226740a8ea6916081c454734ae1dda23376738b92669f8d86e1e8f2900f06fadd447e642fb8156839d33487d958913cd0cedda31728e9082ff0ce40536d448303ce2323d74d857a52907024996b7bb32f4e1038568d83493cd1761fa89ad213a641a3a74597b6ea16a263a8497ef46b155387e1efa38fb2496d804b866ae867fe0b53b16782f0d649d5954b018876df614406d704346983ebe40160b212f4bf61fd06049d8c0a9459849051b0dc080eaf5f06e1e9969a0a7f0780035f2ebe8333c00376267b15ccd6d16cc4b4e92381ecf2a161b284fe67d4a861a37132187ed0b0ef0908378a96a3b6a4fcec55a2fe2703fbd2808b041050e8e852527bcc4f5b737bc17dcf2e28778262f5c42cc134fbbdb7ebb2b54f8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h57bd2a9023083debc4eeb4190da03bd745e03443b4876f1eb148280acc78662b609a676bd9930a9cfc15e0d10de9698005bd4ed60771db1ca65a31b92348dcd937eb49ac154563a262744a3b605a502829d6189a78cb2fb716592a4a1e1affa4c109027c1034b03f5c7afa006a477a595185c0d6334f479b6b2b0005fc7134810efabc8760cda89df17842805540d925af84e6f8f4d5a66629025708de5cfa05e61ba6126df639e34eed8145be0273a10d67ad547c7709cdc7fc5f95c8661aa4cdc1afadea93e1f62a50f6cd0386dea1b253418015c15397d1930ecb20b6aebd20682c9165b4786c9fbb9fe98b23290ec9de5d7ce01ba326274618999f362daeb2ad0802a14109f2e108917a91ef1c1348b3c4b409dbe24a729548ed2a33575335523b442a8c87b0aecd668e728889fa69fa4235add599e4447d38dd96451b551575e3c4d8f89341fd3736f07ae17301b3ed6418593e6c1702978d669f45694743564e77e47d31a8aae7e8e7b69a0c1a485a0f33770d2186e44893f82f9febc38adc10ec101f6ceba759119b1f2cda7a2a38e0b9e604d8add894d569d6f424346223b5cf5cb0253bffced868b8115b4b97cc33e14ba11c2308eb47a64794e0baa939d2b92a8ac2c1c6ae64c976b2bf3858e8271ba86890dac711a053f8c26dc7e69cfa36257509a1b7abfa46fdbac8e64c897df77bf35ad96e15816996df756d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h368117c5efe586fd2f9aadd49dde4f7e636764531381a8589a740ef704ae88526766b75e5bdbfc489b6c92d3c4a53a7dcf2e9c267ae1fa05745f2c1366eee55d30d8f399bcd1f301f7eed9331f48bcb4d3e538e9d38fd07dcba70af187b78ad0e8c501d8ccb19c0a71a9c35d7628526a13fc61d462b2eea32c8556f33c8fb5f34d0d0d49529856e95df15fdacc53162588d379f475161bc087be21591427212e06569eda34702496a449f58c41c3369d18f8702021c11ec5290971fb90acedcc2cca8760a3190811378c8271557708c7129f5cc89dc37948b733829f7d530812ab0c65168dec962a5d0b2d5d69e13f252f17d651b7000e94a58e6dcb8b891d37037d92a0f9ae35678ac8ae00ebf516c00e92745be0b6e50dc0c673cb3d0167a01c321b27dd79f2ca75f71f2df99912cf8cb37f6669d83e98c65eb6a7cd3b1051bb04bb44035e6d0b3f5470a51d5e6caaeaead4d88c7694941111b7a56e4485724ced6b36783867efedce3cf5508d89f37282e56ec5420d5dccf1b0c8691e961f536389c3cd10fa613041a9f5cfbafdcc7b085fb31155b4b89964f92bded33bd7b925e60fa3b846f77d144c7c38fc4aa411a4f61d30e86ef5b3ab7bb0aec02510a1f091d65fc5ed8e69554507e5f3da3b23206b327d682faf4af0970ea8b935d62fa809e25862f09d82f35c1ae9cebcf9a17281c99c9a31308aa1d3065f25710c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h67d4fc4e9c9aa5b5897dab10297bb386a685f30bdbd6c10d40661796ddf2cadd3a503792f6ea3650629e525c10c940eccdb0a5ed8a72797b1d1dd2960536fe53a9c59d171cccf12ee1aa0ec66a93f5bfb338a8147e3f865bb4fe7431abf23111ba07ecdbe2dc5722118861663722ce9ad38c03a55202ede62ac46c6e411bdfc98e5fc3486e7f547900a784f18e1f9b903ce732af236b4e8bfc52541c42a70ff2b1d67179fb292a1d94385a13e9f50c1814622851cba44a356e7a1615d04043271226061edf2c6eeb1f16cccc6368b6011a42fda3ee2e68b12f1e1bcc5afd411685244bf09803ac279bad942e2f4b52b8608adf7d953ec900c3ae42fd4caeeb4d78994a3ee47ab221986c84fc0b8037817cbf42da46113909011998e0d7d91ee4ba6cb2c346069ba4ed71b9dc6f148b9cef5faba8137da9519f97a9ee7418430d0bcfefaef7afffc24c6dba68cf88401fe25d06a56373c7e38c4790a1b78f13ccdc66186e3989edc7d0bde3df12e83fd7a2376c8c5c12cd6c485c0d1a77933c3e5e80707f33f231afbf708d939216475d8f674b1ae8087227f097cd6d2620c1b3b4e3b5478d265ea4ae199524e0dbf371a0589d669724eb240209b8aa2a47e9138a9b1ac673ab220769998b34eb8c1b28cca8cf75e04c93f77048ad36d13de2f191d5e0c44bcdd71139159cb5afda6f192b59769430457422b4178f76dbb24c0d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6ea6a7c83423b4104c42393f19d0899f1da72e074d7cef96b84cea9d55a91ab6f54222f1f2b7873a4be11fa1c4e972dcfe0a26d8fc15f90f501c9119f1685528c4536ecb76684b32f3d84bfbca556d0725cb24bbba9da1f471134ba84c0d85c2d851a312b6a401aa384d9c0d923c5c83c641f5aa0266e701d8a68d5fd1b6f1e177c968a6066390d197a8fe30de1daf67da53f357c3652e253c02b1ec34679144bc31f843c7a13de9d9f634b96b74a5850515deeaf634051a1b6301a6876bd5e274a97eaf197c72dc7044403b9ba98b180cb8ff2c9adf21923de68aa9e27fabac856953e3dd4cfd2a0434a2dba6dda020f734ad9a015033779a591e73895b0f2dd7fa66aeadeaccebf289cfb501afac116ae07b67c9f8c7fa490d9184c17169b5d5c79de0312b49e421b77f269c5abffa44dc3309067b20fa636157889fe76edbdd99166b45f5e12e2a52be11fce4dcf17333c96f3e189289f387445804601dc5b9206d4eb603eb57edbc9e603e7fe86ff494b70ba152948615545f5a614ca26ca4e82e764c91557d21641f8b3e21018aa3ed8d9c7be6be72affa3f7a1a0f9eebfaf5e500fc81785b4606a8ef0562b55708e084c3d044d8e3fa04e39d6e9b9a14b5d3be4a47aadbed75e27b81d011f2f005f8e60047993cd3066285cd36ba2f4c156f7da64c33ba0ab09cb333f40ea8b64341245c19234ecddca54a706d029b8f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h16b9e1a1f9a0c6effdb4d86e2c7d34affd93f7ebcf59d2b44dc05bc970a7111ec853c61458bbe41f4227b2459033dedde2c2bb43ab792f80d33026d5f5b10783c47a31a0c41cdf4440e0a9ee318416a3ab0d56c7a1f2baf926cfc05a0d7884d9cc3132b30f5f8bbcc98ff2f5c3a0a59d589b7e0ed3ec2192c9ae178fa74bdc468e4675a67e7447d04c9e9e1a7492378284b7be49145089962c3319bc2302285934550d0bb269e7119287fb4075e41f9411e30ec995788248c4b8ee810417c663044d83f7cf420727b376608b9fd0c8ea83c6e09eaa3b7638a116a70074f12a2974a68296195f4ede62544e0b6438046a7948dd77bdab5d93dc63e9697cd3b6ca4e9b66a4d0b0c24ac369804e90b8dd42b6b83d9f71fb73ee8c642e2038d3461e090f0eedcee7b1fafdcfe0bf6914f41713b8c4a245f98b65c2ccc86374212528b931ce939694d457c2d351d5d9c524ac43c892fddb654a2ebb93d0404ffd9a705118e57a0c2fc417451cf18ced6f641e702c2c34855bdefdb904a035592ff5d6b8df4bd22682d3a39d53443b1d325f6baca19a7b91aae55b23070c8279d92d2386fb614ebb0960d32002e72ae392f40ccc2b8ec69051c118e110ca1b89f356a20c64fa6c69558dd24b39fd6f7e0367c59e300630491644ada897af7c7351d61d1c87aa0753596bdb1e0bc0ad7cd07c3849000e7100ee43483352fcf8efbd2ee0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc26de1791e5b440be1d125a32c8f889bc3b2e205d05f27658bd4cebeb42cda29ee5d1d5c5ca7a8c028513a0927ecc0df35458e4edff9ee657cba0b42b16ab2cf2c5b4af516e76452c77f344aa33d6472e129cf7dea0a2f49ab66e18f1b793416dc6e19aade7a4ba79a8722eeb34201873d35bca6bd5ec8b6ffa537e279a9d594e093865847e74da062373675ad630bf7ef6b539ac69c2cf798d95fc5c36784f57226e153fb8a798d54dc0fa96979bb8c74f6b1273743de91a5d55963c0ed06ab11bc8ca4b614a1afcd92cfdc4af396d04865bb06708aa5ec60ecb6b66e00f77f8a82b87d4bcda3fc9ef9e38e021bafc07ad03dcfc7304d7014fe208515bfb58bf14234bee2cdc75ad1929064348c3b85eaa0646727cb07bfa531a13e3fd1a435896c71305c1e1dce18390245c759ecce4170d8b2c470620f26c7bd901317faf37fa390466ab8a2429fc346417c94b76b16d57bc6e0b797f6e913d86b2543a3ab5c4d72693e3586ea00e7f362497c9d0aa9bb3cceac5665c7f36ba74414b99f4eec4cb615401dfb380795ff4353983965548aa946bf01cbd3ae056eee371ee58c5cec12826909d35dd75a4fe6a04c8fd6c08f5c2a0ea088b5866cfd8d8246732315ad1d699d0ab1a102e23ee092209cbb4a836843d8273f48d7c8e827688d1f328158a4f7e336933822b7ede466855725a46a42bbb4edddeb0a3226791d7805ac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7bb78af2ce78fb779b3bdbd36281c02cf49fd87b115cf45dee7a00514765a6513626016fc1cc8f459e90c1439c44c9a05b8a589e20ac4bc6e3dbaf9661235c824c8c5613f6b64fe295c1dfc1f4a6b90b81d1f7a1425f9aa9ba4288f338439cf981a7b86d240e549df3fd701913f840dde1340e34db24fe92509ae4297f63410a8b7fd11c1acb5d6d5f63d251636d3d8f25b6cf75900778ff5fd70015c73d73f0cd10e8cf95625bc1f20a68a8caadc0fb58cfabe5bbd9ea2b436e1b126a329f0ad25c6bfc4a3e12599075b98872a6332e59c6fac480ef1bf107a136133a42ec5b68fb65daad8382775e3e58c9b283e7e4cf2f4c8a10dc28e16e0d07cbb9f2c5b028e58fad438140789bf32a7ad10931629e995ea4dabf8920dbf9306e7bce20c0a4d5c6fe665823487d64ac60bc1e5c3feb026a235f8d90ca29b86c98df6ead64146034a0c6b55c81fc67f9823596402520694207249dbd23b3f2f76c7b3f357d302e98476cbd314e88eb27e5e6e1135fe7ae1468d5827fee6fd58b72615a8fa7585f8e0fc92dab4625edf95f01f727099ef68c9012a75ad664921bbf4dff58e48665a0713a37297d009941961ffaf886b434c9c1752e94efdd458541c7ee03558d46df9d234bde37ceb73285493d2278f2a1a5c5d1d890f3f238429c516c8b82d63748feba528985f0a126ffe7f2b945be6b741372c72296e33af9e36fc01252;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6e681edd26de47c8117cf026c782f5b3561108669591f316e8e4d50e7155a47e1a4959a955474ba75aba46bcbb62796dfdfe7f28fc23c4f13f54c6d723d1ffd0d883bc6f13b913f182d1a594c044b2a704d3b29a10f13e56bd2341a65c2cfdbb4bc2523f1b78c839cb70435f0eff093771d9c8f062241607a52f77975585020a86ccaa844825d5f5565d7f2589782eecd05de3fcf4b544e7521ac052e5603ea06fd2843bafb0a58bc9a6f8b6be5920448aa545871549862f1f6cae99b761c3bfbd5cc69d97646c4be10965b086cbd0dce4060d00282e4466cceefad03519451198d1204e4931fbdf78871ebeb18cecdb2fe07575811e4015c51bda812a513d94aeb73bca2f47ddc7db6077590bf6d114c7d34b47581c31bfd8c5a1ed2376fc397e055e849b5b5cabde7170537d1f185664d4587b5814e647370d055f0d38592f59027e31060cc76e6e5850ff6619236fcc97e073035ad0775117bbd470a398aea2c969ae297ef46ec0367f565366ec20bc5edc98f23f09471936a444576e73d5505af768c8dda4ae03e55369c0f2bab0c10e166af590bfa9426e1935a7afd662a248bd477fbdeff03167e414da479fa6e118fcfa066799834e40da5bae16928bef1dc9b6828b1154f5ac378aa53a5d7ed708f64ef87e12fd164d55d95e533e4bf7b2e789ce436ddf500a2cf489cda0baf66f62bc65809065d93b3aa58423abfd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb8a623cd527431f75a805646eeea20d1d77ab39ffd2d14714f3cd95089acb8add9e5535652fd151f77a41f68c60fca3ceffa0711b421de5cd02dcdf506f86f56d842993e02a456c13cb391d996f1ad017b5d7093d365ab4239e96f08023c466cb18c8b4982ed16bc069bf794a247e7f3f504735ec52ada1828dc3d13ebe0ed20d484fdf60113ca8df552b50cb6345443f1f7a54eb2e74011918b278297a700c9849140296196917dc3f2ff9d7cb1836f5d9646218dffe7a8e1bc2721578ba843669fb4970da67c7442844cfb3e7d9b8c3ebe281c96e19391e4cc09887794b8a7d303a23c4779b65e05f8216f5a321320cf8c2934a4850c1f7eb896716f877a146a0ee84d4276175c74dd064f3bd1e32685aa96310a95b73605e68fce9519b5c2f2565276ea35eeee91630a0e6f977e9a7ea6df8aadec611cfd25c71bd227e1debf3fe0902e465ada4a23f284ff2b45b72ae675c0e8cd4d83909d4c1abd6484e1b81037dabeaea755da52396c271620624011ed1a9306f079b55129006749f07608e2aa1daf50e3028b4ec33261a8b0c6e183b67f609ce5fd672cc47d9cbfe3ab5adac425529b95dcfe0ddefb21c5f064bb766a5f43e882d831c72d1da9a51635f774146637ba35a1e3af1546760a6f2ea4f4f9e6ab210bad9e2a6c9266ef6eecdfc0773c07b15483e1b4a213232cb8338e81f421e58629b5666b94d6570af3b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf258bde5a942fa485fef80b09851f8d011bd25f343231ad26d198eb085fae7421cd600718a7a759d94248552ab6d49805f31639f767d1119814fb1d3515b1976a0276b23db6fbf1c324f30db2fb6cc6d0def001ea6fb6298da6090afdf6b4c9582527a66a6f47b36fcba1c7ab8b360bff4a854f0fdbe6c4897680ff319e059619f41bff46d4576254235afa90ed82dfa08f93a32d006b4949de690c71ef15fefea7829fd1b927a327069a4b727176f0f4b65d1a65ca947b022697d6a85664962b9a11eaeac5203c3f82b3782eaf5aa0029ed3125af72d2d14a4d4307e56ed154264894e9a55c93bb92604fda06d3c04af8303567eb510baf333dd17a2e1f4c6e569d22e8e5ba155f93a90fa980f620eed3cf30993ac1b2183aacaa67266ef34a09d1d93043b5d1f35d6bef1f55086961f28aae73a87c8ba770d22cf23f081bb5ba796ad29afd298ff649c4fcd309002fb66ae5ee471d1547fb59732ad57f04176310ed44ba58e91d5b86f8a3386d77e345ec39b5c05a3c69417920de653c2bec3bad6e86314fbda77bbd7b8387d6dbe7804667d2ec0592649c1b19d5d5193ed323f7f54fd4dd8b8fdc2404c6c3a4a6ae381b49ff6f422a3fe0c2d6138a5e50bb8ed9ff90e83d3da003d10c90dcb48ef4cd3839f82b746299fd2993f16379995f35275364326b802a3067b7c5bb6ad04480dafab0bd346ffc55846710c8091b68;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h473839d57717eb0d0ecd223e10daa7dc7a47791748dedd392547eea25b76e9cebec05b5d46a7d6d002f7b70f021f742ae24de01076a6e6e25580ce316b7fea2637d0aeb4f85cd90c37124cf041a4f768a248eb6f7bc8ad23d24293c8798dfb8f56e9c2559983e8f8ec7f8fb1bc98a1459b9cb087dbc3b0648801dae4b88be8e3d6cbc9238e740705af6be0f573ad4982f8f310272a57f8b8e5400b8b08c83e7047ad1931355bc1d6c4dde23b0303f126ea0fb8f2e157f08d53dcfd3934c030a9fe301b03c8157e4043131c87ad8e0ec13bc3dfb8a265a89254ed936630da1d73ad233553c5efedbf94520dfbad988ed964a9c02e0ce456ec04ca400c43e2f62ffcd6f7a7cef0aab8f5d3e92fb960aaaa2dda8fc2bba282eccd82ba1fe933bc2fc2789e316a62d64ba413a0c7c6f9ecb783044c6ea1a2cc73aed5097a4cf846b8c6fc9ce75c768780273ea774bcb630da10b38c4bdbfa69a3857badeb8a81841982432fb5159c8ad83ac47ed6909d85d9eb2eb55e330792069e8b74c061287a32cd643806762d0449e0529ca9a8b546e6747800f82332b9709f61d571c2ce91c12204412202d2a88c0ebec3a71b20214040e6f74026c50ffdf1ee18cb1cffc56285287d17c864ab4b4f60ca7bc15ac78f39a1aee560a8b2186438d1303bede13e4e8619e285fb7e33eae5ad5ce6254161fe018be141ab4a276482e160a48141cb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3ffc31dda54ef4381366ceb97dab45363bdb3bb0c9c36bff8f98a643d49c8c6d60652c28ed2b1d3c842a13a1967676947c46856157682e8a8f5d387310e4ff7e928bb7118a31925a2fb35853856a96dadf773a8642c6f3e77f90af3216e14495a457bd23de1c2f1a8d30549d7a314b7f592e7e3901ef5efc2da8023970c7e91cc79bd2d639d29b3dc07e83c366a29ba5f686cdc29f595a1d16daf6924996795f9e19372f98ea336727418b0427a627b798543bb60652b81ec2fba6b5352e8836d7ac05defacc7518ead65b1c2655a43deaace4504b84e2928cf22f78e4ed8ed80c8de36ab468a23fbe8a8b3a05f6d839720bf8a566655990286528b227af4a0a34a49f872d4fbebb72431b1f1d79e3283f5fcc2727b763465cfb6df2908cdbf04b942619733b7bef008fa7edfabf0d4c11435734e5e3798fde37c18142c746967a1f0abb1d5c7913f2e5f6dd27e4c9d9fd718088976d6d5605dea3f0d42aa9b76dbfb8b7a9f38087fe957a50802ed7bc5c9608fc6ec19150c6082dfacbc0320a14d41e6351f2fa545c0ad9b638e19401f89a37b3fa52b5c555309088911a052d065d09d34f153fd8de620ef6eb7d0c97f78d9553d70ee06146905a0e85e4b958636c8d9b6aa45c5d0c2077952537f60340b84391fabf76100c42727cc9fd6be36ed454adb9e650c536ea75486d082b9c781dadecd56bd62b32f436c31d4ea358;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd52d37b9148e7be3778ad479561dcab37f238ef2a72cec2a5c3886b2643e3b437323a4b76ca48cc77622ea6713f9665285d9be1b05a8e0ed05f4dacf1a4bbf328669b26b91e4317246f159ed52c885bd28ec48b51cc957bcb2ecc3b26a9bbee64daa96beb9e6fe72528d2015678c071f360b742e77a4737cc7c9d56e7718a74915c3e3328dfd67de98bdffbc0f843008899685678861f4de6d5a86581f40f640f1c9d0be724386ae11e5a2ddd26afa93e0db39f370f6dedb5299ae213f3ca4d90ba411e211bd09679588984930ec34fe4bb9eaaf8b372453171f5a070cb478f6add093b3754dfba7241d7c6e28dfa082b2a6e480e147e38c39eccfa530e38eb13c0e43bf1bedc49eec9db519cd4716681a7d88c0515a6a6b91af595bc2c033a80249b633bfcbbf20d5070a0573773d8f50eee95ea8518f3ae532f0aa5c22e1a2232f6e30b2840ad693e562fcd29e1b74aa5360ea6796f5c6d43da3a36a04ea8d1421d37e107aa28ec12cb0b090038c585d4ef6e060f1062cf58f64b7ff0b8a7fd807842328309f3a4e13e60855f98425461f33080c30c262997f72f9168ef45fe759752a2b1f7db9f4c563b646efad3dccbf798446e934a8f5895561a85d271ab9ca33dcbac72a7d24940e80dea135a271d775b351ecc724c14a94ee639ccea45c597ea88f173c74d074ec40f43a981d8efab8a79162c220b7d7cd05da8c735a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2258f30c089058fb322e4063f79c5715ac2c60ae7588a6cd4122a7c4f2a0bdc5dcd1fd548c0dbcdf431aa5f52b74d9551fab3b1c83cec33ae9e4af164b27b80a2077f44b49c558c89f99c4aeb1dbe29133497331b3b1f46af3936597888323bc43accc79598f9a058e386ad412f6c4c26a37800da546a2a89b9d9ac9d3495794bd1372a9cf157172eee9ef1ea88eab9d57dc3a03068ee3d5c5397dc07f4bc635547c2acfb80071aae91bc1315f0a3dc6821679d510bc1b3495705d96c3f6b8f98aa29a9ea2f64c9ec69f8f58ab5cae758d9121bbbb51ae9566972454e8e3cfe38d7d41b4cb20a6199493f4155b309ed6efc2fc4857cd1659f69e8e8c6cc817154c4f61132d028a10598b11860c1d99fd8680e65c55c50b66f78779acfcc58fdf09ac6d3597dac167921c92e7ed326dac868542b113b9610b4a3659e9c51fec66414e74187e24df3bd0e7f90446fcc6ef61284b28f3268a0837d4289036e89b37a9663593e67f8c795722721e32c7acade2ec36e8d3228aaf41632421fe0c72243ac98381805fbdd2a7bc006e55a347a90202f02ced4c3a590d6944e6ebb033301238602cd86add46e83c105dba24c0dd27907f31a206a2630361d726ce6619ab6adea74c6712492faafcacba00ab06545ded499863d10a99721fe00d5fbb3ea101dcd3adde137edfcf740ced49935871723f7164bd41cb1c38540d32557cd2af;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h789569c9f07b968730d22b806c6e5744a136dee819b9c05b10d0aba59747f183f3c36dcc3f0d858823af02e87f2921d76e27d0f09a1a6f3857156f299316a19ef19242c70ee584f295fcf6646de409ab664097df22ee5c8404ca776b1685bb3f671f3e6f8d861e9108d561f872cf53f9217b6211e5181cb8782e8811659c7208194367c2f7e304576c56ba6e9efa6f7b138ac662ef769eb35144d426753251aa876221e1087b4a11309492b6bc1dc674b6bc6ff93ecc4d1077b2a96a42e85a217bd5dd775183537d80562310f2e67433b4c434b08966014eb8900eefb1f6d8a5b7952d555575747948f8d56f47aaaed8d06a8e2ddf0d85a77a00dfdb630264a463d40904527dbf4c07d12143435a18c1b75cc0b8f6d29c1626a58214536a543de2364fc89927c239276151ccc6baa94188538608d5203230d41907a343d5aa196d66366e265d2b9052a403ee39f6f12a430976da261aa640af2bd6e03d84a585a2e8de738104090a58dbb73a1324faab82ad5a50cc950fa6a75d44150d69f13780a55839f52446a7e55289942e038a52a4ddf30180cbb7a13afac17acfad29708c14bfa00f4ea7c2bdef496b0a387410bf97cbf01620dbc1851514ae46c4b98a8129e0b81be0c414d05f1e287557d3e3b238fb528da77b569f6d5b4ef374e62ae48ab776f325edd0a31fff59b20fc11b242c5b57aa4a2948b28d870ed32fdc9c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h478984690f21d41ac1c0d721f6a36ff758ed13444790e286f1419795d92a77e1a21280422c9fdd1b269bf5e6a1038a2d6ffa38d2bba58f09a3e1012122a77fa807f8bb4bec91bcfad521fe89952ff0ab83bf90f569913e9b1f10e508e22e33122d778f1217395a6e8e7e7cb79b35b186e5cf3dfe7a0780460a6715be70e68739b72cf64ac3af6b56b8de57137ea834dc51e29b9ff21924845316e07a70db30ba960403ea75c0b054c28ed283adffca90434bcdd5f8a8ae33ec22cf11fb74d58db06beeae29284fcb68bde0922398894e4dda7445e3bfeb9c8f7adb571c2023ce02075a0d6c326f227d441f7d5641d5ff532197bb0a31cff32fc312597a67de1482607cb3d5a4b894f0f706aa299f0a91ba14f1619ef3ca962f23b962268b40657c2124d82b59e677296e4478eb931561fa45432ab8530ee9b142ca8cb2016651ba2de9d9dfdbc4fc20b9b106e1b3a6323252a7652df9274241483a8dbf35fd90330a1ec2a8f4f903111cf7de4045a807f430cf45058c26b0e986ca0815507c1ebb0a3a86958a26450e5d32f028553d149612d3597fb30e6ae9708c40e0669158e3dc08e0133585ba46a03fc4c5ae6357be8d167af1171e7f31d4c0c7b9aeeeda5c73f0c93f07c3ca6820909e096e2d1831bb7036f5012095c74a2dc0ba99023371ef8f8625758886a21b79d72a2c8c8f62e706d963ce4effed58c8b163da5688;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h3fe789fdfba027c39dcbac5ec54eb6aa928d8b2674cfb64f99ad26c99172c769cd38839d3122e9c5d274bd3201d2fc8bfcd216e1c70cec1f49bc25d766b3863f1b660c052b1c1ef890b56e1a5e7a621852f01756591d84c5fa9ac5eb2f98855d0397a4f04b82e3373e9a95db19406aecc8c6314157445b891df7cde8bd50e3deb6c35e0af16758cdfa6552db1d120a3061bacee2598d20b2fe7fc4b4093f46cacef81293998833ca065d1e2054f59164495bfb327542d0ca5c272dd2d3cbf99d77fcf72a429994da3bd62a07d21095815ba54f4b786e0e10807104d1cd4fe6a4bc4dd2ac407d1d9d917bd9825b396c12a0d2160852ea2af6027067923aab857f1c7ef8610611a84390cd22d58930f08bdb3c51a30647c0a76e16554b6d62735689819ac6d9d3cffa935c2523fb35162022b08bf5e9cd3e06376a606886c2cadbd6643755ebedd1f6adbcb65b8507310087e2fe32f29494ecfd55d27d5ff26f0649f9f1fd98f58d267b374dcee4b0901972c92b19239e7b70bf400b8ac3917ad036fd1516f02eeac4b0f3387f23d54f18d2d68fff7e51a0fc4f0beeba2bc40334e7472b79faa3243853d964a962674e71384917bf4634f5a20f57b6c39e1197ead40deae340178f5815476e9abaea692f08901f8f9a7ff1445ca906a45b02924490d281786a93b32bf09a03c52ee5680b7d47d1c970f5329a20d93a9844510155;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h841dfec2d92473a783e4c4d78cbb5e734b88420edb833695b5b667b333c47bf703226f056ee986f56d55832793bd7bca28bacf839f6c10d6e724bfac89c2e62be1c6c17676e16603304964d444ad8f2fe5d1e9119523dea2c12f59035c335365242f289cd3455e9a71f56b3e0ee5ec404546cc70e8afc6d51e7f92f93a9821c37cc72bf3667af70bac89da86d10dc5d14b1bd2d33e87b48c49eeb87bd7ce3429d06b4382a7ad2b18cbd577a93561e3b7fdaa4ef36e8a02fc053f3c875d43a71fa94408eb14b79313f6ae050b3c9aa68011ab224bea7aed38ae8302c60f882b36b64cb161127ba3a0a87302e4757d75691af81fbe8e1981920279253f0f4e9f0782cdfb75e24780fefdaab9fdfee2db12145cc4b9a646982c00faa8604cbf2f95f9df84a59678ad6f3052795482db0dd187d2a61c53109bb957258265c9f7aee16b520ec43ddc600ee5f5b709c24cbef5489f254812da06a509004acffa2a70ae46d94a236214e954029b0b7e930bd833d7e4bea995f8dd20f1794bb5eb8ec589db82f82d7051e0ba91c1d10e17f131aaffe47b287b0e2ab904e44a1b38e0ac785c12a532dbbb922ce55767e1505e228c14a04e27d5a04cfb73d7fc08eecb5f936c387b2619e8bf15720c647d5e38da8c5edc9df760a288ad2fb8a6a3dba6bb4bff976d12f17d76e6325a309f0e4164953015e508e261b91feeb38d7eb780190a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6932683ac8504aa63818882d6e3ef809ec295ed341c20bb4d76f3cced3859c9e8e4de361d295b7ff7fae04494acd5d07a48788f30d6658bd9ea6ff1802942a6d134a2ae114ca2c29fde9c29887450aeaa8f5772378afa38f6566ef9285bd5c1557c54d2b79468b677bb0edc9115e40490f3cb6ef4549341133e564b66aa39321c81db8e0b1fed9fab2e18ccef5160b84a46ceb4035da19cec9511733441287e92172fc0c11cd5c8e2faf75a09f1d9cf589d5d3e1060c772b9497269d33dbc3986166b3d67e7ae015f2eb6d5dc7f0eef1efe79b510e111d52a8dbf3b45f42667dc3dade99dd08b3d76381228c57b4d4bbd787cd3b8da38bb460bb9b561ea1b160c696c54b337fba919a21523a710b5e2ab74a7af45c82244130c3b787f85ea3d3c0149898ec8860f04d03e683e2dc8412d7d101365c22eb67e3ec607b8794a58fcf731db6b6370716cf0aeefbeec2d7012c08338d74984f44a56dd174a1c0e759db0ab790934be72741d8c47882efe3f86458ef515f97666c14b0c794ad5e404ec63629df3a8acc56bf93cdde6e509f4059d946a4ae013303d33654be1fa90c6b85bc2fe94c3391078fb8a0d3ed730ddf02a5f1d4377154f956050001244cd93adba2b5acef96e2fc3babbe694108e1276800f910225accc29295e2c771f6b687865b3696e31ab9ea3c40a05d6a4be603defaf33af36d1b015910b492f0f3bc0a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc94486724f812938d22a4eb4a39c96636076f98f4d2a3edc1b98f6a70c4c4e8691ca6dccca0b6504a6923941d7d76743638561c4e708e1f482d046e12a3c823ebd49a11098385bf23209c8b95d04c4130601ee5d2eb9f6273026c4c6d9ac489de4d3a92c29ca3e932030988a627b364e9fa020070588fb1a1cd2aab8f071f842560b762c66c50ded514c289cf89ea753fb1d7842430c7f6cf66f0722e2fe3dc918a87f3c3f6d4401ee3fbeaf553c09e999ce682a3dab58da9094b4f872562727d659e36635a51f69c1e6ea4b5e42a94557dbe9c85ffc97d030a89705f0f6929860c686e84d7e7d5e6f3316af2ee234c13cbbc41bad62848557bbbd08acc727341d2015cac66b834fa2fdd65dcc833b0cdf7b323faedc87a4cfe190f295f3db3f164b9ac6b43456eabcda5c461974e60f3efc14621fe340446cff6bf0fd265301d46168f9156e09efae5b6d391bcaacb27581dd4074edf1bc1247cf0fde7a978bd93c1b88016465d709a41eb9ac472e317b197dc7b7731f4b0683d6004580046bf6ca822af4fb5257bbe8fc934596adf91aab602e31bd8a0892da68abbac2986ec4ffdb9e2e67262abf1eec277a5e4eb2c8e3d9880f17af2637dac560120f681e705fb83e7b576a46a1974e59a5196ffbc15338dc7275010ea1829d6daef00aa07acb81df62687740bc0a74b45e928370691c26d33d58cfd97cb96c364417d0f8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5bdb390cd8493ce47665cfb4dd0ed566761066429190b622e557d30c4efeea6f0d1bcccb868efcd8c8c4105bda156da118fb5fd1adc33a6d7b9ebb6f02d5bf9a31ecac33a5ed6873ca24f1446edded6d187d96dfe941c94510b29115feb5ec519e85675d94380bbf303f830c722b9b6ca997bc2ff4cb4809246344637219bc0ddcda76e411eeb19632da33de4837832fe28849a483d153b06625e69e01a71671ce2775dfd7ee51db165096e6e164c7be19a995a196ee27c0525285d3f6a2c80486457af56afd8d8dcf9bf7e615b8fe5f96d78288e1274f8b52ab5223627dd80584030daeab7684336d7b50450ab4b9a651efe1f295dbeac0eb36a5b32192adc28fc989a85bd65311fbbac728548a688cb0c808d60b4a512b3d81ae1310198fa9ef1a539d6ad927e7dbb2b48f19acbb5d852debaae07a7070624fecbdf863f57385a09a01dffa8d6fb79fc25c0751a251f8c1a570a4ee85bf7cdb6fe14fb33b594b83b02f8b6581548a84ec76aaba7d1facd271ccb73645c6b2e2668c356d5b7a67ccf57e78148b8a259f00d33d2ac2c4f206694649a43c06ed29a337d5eefd4645131d110c2b8d0cd7c4d8b5cb5f059c286e4c50e8c4928ccc186cf73faadcc7c0844e99d76848d4ef27d4dbcd6212b776abe19c0e80398ccb8cb3cb77dcbe60e6f8262e4ffd13e357d15a8f7311109f3f5c36d6ebcc859aba064c7d2640b5fa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb51ae765dd6f73e29ead2ec531f7bd88df3222c39627ffc518a9c56f1d1c0ee4d7a7ede7667933d4880f1b2c486c2b991fc83ea13b342fdf251a0b3744682564f2fb96dcd73be84be6c7712a006810d0f6db79f6e6d280c651f7f7031cdb257ca0d818edba145a0c72b34b8604fdb64047826d8c145d5ff86b6e6d881c1405f7ed34236caaf130fddef6515648b2431c3a14e0d715211cbfa94e8f504a140e7f0bd99c052a6ae57652f0e1ad61374295d01bde13c2b5a7b451408fe9eb6e2ecb378f15cbea937856b3fb8c9e9619660946dba29068defea98eaa7c142c5ea2630e188fe96e9c4d7855c1682cc165eed2b85d14aa1722eb09f55ff73125ff90839798638cbb3ce38340e2d8c13292585864f93cb5a2f5f98d1eeb3b73c8b927b6b3b8f685934f3687339e819634c7b0c3e89232981d735fd631d39cc5a86973cb042b64384eebb6070af8ce4ea6dcfe39264db95ad5a3a6c2fb1735c22b884732ff85dbce24419df106808ee042bf174f388e689bb1eea77bc59ffe081b139f2e6dd4cd3744ca45a5c191f8af055bb5bd19b259242bbbfff3e3c42bd84ff650c1b0d69738312d0fd268d9ff6a468970c6b61a8f57bfa2f97a6c1c85ab2cc3d8d1a115b621d98c4e07356f13e2267b5680020ce0a0f06aa874058605d60b03966eb02aff6893a33491e6739598482a28ef72040965020eb647a37ee3a2613be4a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h10c6a7dc6492018d4a6ab9bcd45ba36177e56b751ed9d6944d4ccd06c889e8b5cf81ea02da722fd47a36034f0772df4de30fade5f9a121fc39f1886e4874abaa074e6220b839acbc222511e5d94edd64ecd52ca026d41ac298dfffc597bf7a7a1777c9c52674bc7a638ddd0d69ff2d07fed4cb8a0c41a75ba7ad8fe2aec3b8478c4ddad55f0ddf4823270e8b4e2b16beafcb580df2d60fe4fc622bd3f00c197cbb6965993bc9ba67d57ce92e2f5957ea6540e0efccd3c233db4d88adda0847f24dbfccc289a7b9b3f187b342ab8a97cdf738ac1d7feb2fda46dd2fb2ebe035230321ee008ccd8ee84fad920353a87683dbf1e7e07c7b7618ab8bb79daa739f5abcfc9696a6ee78c4ea776c19238dc7f701be1c4144a02b9baf9a4c2e4339594509758e8972f44b1b2f32c855cf082832ac466add59d2260d88ba934193c8425d20df3f24beafdf84ef763c691575c1023e8c4c5498813e18d67a62d5e1c9b3ff60bbe3940b0eeb08449da93252f0317ed77c6c95644f100a057d228b608f7deedb01c86d25e06a864390657b88de4b54f008df3ea06721c3335a112c6a54c58f5cc9fac684146ba25540e4828430d465bda226249b5f3d534ae4023c619bd87df3721b14c4440210e38d1893279187853741b2bf3f065a2a2758cb5eaf3fcc506bcf906e5be879e5dab0bb6e74022b4b2c83a2137be93bb0f30f117a6061fa5;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h776ceb30b704a27f2e820f138f130d0f6753d0f2249b77acb58e7fc73750d26254bef83d0eb289624299a2ccda9bd885de614c0e64f4a40d67e56eb062de9c85831123b808ddb06afd7d8f82f37fa83694624744277b7e5acbb646165b3f15229053b8f36b903c9a805cf82b1fa5b7e364487fbd22148081d64d11c1b5c19c102058f895930db0334073ec952a62da209ec6bbc48a976c0d040b4cacb89687fd292981eb50a4866e22f11ef1eaa4d4558730ca0b76b506a74e86c6c4f0d3a9ac64aae4c536f8048abbb73a527fc3592eca6bd6353447a7ea878bf6b32ae9cb025f9cad5568cdd89731434109037d00eb9a89b30f912b9c2c6eb77ea30d31b711af95f15a03516de0303fc3e4757f829fd3ca59856b88daa3770b1c6b505a489748366d1768d1371e34816502263d275273eca3a30e796b9b5361abba8711b3996edb5126e49ff69f6975f78ed5300a7813d33ce545cff1492b08a4e7e7bbddb5024fa2a1372a83185938b9f406332a47bdd11a7fb8d3b12d4267041c306c0fa225775395670998d39427a73c0646f85139652a82e33f50ecdf3700832c9340ca0963c6c8419615f4af651d44f6f65d832e0eb02803e5da12bc37bf1e6d79814788a1da782e568370865fbf15009af186dc7e3ece55587b049d77ccb24da453aae9c4f61f16d35161fefff05f9ac078376052fcc5e7fdb337573253d71f75fcfa;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc23af1cf903429bb8ca6f2b308ae8653bb93f8c024c79f085ab9c68621111a9da502e996f781ea9fe3f814e82c46d41fb5126bcfdcc11f53e0af6ec633058826719089c894de37119444545df47af78128a2bc32b36b63e9e488adb27ba0b958061121af11f784c6dcbb1442d4adc6efcb240917dc16cb382c1044320820f02c09b6532af7c960b26bcb2e84299bf650cfe95e2c4e621fb12503e6584125a1e4918bb5d9a4b8800b3a1c565936b5ea9c6c435042b720b4a4cd3095d7cc9e436d8f1d7c990fc97ddc6e3fb4ca4354926d82c20eeeec66a287cee75e36588c46d23d7dd6298aa2e615acd452aed4aeb3ff8313a51684697930ee14ad8e3ec59d32e3adc769dedc076f541efa621d7b66ab91ec64eb860b3719ff6dd3823ae703f8f9a3ac86d72ffd98f4a0f0e55c344d1874b27f594d47855c61071310a7bb7699df091bcc474f0c975af8e32edbe43c907b4198e24ec3f21662c3ed7220539bec84ec6b453c1508d9bc0745e5ccbf76a1fc0769613ad2d045e9b515f42d4e302a4516c2a7dba957a15c57cad9ad9a025af51c0083e26f51187338a925ab3aac1da8d8f33c66ba7fa13556c849e36345bc52770ff75a68b1df2cb0906a144e96ee1942fe4140e52c2296b5e46cbb4b657a0ed550d8d8dae4a5323440b3b0c2276c89d690a912e094be1cf7ad001ba4cb346eec954aa9d45eaaaaa04c76d5bfb521;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h91217ab31d2c053a41d6179a0180cef6d8bf11db135eba448839f141b82676c7282eb2def7572d5be55b4821559bf143a276ba0b3ea11f1915036efabb999740a76887300f19c01ed3705c5111b744a80f1046b3fe69801e376647158adba2c66be43237d9d8c6bdbaca0b3648e995978e8b5c2609bb55025328f40f93ae8ea268e6cdfaf7f2967c99fdf133db5a77e59fd6fcfc4b6de0d0a3dd0fcc74488793da1dfcb64e7876a658de4f48ff79a12685ba357314b2b3fa35655d9f2c9b90eadbc5c68724800dabcbdc62178300eea78a621d4fddf5f819793e423f4510f6bcfd57939bffe18acf64f06ec3a14b8f59d7e3119184fdd992d8fb4a764b5e8427a368460fd08cac16fc18e9078ad4563c899ec2de4bba5564bd6fc46e10ef6c902cfc0f21f005c9196f0bb6e856778f5db2f029d5ed5bb99acd72f442cd4b57594302441de6c62a7f787e2501325401ccb1593b42e4195d49f04128d26dcc9cf6a0b89e6287c6053c3d0121ab35cda812123fa40d0b3a4bcc8c75f15c3409527b6b76daa534cd938202247a9fa9a314470c53758e3412c82d362c493cb731bfbde7f9e8ce035dbc672b21d68ca1ca36227ea37c8d2185b90639e60be4b269e883878616be0197d72ea4b03f963c43a9b6cf2e858d4aeae6508c798b646ecd447b724d552a3c4e63de7a0a0813888caa9244be383fa2463f04eb11825854cc261b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h160e9827f952d54e935e70af33b600aeea11bfc488a13d58e44a87a6a51f2557fcb1fbf58aa1ec0e7e8dc44657575a645f0842f1f61f95f06608b217acc4d16db8eade674533ecd2752e51eb62403fdce84f43ce3d98d3ad9fa113878cd6a6dc3db342147c0bb747e726c13b502576083f7005322429a0eee64f2138d7c9a19826d47d9445c59ca5b94f85956247be4bcabaac0e73b434130df682154f1c4c1c85d18f522e6c1bb59e6597f5e2a6cab5dcdce7c77f66e5b94fdb2a8d05a70b0286d9908c9bad51ebdd64c6d9e31dcaaac8983cf8a4176faa4ce250294c64cac192794440147d2c30db98387774cddb1134d07730b366fb212a7d1ad874b115a82a9790cb54e2e8554b13f092a668799c24f94ce47f94c477a5fca82a13e2e831277be1379532f890c8327e3a4fa0369a9deb77bff8e6f3c3f11deb95a19cac0d882db03737110cab6e9104de74eb837e0141b15ccaf8e058731ed6c11cd9c7721b925d2d96666a5fe459b24faa66cb44d4f827e64c1be97a545ee3e54c969fa6859ee33c943ba31fbb6282a84a5076e0544718325fc0e583b7acf54e245396b3b7f5b8acf0586f1a0f3b3a05b2b9df1060ce3b7bc15228a99afdc8ff1d15b5b0547b68fdcf9b88bfb586cd2db43e6813a4813315349c81a75860bb5b1327b7ece96c02ef6a7c04c42df6f247bf6223a680c5b83fbd010d68fd76be4e61909c5f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8c2c46b3d5405fdbdc994b9573d0136fe8ddb2f71207b7aa0c14789b1363f390f228ffdf51e7c2757cc7fb5e52bcfc3b42441644c8f804b81519c2187d4882ec0cb293239eb6de8d8f16579d637e9c3a9d8edd8a76673c360c46fe0c5611608431fe2c41b1997e248db55971b9d6eb01471a70c12c34121aee0aa3b3eb132709f59f2c9df00e15eb1af9ebad1b1a588aadb827cb4af21a404b68bc8bcb175fcaa1fb841fcfb122140c2eb8a3e292b422646eb2abae50aabfc95ee66dd5c0824e40c51b5fe6b80c88415238febabc388623a1083eeb47000f0b560e8f3d1ad9284667b3a08d6f200d24ed98b4c5b7b5f4db1b076f8bbb53bd6eaf35ff9389cef3e5938b0b45148c9846ada1b116f21e4af2b1992a51421bce720ea96413a2784e1bdcc52dfd600b7ba8dfb66068c1f22b4a3a535f501f70f99e520d639b01b9a80f9c7f618689d26186ca8cf5ce04a8c31618746e5b8b565a58846e98100584a3654da296e2677795b8998d65430abb2600faefb6c38d6f02d4c9867cd0198a3a3c5875cc060ddfc81a97ab1f7984149e91af9209d3750d930bb7288877d8c64aa37dc30f637c5dc88124a0596f5087ee6afa121372cf6e51006a5cae99aa5110ba66b12542573d8551c7aa1833a668c5917246d6edef9b0c5c1054b9c0b3934ca8f1445ebfdc8dcb7f78d55d19f252ff01e64b4e452494a140176379fd7538ab;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1db5396edc565f417032601f5ce3df0e97bb83ab9386caccb46d810831865c1b099fda0ce9ba2398d8866e087d1390216c8983dc8673b2b5d7e5a1848e0387d40842c7e7080ee8c6a3cc6560a6c6e417e52ded3f19cf4766b169301f7207d9f7fb25bfb697befe13377d3675dc3bd4fe6cd8e7f34ce9123d40c63098334304976edb528431cdb085c349c1aba26f788f2b9ee964a50f673221426d0e5d97b9a9ebb03881559809fb02874ada8070f57a71038d4420c0e22a8a3c59dadd10995bfee6bc955c3d3e6edd731966c9cf8b8ee318b806a1c965a3a9dba5d09522812abadc3c3527fc6f84cac57ee272075615ae74efb41b9a85275b4fbe846c045bac84b1216eac7e7abd872f3a95a4fd77942cf847da16a9566c0760300e13707231783412ced6ebd7a7425294573c1784872370d0e4ae41f95d0093db32fa74742d9a7f95e69a1793630f48bd2d084777ace68460ab395ab5ea6fec9230ef7e2b2553e3197634762773038530dbf157a69ea232d498ef85ba8f138e76cd2f8ad4812016d4655eae18effbfb8d4e3608835b9506c885d1519b26d5a8d1de043409caa41a3d21932e622adb6b2b200e24cd3ab0bcaf76be3abca845ef887fbfddb0aabfcfc8a3981c7ebe8d8decf748c916d448ec17081cda94a40e91a3964d74bd484058a71826461a3f480147dce4a89381a35f32d048d57f16d3d5d7cf3322e68c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hde3dc6a2c3deb338ff8153d5ba5457f4eca1b8a1c007cf517fbfd94054e861e6d82910e6db7de9a9d5be5bcd3507f2f9c716217168f72ad1409b7e2134f230046d132b18d662ac6c2ef1e1320e4474bd1d5e591ed401b0ae7dcc8faff4191fa537a5bb4075a18122ba7fa638591c7d9592f860979fbc9aea1eb2905f3d02f07f6b29400b41f095ed8624d6ed641828c9b48abdaf0243711d361d40bd75ed9d44169ec4d7c08e66553cc93c1850b2c32aadf537b61bfb39b15844f66cb7f98cf0efc9539d80cbe526eb64ea4500c5eec3e490b21bbfaea63ac63008e27c49aff6b70ae7b97af5bc6e7ae0bca3632e0ae7cbced558c37aeb6e9c1a00f83176302a0a9fb569995fb83aacee80b432a6ae86b256a5ec7125b0783b9682c378d7af5dc29c436d2a86b6273d169ffab714e3852f1ca3c7524287c0972678f7471933fa911f5d3e56595097501d7045813bdf14e775b0efb88510abc0ea974020f8a806d13d1ffdf27f2845229ec01f76b96fde651ed3141a842bb67905c325e365a2ef09957505a89dfdad35726b57dcd764bac6f5a2cdaec737c64abbfa6e18ec4f82fd091e2fea02c40162745ec501f888d0187da7b5bf2ef153336b583f401814e3a65c40fe8c944102bb39c8da99ce7d4879e2624afb562b66a953e422afa6390709b382903aa3ebcfd6a5b895bedea1bc356d48067e3bcb86c54fd42b5d771e14;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hcdcf023032bcc7960e7be0fb8eb23538d255d02804f71307b10c18278f6ddc84bc7d9f65b637c88514135d98762a75bc48cdb3c4fe301536cc4da9126e63ab5261464569297015ed2dc20d1a96a950e852b41deaa6efc1c51f1e0cae0c71d3fecb00d82ca550e452f18e5817e15f88436a2aa7bd0de174dca364ca014960131464dcba94556b38034c7b184bbfb6b36be07f601d50094e07cab9de5a80e1198a3ead38711e27d1db4ed12cac43cc845393607976c6f55f4072ae70290cd67f632d548cd7a80d8d63811569e95768a8e56f743a9004dc179d4aabf6e83290e12f09339eb098fcf6fa255b30fd3b811e12c2fc8799188ef1cdcc9b00584ca87badcc48ba30e7dbaf4c84599d93cbc6f9277fcbe2578e50859c86be535476a54cd7055cf456a35694b3314ab9967bc8f250beadd71c4f481a30a6977ae67f039d8e509d6108ad2cc37d9bea4f936a9e834728861093793140a21c8596fd1bceda968ec69947d0dcdd5649993ef8dab54582515c94a55b7da95bd9ae63ab26593b05d879491e47b60f37e9541056388518739c6f7c669855553ed8dd5f19db2893281cea170d31a540c22aac1494b38eadce37a23a70a55ecfd96cd1dd268adf77481ebcc6619b56b4d8cc27843957e76e0a1cc0e1e2b150a2c819a3ca360987d00a80ebb0091cb7fae1ba6077e2bccb1e016cc5362de6fa9e0730ad87e9b0edb710;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he6ae7337f8e5da5608188354776469008a2069f2208051a7734ea3c9b596cba3e0efe52583661f3ed8aa79cc30ffa5419b2db45e79f2afd2fde699d4fd9c8a2a074417ba01608aaed94065b79305aa686b1960e80b2aeb0d8168d5e04a5c193ff47e245347c2829a4cf5d527beeaf5a57680763adb323a968bfe26c7e86ffd0a6568818a5247a8c0e83b055924b85f3b88b3014059f71ca60119a1a325eabb28d2777d3496eb5a2d50883eff3e8b422edf9dcb581a0da9e38c72f1d86c526cbe34f9dc1223b2c8c4bf90e5206b36043e94d202f3053240d73761538e45c7f8e2236abfd28127ac0237cb74e4ea1f20a48d3d21da9d902c4c4aad1ae98bba7ab633afee8dd8649e099d60954601782a7e55687cebf132bce35a43309ad03554ba4650993a363db4208de3bceb1fa27c7df0d30150497d7f924741b54714bfb00a02659a95495ced584e5c6ac60b8710dd0c5f1db25aaa92f949e6cbaadfcf2e5fe7bb24829309e6325758e02c46498cb17b904306c1961ed62c9ef249dffcae25afa01427fb583a05d5792b76a48505cd1cae4565a72f84fc321200bc3ed24ba816c7f053a0cf488210deac69db9211449ce858941cf9af63b798581c487d77007b4f752e4346e0928125a808bc450ca44da84fe9a26bde553ad93d64b1e49a585366f128266cd23391942285ba1b934cc67a0fb5f8efd9226845ea20752e234b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8f5ae401bab70e22d8963b160107739e3ad6cc14b6e343da01175c4b99cca4cede5bd189a7ec3f6e6a654341f61e1b842000da74c4c0eb5dca958b88ae4ba55e8294c5e389cb8359c82ec44c93b0cac85742b73ab191d87492501ad1b0caa874a1d036550b264ebaea5794cb7fa2c32a499e1a998fb0e06234309383b447dd813e8abf8adde5116c19d002a53b93d88e1178b1bb8aac4f52dbaf2fc20b508c868c1c1967d1f6e0cf81fbf72cd94f45ae66ec7d84518148894def9a14fb91b2be46007758c8dfd1a056e33f36a5ba24433f10ebf97c53ab6b1c491cc209843cdb3623a081a246d6b6858aaeb129a41e13a253aab77db8db56f7eac3ad38cf27a0d2ab304cc63c26ef0090e41b562bef4d9d2f2d02facb02b241209389fb751ebe373eac957f8567f8825b1b1bba319dbe781e36972b1b933f0d0bc6fe573b7487c5c5de88e2c309ae7832277dedb1b2cf72a19e515f369874bf365052b19b9965e19ea7b71443cd381f3232f2bdc527d155460061872beb73e8ce5ba3bb3a90a26d962a0ea2d9a25e7930f17aabc2b388f330eb60190db9d76f7365df11335bc8acc874dc6c7b2cb4f893b93b1e5df6578d14457e22b340571d4065e156b5291791eb4b33640458e0fbdd4eca2824f17015e77a0a5537f0334354793a706758f85e79de065280517bb2773d6de1da945f520a021271d471f11e9a1a9810cbe681;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h58966829124dd70edfee3b5f39761e3db2d2e9711ee61ff1ba007b6ce53645e3e1eadd133f7cb70849f6e28f16e581c7bf85e7774bc9c55c9634adc93dea933e8e42db4c5fca4781dcb8c14380f70d960403d01ebb60026ee686d5ea48d35cc3dd00f694c0777a927a6657d7c2ba01d5b736ed043cc3120f829d14345e3b498514ed72dd5f991c6e02f77e2bfa06757ebe531d5ebc05b7f76dad4bc17bbb4e64250e24670dcb961a560129b0b0484e00dd46bd421ea1268ad8887b066e87b3ca977058102840ad8af024dba52830e96547c58f9e0c053f8ed11c559a444ec4130c8cb522b399601880d31739e68e9a20d6484d2f9a25e641bd0ab2eb3b1f7318d0c92e395b8f896aeff73aa6f958f145919616997afd6f431334b9cfe1789a2ad5cc01c63132f7a65942bf928b96a33fbeecb1f3c338ec906b6a258df2a62fea1a5226d33946e39d4e910873115126cc0f1e7cd966272a5be373ff72815e9c45210b3fda39eb0a2709649187cd1778973d51f03b3a42d7d8a0110b471aa9837d227b1075083590cda3be641ad95ffb08065d3c81f04d09fd3796f8cfbd58f2756acffacca23efd6d48d6ec9c218ac127084d7c7d01902a900bfe1e6f8afa6b381908138587db0bf441682bf97eaee9c2133c227f61c39c9a7a4fdeeb1d4c58b81c2e7b782fae870d76c444cfe8424af280e3d8e01db9995df9503b2c86ea90a2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6b156d519f1cce3af0b360908968e2b8f96d508060c546900464aec83277118e6c75f7ae6ccba9ebd66206a5e78bd8621291bdf7b2ae0cefd75dbc09be9019bf9791ebff61663898df0c2497f00513f3dc1252688ba7e464d9c9a963ea1c27e63a513db38c34bfc0748f59a2c11201c6d49f4a91b69605ea912ed21732402ee614b33f531b9a31b3d6c7a15a805621d536d3911f49270e70f12706dbe8dc911c6881a28e96b55626496ba1d3276d876594d6e1a35b4a73fbd829327908788cae0c94d83874367fc9fa323ec11ca9afc9cc3fb3be0e47ec7e4e2122a02d73585cc27f9ae763ddad40e059e4ea0108f1318f0f8cf9322e9c5f25814d9b70072caa9f10e5b2a67c5deb1f1c8037cc7ae4ddfa6d1c1539a12503d4d3e84916d8e51e1ea8f7a6a5a9b3495435f49c4fccef3949cfeaacd135df5c79215c2d8cce7a12de4f7cf9a0667e186466471082915806e1609bbf33a297db4348063f8c6fd50247af559fa782262fd9451245f6569b78c85c508c8f191b46d6bc946df9257cfe8b527fd4731e551c5344b991d3b661a3bb6bcbcc242feee37c8e2e3657aa76dcd5bacf578aa7126abea709475c105bab2a14eec82566639cee24831612e5d073ec4173459263df3ec67f33114d90c252a9ae8fc3f421ab9dcf084a81d06271d87410d0c4340227e01c564d209315d04f3c2ff48040e920184ec353f9e5f60c78;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7a7d9feb2b08f4deeb18ec9f6c78c85c88961f4b7eb8e69a6b0f43711e77029d27e600d752756c3e2d2eb4502a8f2fb150e843dcf70673e3f20fd16083fb893739f50d5c6ac104ef432780287565cbaedaf2ef7468c8ce5192123565349c024ecc2e2f5f770abf4535897aaa424d9a6820f25dc5ee522dd7f662be428757a96b0efc17206496a7c1351d8bb28fb589135d96b0d694b5067245bd9b204e98218b57388eee0a54fae0ba85d16d091b2d5d974789da1b9de34ddeeb339f0cc625e0815a116b75f5b57b4d8c6c8ef393c3bd6c2e599e79f5e232f21331b639bd6754d7d736f3437f628554b08b5a3a4f202cdd665ff8131f3ac00353ecd137adc0a68222dfbee66367224939c3a2215d302e5bc915116b3a3815fd3bc6279dca8e5cee9bbd48702358b2fe03b669ae93373760baa78cf4df1a9e23a2841d123ca5663182c44bcd03c4ec17f9185c2b0f571fde880bd4715f6343026d6fd581b381fa9756da74f2a12a7dc68e791674b3d5a6f92dfb7a8032f9bb1b3f153a4b62a0675004372c524b376deaedc68f48bdfb5b3c643d35a72164231286106600184607db9cd717c99a5d6fb289b4d4f22ef00e2aff3a171270cdc218b4a9ef27887ebd81fdd4c9d2fbec21fc5fccfff1ccf914f8353bf2e0a949d04cf8d136bbf2f9858397ccdd6f95e24f0d15a5e1406449c2f1acf889e6a01397c324bfb851818cd7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd041ec1fbadf0902e742a76996316a380e84bfbbce20e6c0d8f1fdd329c960b9ce7aa2595b9754219c540d240f3672ca885fee52c47f507f50faec1b2b57bbe735e83c85b1bfbd9413ab2ebcba18b9c58e9dc48dcbd299e2f910c09f69da40bbd5c8a54c137bd79f821d2568d9aec2fefe8e2b50d958d482d5ce92dc750b8453bfa4a52b08ca91e2c44e4a38164039dcc2d6ada7838c93d547d9d73b686ac65d12fe20b6a1527c36b717636115aab08a924b1431a913b157e682603ada7bbfd0573ea99067c12419f3c5385d0062fc37f6ea87f761e8d069781ab19059e1b18f6a36bff69c12202cd9ee7a1503f7f7580a37ad0701e16bbe2b4477b8ebd6d76f573ce7e65b63afbb1213e9b1ddbbca09cc6a7bf53c083b5cbdfd159cd21d7a8c004b1c485f0cf1f7fc88dc21a3b72ad1d58d005dd4550df93e5fe07ae36e4bb4a74987e3c7f39f21e1658954103beeb8a6416b6216f898192a401f10bf63deadc97aaab5b0c25c2e09089c3aa3e4ad2d294672e1d13f801e25c8bd39938c3e04e765d3eb850a6b025665c44f097d9074773c722fa34940229b3772d6f920b3e6bf05b176322111b082f5e1541e9d995ca0c5c8e76f3948772a76144ee03f734a443ba4e1d4ccb7eeadc29668403e903957ce9fcfbb8aed372380c7f63db055a9ef212bbd918c17f1bf6c8513752d86c76b7f6beb8e374c63b919cda546bfba23;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hcc57ab7369605eef478681a291977a6930eb7db4ab1d5067b1a4dbc4a45309f4a8da5be54f0106cc0112d224f7a0550545319c1ac9268c8d3af6138560d24d9a1b4bcf78518b04d3328cde2df36aa204fd60791760587bb1c9b4e070c3d78b39d2938e4aaef9a34029fac5fb326e95949ca8a5a2f1b38d3815737b489b433dcc18f27a3299a6bfc7d8a78464810b15eedc21b8b4b1f8190f2185d427589e929c964eba74eb1fcbcb93b2ee7d7f89e99e05fc5bccd1a690f5870acacd4d1524bd7be48d360b05510f7284a5909e5d52f9376b3e6670ab1dd0a9ec18d4fdfc9b9ea644691b02d55cf0953d127fcbcab21cf9bc005b79539ef7d09d88211d25d672bb00dcf2a05c3ea9dc0e1db121d9c21bfa7b6de6d15a1423f5e3490be0d51852893ed2096bdc7cb739bb858dca7010181aa9a2b3fd94b186b8305ccfe8ffc0fc70cf98b5388998e8366bd1e0223fcb7d66044a75002211a4cb925a88364dd15a60c9c2618d2e03e5f1210cfff25b18c7b9a5d6eaf838c98de700053735a2ceb9f356b0bac92f2abe7ffdac71b04e025905ffdbd378f0eb774f6354e33b98e24ecb9f74253a3d72bb689afecf209340eddad96c5a3ec5c986b9456f7b376b93f7da476d425d37affcefa4f4fc5bc72be8fd2667e0bbdf7f25ac7e3b559391219ed0057e9d084038fda8e2ad74034b5e83af40c57a399f4ee7997276624322a3fb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd881df5728b2e761a716b09f571eee6f1b579fa01d7469b953166205826c72ce81cd951df4fd4f5cf53a73beeeaac6147ebad2954fcba3736556c8526124f148d8fd50f2c7da1a070cfbe65c87c9da04c2ec3b1b630cabeb2881084f396c9bf138dd035ea3909addb05750c1856b8509cc1ba3610706a53b7b8b32fc1c5d0789cb619580d1a93270b4aa130087e83d94044b3accb5c1b3d1f6fa69f7f84d4d615ed8ace1de489ab7968943b9fcade45119c0641147e9700756e27ad60c499efa931812a6475907dc10c350c42d1d5af975e81a8450c7c228c5733957ded2e74e1ccd4d3f6a4ab220ca892a3129a00ff5e6ba6cf4b2a73b29996baf99bf3edcf8d8a971d202301ebae351e0db681d598edfe07a09acee28daadbd882f1228ffd73fdced5944bd1d0f40638b8c56669eabf6196e951b5a24f2f3c30b301b265980d34dc03f80985eb9fc1003609e9f314170367a00afba804e765931d9fcd2f977afbf58421aabdc4a57c2ab0dfe90d885c1dccdb146274d74356d33834145b92da406bd2ad4db1dcefa837adf984e8e7f725b1c017c15512bc1894988622f95c29315019ab933ab193e86b8cf74e7e68f21759a5c9bafd35e7009c3c112347c66cdab7de1e62033a9f1d1dc93349822dc84b7e19546d745fef6a99d1696e92cee48f75465a0d7fead0c88bdc88f07d22c3c98bb3694ec4c34a63a9c7cb11de475;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h4cf2e6c703be7c1e18556599faaee0c017bce3bc4f77ca7484bc919882446114b3c815bc1f90a2b90e49971f7ebf607991ddf1b6d34ba8b632aef07711b8c80f9ab9bb7816f7d20d0dde973b2e9816c5f6ece27142fd86f6aeb442a8b9331a2e99c6172039102cdf1ea68b42d0d47920bfdbbd1a499e5e5cf470163a5c214cb9da25dceccdc9b96b8e4927590596f40c28bbab1431a619975e98160a96ea5a6925ffc585965ecdb59a25f1d8529fbf86f4fc84295df7dc991d1113451f81d91324cb977d44e3a9fb3affe558d56bbcbe20b7e3962263487111526b23486752321817210aa5254fc9244ebfce70c83aa4d023e29d5631098bd2108ec8ef00744ed4cf6d809e4875c02df22a231097f50725a90934e8b599730d34c314caa4d27980f84058cdbaeadc6fc756096b9769d9cd2c8defb6795b61526e33021f687926eca68189ada6cd9ba14321e93c1853439efeb0e50ffbc23a9fa84b47316c8d6808b4d7067e14713ee1246523e4b6b9b39277d34654d249721cafba3f4a1c819a5d28a8aa91d2a2db88cb6b795cfd87d25f28fcd01eb985d35a1677b2a63edfc06fb52a1359424063696ebd04d4044f155d2e8a15e6cb215d85fe3b2e83ff8d3a12970f67be8577df1d8f8abbad441f3e4fc57cc84b79d3e9d765c1ca4fd57f58df2a6208b5a79286255a890e7ad0ed33a847d1fba88b7ddb464766ce11eb1684;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h99cfe5519f0f22fdb4f86554d72187c27efe3a8cac4c6046703d26c8dbb9a897695b1cba72425b4fd5bb8aa5929e3bb2411ff386e6fce023cbcf24e2e6b36bed9414bb9864a217f9e3dace104cf500f9098d5dfa3f7531486d751ed50c63e4479a7c6486dbbf04a0a04bf3ece738a881ff1f95a9752fdba432d9e81434b865eaaf2589f1a340e8eb30fe577edbc09e575415e2036b8a0f03e8d38be48d5400a31788f044a3ed5834adfc5873c30f27460b38e01c3048ce6f46a982fab36f45214ecdceb0b1bad696d32d498f81f229318a217517438ec14a1ab40947ccac9eb1c3acf3894cdab393fb4c85bf5b0ea1ff9ad804fc02131f1524fbcc6f0b8f04f5be3677260189059c617bffc1a383926bbda4d8d78dbd5996c4234e2abefffdd184a3bd94aa1d9039e99a6705664ad07f6890f52b2d36d91ec734b6898ac4514120c2319f133e3f074ca5ac4553b4d6430131119831ae8a5602d96dfd7e432164a8383d19c11835b6488bbd83aefa153d2ad7271eef5b7f96516a5c98762cff15035c6127f431e63176f22c4e2a35117b1ddcf47784eba52e8f7323814bb25c376d650953ae3d914066556e1b36f4915ffb9f14c67eef54ca37c4c10b3fbfdc782902309e51872e223f009c5f170f81958d3fcdd2c117e65ecf903609f4b3243fe0f4c2979aafa746ad0512877b2b4b16b226a1b1fc87af5e99100c39d1ed58a6;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7a78c22f55dac0e6e05a5ea1a61d41b2ac07acfe7a0ba53893e75205996c2e7824ae5d52c28fa2d4f846996b5c3182b48f15502942554c2a388d67832419b220c6a64f7c0871d676f4ce2412c6f129c8ca9083b6250ec3247056047162694ec61c4d1179ec57e61682af0722952e209e9c9190c11bfe7e1c0a6658c6435fccb8949c5fd7236ced77b86af0b924584727bddbec0011dd8cd8679aba3c77c3c7d1f928380ac21f659cecbd73f1ef3f09ce510229ed188371bd1463a105a82ac4fbe976f21a389e238821589ac21c188d1ec804bbaf692af7b81570e89b601c95687265f85175774bf3efc3e8f3e645e73aaa7fc3496ef1178e8647d352cefdb05aad71701a6de2389f091cd72fa39fe6dd477909cbecdcce42170b699ea4eff363c8bc21bedbb3f38f0f69b17d0f487bd215529b38f861c1c4e83e379e0132cca6460a208ac1865686800095bd7f94b130ee510ffa3ac4352f84ab969b3b72ce921fa7ddeee74205686f8b1c6875847209563f529e61410dbb522b7ec4f4ba53f8c40d55d68b9ba806fd86b7be89f693f3621729b3630da7da91996fce3fc7d5b79270592f935dcfe347662c51951bcc2065273f4f7a6c61bd874e86f19b1b74352973b2a0bfa8681999fdc35c4ad795b7d8a49d48b07f02f0f2f2f9b71e6d2294ee75d6469c5dc1175922ba069647246d870028c427ddfba70051f5c485730ba3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hec81be0a8f31c4a578cd957ac15912bf8eb392332e5e6efd2674502f54e6f886a509bb1d019c793ab4ab5626bb1f974d937ad1bdce2082fcb330a95676ea3a37312353c0c350ab33737aadd80aa3aa3992eea3de89a3cced08d5e1cc84637f50f10f3d8dbb2dae5440a9d194a580bc8df53c483038bd4d22b2afbf68235a85a7dbf82c7352f3033eac1a2f47074a09fda072d061e2d74405dffe6522aa7f7215dac0ebd5e61bf3769af1526c17c099d38c1003c3a9728c2205cf05e496b7af1c9fa6bedc89c9d247b18b46b21a6d1e07a681e14a03f77e148ca7565c1743a8a0b65096b062ef6f7bb9d83a47b90a851dd60a30d1aca676de92315c89a1b0c80c5bb6396cdeffd8d778a011d218a41b93050e1d68f148f258c153443beecab4aa606d773191a6ce5e59f689714c99eef52d61a569ab4995a7b967929f528328c2eb85717ca8b68cf61078f04328a52f3738958720a03d2d257abef24135b0ab3adeb1c6c88e0c3fb58d70b9dca4131d197ab09c890e3d38929f036c2505eda25e31c742e148c575f8bbeb3c368e11e146310ffec2d2299ce0ab502a748a87576ce9afea4dfd2554b9e162fc6771f6fa37ab0666d8eb8554c41eba4691c67bff2d3c493bf15ae5edb3097e0decd82ba7b0e17922c8954650f9d8513b26b7d93e0bc87fb2ee14aca9ab1f710d13554e65dce6aabe18b5d793dd4fb1fa2671c254d7;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2fabdd50e0bf08739ef2e6b5bd3f2560b889b0dda8cfac8cc21baae5e781ab30a72b7f00adb9b5a38525b4b4edd64fa3c6e0e772cfd7afab24fa96267dbddef0b4d4af843ef0f329274a52bb60f037eb4f8f737633690d82a7a562dd9b7fcc918ecf65f550cc04d54076172e5124919f0ee1824dc284cc37fd9f358050c2327c2fb9b6eb5315f546024e83da3455600ddc25fd2bf53228d7b5745fa5366159a666b8220039e08d96a670aed344ef7e5218aa559a56ec164efbd01c3566ba3b881125da98930879ea4a58a3f924a874f88c87177595aac3f15fdd94a365cb5461b14f2465220294adf0fb13d03a51295be840d5f51178fbe67840557b64e07f5b1283beedfc3cf1cc7c0d878c3773a9df2ba7ebf10b384d2717e4067b46938dbdc101c05b5c0cc37cf3a54ec5cf4f3380db5aefdddac7006b0e19b0064bd5079b8344d452b0a150663ed6c3c5acb1fd073d26e748ccadc0d5b735716177768ccf151811c0084c1eee770275896b7d6bf949f26dd3b92073b375761e6357efcaa5d1f88d67f7160f89508f1fde70ee88b07bf3c254731d2d509648ff9d184804dc6c48a2dac8fa30ac4eabc6da099c174132f0a0e57b66d52c9e55a0f5cfa2d3c44feefff98ae7c965d224cf823b3fe0a3edfdfffdf37a51b6873acb605686641bd3894cade215527e7d52c78012ff94d99211aaf78ebb8eaf9b80d909cd0d643d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6cd0a445ab8687a23a10960352cc1dfae6c41da7b1a7fd91b80312d329bca98c526520329a884dbf4bec9781eb9e248c273dc347631e6c351e581effa1dbfad110271bbe73da5376c2fe7727da5d524c28c00dc358a8fa1ee7a3e4a5b64b1be1cbe0940dde8a2b1adfa9c21785c623b71a1c2f0ddceabc70e3dc4002067dc54a7688faa3acc81b8aaf24ad2d5fa606a9cd340435aa710c77542b0d775bff5bead3e1715c0283af4fe5b5e37a69b79e13647e3f4e21d736b40437e15ccc58aae52d705e0964a724b008cd4f5ae64d39da7df3a281e495dfc7a24426caeb98bf3b9556c629547a397909f504e112803172721fcff4ba12d375d3a0249a0ab29a9904b8b623620bdaaff2fc31af1d674b73b174b946defa5bd78bcd672a4462771f734e6fda9d7b51b205982b0a89702f2f986841f9ac31da14302dc913b0ef5af7699d44dbbdf15351a7c6b67f43fb94d907da7c2c239b6b226d662f78f327703444ece127e02842a0feebb5b0b392c198210a4e349d5a9f67b2ec59a12c5a8a6d76e82c550915b83b328ecfab904ce5a1aa5ac2d21a87156d1ea70daf707e203ed90b19e72bfc35132704a1a8baecab0cb453706f9d44b49f0543a9d11d935f8830e1f75767a3143f61799db982c9e3ea31799cb45236348fed3dbccbaf0f06c3f6172daabadb3b73578fa2197b493f2953cde71cee4e532c1d5b16d0f7fe06a3;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h164d009b0eae443d9ff0a145d6009088cd1b66354ab3cfa8a696dc58beba76682bc90e5bfc1d54beab61443a7f97203f98f4c2187d22e5e9e089e035536025903a376cdea85608573bc655deacd0300af3affdbbcd3499958719b483a75fa40fd4c1086581786e6bbddf1afa7507cb8227350b03ae7f9e677c6a7d730a9f8d246a9a307bc91f744022287e0eccf020a8aa10c735eb0209f9ca47ea4c932a06b002f88899e6fd51e33588c6b2791758c0f23c0429ced2bf8c9a6c4713367f1b067afcf2a061e28a2c77e86639a9b8d5a5e8dcbf2d0b0f1ad25290c446e90db792b1f3b0ff1fb8cf15324909e6bb247821a3648567e7979981ccbc1c67ba9c94873b368ccaeda7800b66cf1aae3ed0be32197c15ba1fd4f3a59760a750ca613bbbd978c1f935168493fc18003cd1dea2ee1889cb72f0858d30becfc1e6dd5df56d1a950402fae1ca142199dc8a53821dd873eaa1173c7a86b991881e3cb3c0b6bea53ace28104a42389d91ef6bcbb4a01177dccdaaa6a24ceff491342caa13dca78c2b9ed513275e3b0bb08d8bebef65878738309c94165b53b5e89ca84d5ca10978d724e6b0a6f635f5c6652925914806dae04f745a2c65e843241b2e364a8f2f8363f70b434d68f7de518adf3720669beb44d8bb99e8619e9ae2cd99be835f63ffdbcf664a580e1a95630056791c0f48172cb08e228fb8208f48becfb7322f5b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h538804a9828d0dba9ad9f802ffa1c59462dd873de50ce8a606a05d49e98ab46cc2209db1caf3e9005d6b9e72b036a7e843525d07892bbe10240e3bebaaf20746f091d331c1967660f6bd77917ad23fa45acc004de36bbec8290653c47b0216cf0d08595c6a0175ee353c00ebac505011abc1b1d768214aedc34e54e263064d07efa3b70a61e5a935029460e987efa738051a7dff1e3dc7a8fad170201f1191e469ce36066cac062d7904abeb15084f34305869512f7074320c0aa93981c4607e26978c5934dc66fb5eac78d02738ddbbecedb0d9e7ad8ecd18a44d78cb913bedf76cdcd5fd84524cb591bc1bcbf26ececcf537bbcf85470bd54e7102a78f58402faa8526da169fbeef530f28f8515c85802a0212c525f9adad9756f5f39abb04f5065ea0dcbe4c9be569fc61fda119767e39751256a5638fe2f6d7d33b8d1846272d3dd1f44bfdf117ccba08acdc59dcac9b278ed07e85a73cff6d61efc8ba6e56c09fc37f20b42913ea7c5fb20c5a0024d28ab52644341aafbbc80aa62a29fb91ff466221b6a440780b11fc3250a3fdb7f67f215bb61e03bb88a59f3114b9fdffb94d368914f6acda423f2d1172dca79fa6a4a8747c9d3d8f89499f24eb1e48977614f4f278168599da11f55e6e0f67b1c70e927851183755421b609848d4827fb57843e2f3fcea592ae1947eb9e25cd3ad006628abe03bc1a2cd9080792e7e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h28cd97ec84316eac91a4ecf6410b5a946cac9a3d4e4a575f941b7b7bb0a8c55885a48e33496d4ab3342375c59c8075fdb9e87139e84da66dc07bacd4837eb63ef612e27476a6a2e5be3d6114bdb4b9506f649db3d6b9da0966a98b632392e2a4e0f28f2294d9e0c08901e9ae5d912b908dcf49995f750a93ee3700984ab49e8516127129d20dc05a931dd1b2e941fc808973b12fe2071a83aec7d2345a9b8b4e3696a0246112c1ff34859de2df0400efd9eb3e95c510509dae9d49a1c639b5f0bba3a0954b1731951fc6687e27ff0f11dfbfc30a86d10009a4816343278df5b4e030d344fff784b7d5d7ec12132f64f6730f32ba46c019576c11980f6624aaa28539052e5025a224f4d34e1578945e2cc6ae3af326f472eea461b4f9f5eeb68bcc71d7967fb7904c77fb935cc2be659ab94e7cdd46b9ade52064ff7308b071f9e2b61f8396287e78273217c462be443b20ac1dc8254c46f75197fac12f811a24f8a8fa6014634472601bc5f0fd3b090607590a813465d5346ae5458b9fb00fe28f3995d16a87edc911c179469676be6272ab8c11a1f168bf845590b43b9c4e648762758d8785af5af4260db9266dd887c4f8468b2536084d1bad5228d6be839c7fec623028d0a632dbe29fbb6cd1141442136e4b9038dedf0ff633110c6a53d0c75571efb13feaf5433c10697531a13dedc28e4fb97796c43edf172a89d5eb9b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf22bb2ae4e7a9547e94bfce1f5aad88169e05222fcf8ce3c7e04aecc7f495906d6854e79c5427b114af4f3bb76cca88c5778eeb1ca04555aa1d7b32a154042e88da6bc803042ae890b53a295ed558dbf921195643e8a0a6d948aee4e03130e419d55817055f70d70d330259cf4c085348b2502d5292b658debd606042c94961e6be60455c73935a8627453f13ce98236d17033d67ffa52c680738917a768722c329a2b4ea5421350cabcff835549ffd2d4d443babaea656ebc96a79e85128da45fd1b08863f29bd65bcb682c54b5910a5f735057b3769bd46d1753042c440de77471d97ba9b658c2ccb85ddb3ae81b47b5bcd299bdd5d24d9f8d68da90feab6d61dcdc992d14f7331b5564f9b42533317cc7a57c804b98076f990ae358084e5b8c1450aaadcd4f356cd74d2261d878b0f6899725a7446557e46eddb67fbef1ba804cf51faeeffab1bfc4aca4f4318c630898d4cf00d0cf02e46dafe9f3860e417f581f8c479ba282e4d4e6464f502ac6da03dae09ba6fc63fd408363e33f8d24ffffe6d5fbb95b6249875b40e71af993df4bba25def2aec0fd87850eb3feb59d103c6d9d5f100752dc0539f25e24c7347cbf4b2e8ffb4ccf8c3fac3624acf87122a5940935fbde0763abf1f4c55adc03c4b1a6ade26e9877ccec1c45e365180b261c13dc9fa23893001089727e484bc6371f8f2a92579371a30a65ecf0627e55;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h114fe08c4f859adf2c7bbfda89dd6d893826fec0d738ba539b626f48644bd45bd89d5c3eb10768098724e77298d622bb5bc57d73ba4af13f0ed2b404b0ecdb2d14bbc6921cf3ac128fe1350c1023a7c8dbc406c4066cb9fa1d3586393a98de0d350230f0572ad175a424aeef145c549c3580d23061dfa74ab28a5a3c201d1e6f1386fafed117f9c36ccebc5016a2d704cd535ff0b1b0c70fce3ebd4867b874b503d375557aad67c08b850cc884644eed90ac2be337740163e4a696767d4e03abe69fbd1f359d213c4d24a135680315b584fce3cc6c3b6dd92f097ef10f10ab1af04c8ff71982cb57e1b7b739d26f16a59d221768db110b23a8e724b5f2e00f5a435123cb1c5f4467fa808d79b367974342a6c065415c90e9a48584d0de6d7a20fd3fefd576f47ed416ab659d3f66c9cb21440f127bf933d756b49aa2adcb9b3a797190b3ff0f838fd33b563d966b23383876d73ca4d0df8270504a80c5c41701b3288dd3d2c1061d48060ec8676cd06e7b6e46e24fcde12412de181f9b8283b8ceb1004c5dcbd8053fedf5293abd71b80cc9097ff9170259986963da5073f80d15b0c73e37ace47e4ffede3c4e7c7cb82754d54c5ba1d2bd6023276da6f1ee7acaff22f165fbc6f44fafa6a4308dca3d2d4fc8220a446b6e5756ce90c5ce59af29428a5981a10edc6378937e4fd043cba80d38b33be394fe771f4a97f598d27d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'heb6a5d376a04fe157cf82b6aa50f92ed07798e0c486f02a4e6a3670b43df209a338d4c36d421219f2fb84aa4f700d89082dfc4f4eebd9d171b205ce4350daca348e82e694e381cd0a4f1065fcfad107770f2ba68ea5a522c0428f1b4b6bdb24cb86e88d4dc6fbb62d8b75ded5340ad0d6decc7594c04f00a4984c4ad21701ae21e7917fe6e0d41b7a775bacced6749dcd1f26a22a3ace15a0c854cc04a1b5cd6a34757b26e37054eac9ae452a82e996ba3a18b648295b9a8f5401c29dce48a63300299cb597e7830179f1f765dfd5b6a0e10087adabb65853a51b7de11e0d0f08df1fe4fc1b5a35e3bf2f1655737a6a223f29a734d9e21fd8830b6065846c2da0eee94b4556d0704214fe766decf196c2df4097893471d531eca61710bf5a7f1337d868b5f2d7ff0a0b11feeb8c91726464c8ae4e23732fc7ae9bfbbb72a1a08d019f9bdc03548a0b117a6c9e71ce09744349dfe725fe1a547e10f42583c1dd4ca318dfecd94648dbf08da87e1c27409c7ad27ce44555f2f7ba5da0f3bdb4dc34af13fb8d09fe80ea726339f6d559b861890c2f77ab8c1e7c1daede034190cc2a10fca827ab441aa2b6a01f7cf5d893b6e024ec7be5a77259977b5b08e584860785bec9a81985f132906f52717cd65197f60bbdd2a4309af3d9679bc976708f42969d115eb5585901748fb231a24d20eca08dd987e0b0a8eb28e5ec81a2dac70;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h584a5fe7233ca546a0738fb1616971dc9f455371151db3fd0049bb5a2225c68a815064f8061a004cda73cf93ac41b46b69cd5b1f597c053c435e76b999e9ced39f2f4ebf407344ee9c76632b5a1d80b27e603583817b559bfeb3cf55786b92b91dc6523ced98f3cd963bb4207d5a52f027365eb6e901217426269aad58f2e9326b54e2e17d89a1752a83b2c082cd016d5ba8a16b0611a896cefde34f662e019a1c146a06227d4110fd9e218e00dcfe81d0e575c85a539232dc29d0cacefc947333ad2c2737cb282d37b5e3f464fd5185cc730d6c576fecc5dfe692266f46258299ad52bea986fb42717989338ac6e72d762473349daa129bcb3c0ad2c36d637fd1fca6834dcc1d462cf093ca365ff12d65401a7bb706c2a40866a7bf928d6c2ef15c1a549b93836e85e0eab29ca87734ed97fba053e3b68fc8b87455e7f21b75b21bf934b380edc1f88aa72558807649ee097b808597b3c476ad8746a7fc9e96d05761db4147ab0d4151101f1c4b7c17f21e0b55a2eae14b172e98de9aa489020c8cb6e868a0f6857d54fad6443189386920fa466025fd7c4dd9f2e92bed63428a6861680a02365b84a311f9d32f2643931e743c226a28b624799a7ec4f90690142c248bfb7ab809d71327e6f23418c9b666fb5410ff69ab8296691dd9411862c19a546581a813e0f9b94f5339b2710e665e8d10703dd0c23bfd33a53ebebffd;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf6b0100ba3d43f4d3c10240cb14c5f156fa25df3f0ac6d895749f027ccf5b8f35a75c84d1716b72aa8727085e22633e127bf4a0b7735482bf2acf4c2ccf2f937004dcd50d916f15c409d962c34fd794718ce88348872ec18d4963a66196fe517a2bbbfc02240bc343f7b48f171e71f05b5cfaeb34a3cd4d83a74be707fb13504b4761806f30ffd008c17b00dc7a7344e802986e7b300803222ac098c50860183335718a10e0a202e0ac681de33e4cee5532c8c72161084358031de4b37dc29f6649c6d534382bbf76e65163cff19632d5f5b2479d9c698c42baaf55e3806aa4cb0725b6a1bcfe3b2e2f7d2336ca13bbf5d0d14211b85e7ef66f6474472b60005430d67fb69f9c18bf1f26012207a393f8e47798fffa7e20d4f6aa95f7112d5535d5a3b98cf5d8a6c4662f8c9af28db9b2fc047b4c3f0c5724ffaa8a2aeb22eac69c77b5859c9f6cbc7541ddf1a6a1cc9096a775d30bfa2f15201a77c174aae556f59d0d101727a0b50f54f339bd9c611e0e93a1b95fb012e78d958b4568ce4c34ee93dcd60819dc9f6d846254180f14452b9e9de3d49b9fb9318fcf7468d61e7d1d13ad5b670e7ed8bd709a54dc2897b0e36c53f1c2c41ec1192cd03712f43f3cf9ff797987710fccc6e0c44d383edd1520d853451db0af2cc4c4a9d44bf0108f6fd07109fdd2bbaf3a6a7c2d6507403086ca72837ee8ebb1359cf7a0da17c8e;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h6cf25190b2d743bb5862cbf1e7eccaad59c453722329a0c8e412755fe89f032c5459b6b3ea4bd3dbaaca005f425b795d9f25c43137671b4ff291837fc2c56568462545557466226c4c894913a4cbe30ae8835f5af6cce395365017dfc119ceac3dceea247f572c561490d1ff9f8560a787f06354095af77b2033cee48b79d55cceb2bda2dd6e8398dc57b40ebf960f7fb07869bccd13b60d7f980b80d082a82207e3c9b3a4e53c46c5e1ef1333511681cda24dbbf339f0506ffa1e8c45f0e2332a84179f8e0be9d31422f338b359909a45fa490ddc2052fa7fd62b29e96feb141edfa959248397b97e47dd6c421c91b156779d02376c97d6a740d9a6a5ab6e17e08374d93b65245510eca97eb7e33b21aa0c18b050cc63ec7109c2794f71c6b8a52fb95a0830cdd16ac744786656f00acb64e86736f698129d7bfca8b4dcddf161cc571eee4d4a72954da8d53ba4abbe43257e6e8199fd0de177ae1901ad46006f15377d70a78e4b87323adaef3c181d0dc920637d855081207c340401ccc0e364d53a27fe3bddd914d1775ae3d345989ca3f0be7384eaa8787094410df7138f024234ee3c8a0b4d05e151fda6003b7c148c31009bf51fe4712d73e97e0ba0f96d6cfcc0922f09c3c818cb405113a22ec1bc3f6c18c061f435ed16bc47dd4a676f030ba41c65c47ed87f8d8dae4445c23c8c67f1fa98f2d112780f4cab445179;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd3613abbe2a07179ee88206be10f8af335757557864694ea89ad95f757cb900cbdf27cdb1d3dbadc1ec33510bf185e03c4cbc509fa994655ae5f6000e96117871b844ddf9d6a0ffa4c263e653278a1772d565c3b86631716d1989bfd1cfd465b0e9162558710fbc0e8f134ce60d584941a4c7f99183adcd01c94736eccc5911d0b50654971a411c933cbbd55b877421313b0a411c640a9dc8548553c6fb1425a4ca39bff490e695db26db490b6e3a3c846fbc4ce6d2f915ae89367c18b53c0a215e707800d3a8cebc47923f7b833640718264722035b2b4a76c4bb843b35ecf0c0ce295fe8ee105fd5c10ca3fc98413718d3ea9a7878c892344f35c3a3105737e06a162a7fa88d5211f96456e65832bdf8b4fe23fdb03466774f125464b4d6e7edfc44929ea0f2c4089bb845b32ea06eb95223c05bc1a2f32cdd782699ad220fa6e5b9225b986e7dd7bef4ca5dffcc541ebee39fa3ce78ab0b888ce80499cabf5b50bc06cc7f5b3eef423b05c0c31a5a3c8718c761ba0058332fc049f7ddd212354ee88e12918140c1bce47cb7c2ce963ce3621c1a90020905d7b7364ae45e2886457c6c314d08e3efe34459be19d1db18e18522e415063d525347e45dbaf0fa48f32c2e45a4f25604326c44aa1ef41d7cbbbf4aad61547e8f315fc950b4197e60b9af9bd38c6e0d59cd803de19f25a2f846c443227b6ab7819b3026c1f05048;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h342adc6e0d39f5ffcebc05b4dd0e96c594c3b30b7f9dcd041142bc036ec904f7fad0d7720cc784647b47e0f9cbdb93a82e9d673db2209cc8de0847a0007654e7a9c71666dea849bc4e7087724c78a46375097ee79d03fecf3723c3c7478f88c018eadfab94d738faeacc52b10e364330f195a181c48896d72cb13c0cae90c424cf9a14e60ea3b875c584eec84a2a26f8bcc078ccf4fc8d70eb083f3a6e8c2effdf322457fc6626e759a29b27d1b6e97e4baae040cf6e429162af16948a2ccf8b323547e67950de7fb70365cc859351cd007edeabb4da097afa8cb15348750d81952307b271832dd4ce516f52950922aab7280c9f15baebce3d39ae8dacff40360294761b3ee10b31504f1d789b808891bf98fc06baff183f61f2f051c774ebf0a411ef375a66956642e689d40deac4a644980fde3218f7544e134fe13530c56a89865bc627ccf80dbfeb7ce13f83112bb2a170142d49ff5c098ca75290b975d347332be74631d4e503e4e89a7f5799b8d88e977d53a294d102557429ae0d0076fb48d472c9e5b2b388b9c5d55308ca0a1543b83bf1c726074827947db050619c118ee6fdaf18a832c70a78dc5c2f0ca5ec34afddbcb5d72f221e232634c8caf197b5e4e9487c96124bc80d8529ce5c6cacb1dd8d2df85766f3ab70a4ebc9bc150dca76589c9a286342d542e0f269453858ab398ccab4f62afe94a24cb03801b1;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hdb1a7d7324a7dab3a0cae4027f949fd4d93ee8d628dfbcc4f6ec49c4a084ce6aeb81ffcf6b3b184d7b9845d3e1f40a7c6a1705babe0d24ddc445172c4bc13eb58d0ad951741cb702ab4330f617e4712e3bc4aa15b58a0065497d947bdefa92bb820f83328a247f373ed9a30239e4446753a9bc576b934e3f1797b215718ef9b450bb7bd926a96137312114d9fee0b6e2e5957d1b1e714d0d1025acab79cb26e25d8551b3fa786416a05b07a08ba9b1e17144e809cb7d9f80293242cb8c94417251ae469e1856c5905d6ebd08983eeea97467b8e4662c6b3464e06d4ec448abdd60eeb487a77bad47712e96e38707fe2efa730ffd177146cb31504f8311dde82fc5d965eccbd9670f9bda49090642512833c3392d507c81234d0eb0434cee44035ea3612013832ac56a35b43648437f875849493414c59c852324d300ed7b0d26c63ebb4e37332fa2ba0207c859a2d8ba6e5df90975530dc58c51ddfd6a4968a0116a8657fd6e9d99a28850646b285b159f491a78effa4b3ccfb1739287c07543432f7a885fdecb78670c5e084a69fb8c3ef3bb83f12225fc62ef9bd4a2eef56b175b4b56a66578df41166b5f0233026d514472ff8530b6222593a4a5f861ad9578a8820ed6061a9152e6ff5f2fe449aa5eb4900e08ace0fbc71f0981b7ded7d5356ccaaa54d33ec0d11350e181e188e8a4acdfc098eabbab941e589fba912fdb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5ee30bb8889fb743059e08eb88b53e0f246979377bbe1183ce0192b09dc93c70659ab0d26f7f2650a1a6990e6b692b53d0fc9938a04da8e73f3e27530fcde464fed7b25b6ad7d5dfc476bdf11151f8ff0e58599132c68ea2ac393e84f6f0f52d3a8e88a351825e32321865f0fef4c2bdd1920a4f22c3766fed388c1a5ffad5e92be7d01e90b7b4361f8a9fd2a00b585cf10689836e40a00fe91357a6bce89ecf90785ac8ea0d2f64a813230be86ba8281eeec367778899b47c231a87eabeae435805fd363c292ef5e2c09f79816dab59f6a6b23c363f7ba07b726d5a14511cf6e28d114e0d9a6967709a1beb5717e5bb368567d0efd4ba141139ecec8c3bf2e2aee161626504eea92f41d2cff502cf1700459fd567900fc7862d1dc40dbf08841ce3f1910cafb30a8aad2dc55eb77ec019a94de3bd7c1b397678ebfa697383e68879c48c8a4c59f6d92da6ea48c562ac44f3eab3b398388106d8f09d8d237639092c035c254d7115b317b79ac3a08d697eacae1e5cb280a831c05eb48ed9418e266cf78af926df3c8d2c4fb2190d6f820b47210f1f90339eff51525c471e3fc5c04c8825924123ab13c42c7489170810ba61172566373fbf9c10a201a3790b26cfd78bcc3f2745e82b6c32f6335bee9d5b3853ea3069355f3d98112a454b4605a29f86e4056661d5a72a6a4d9065b09681d5b63ed13b3e7fc0cf6f97f821ae03;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hf9cb3f8b76e533f5286d8b674b9a744ae5c80d4ef1fa6a0bf74a380193b2959c34ee88d51ac7d31790d69723bd5a397e7bbbe66615c2d93cbc87f7bf8fcd1285ed930f64fd45720aa8d3b6d5f450b83536edb59a96383a736ede241ab6e50b36ef4162b5d3200018a05754a54669f31f020f82983c1eee0f34472f8ad6a7b1916dfb66b95c71697ce0fb7739f121576e621d3574ef95556605be179129fd691315e6de2d44084148302678901f4e008d64fe76d2a534ce8da9d8bd61512dcd6710a0b961f346d78b8e306eca5df32b4f4decca016b22432b08313b61769a827028b8608f3f308a3669bb409a6b4dcd206458577f5894223dc3c57eb2ea83c3602e4a9cd4beb3e33e7701317b84419d5e60c3e35a56ecdf95836b7ead2fa8bb28bf3ebef1386609affe5ea67e9aa78bd1f0851a3fe504c325d40b79bc8a3247c3c07ec126642d5f8637b4eff6ffae53c8a81ec39b5cf6351b8942a96e8af1de9e6b550e90b7c4c74b38e4fe70ad1b4aad386775daa38fa150fc601ad870de32414224039608475848716cf38806ba2a74a8b6c5d4dff705f46de411ff36570ab9613a9737fdfbcd9fbccd8dbbe3fe87d1e6f26dfebf02b0dd900f6051fa85242a458e4a3344110084f9a5d8553b22dbcc396fe4f693014a54e0a53a2d964c58e78daa7243c346575700d7faf98574e353bcb791181d406cea67fba7e967856116;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h7370536535a5f72d526964fa0f59c7549b64c1a3b0950e1c282b082309c1108ee6885acf7a73ca20b54241b9175a51a45c678d206d38e6241f944df3b5755cde4949eaa0a5b0078d9664666cbf5a52d9615227dcdfc06deeb907c2bbcb4e0d51530c8417c5154a5a29210a38b67c54d5d8c08fd81938e815830baa2f0f7d0a5d221650ad9e5ef5809bfe95f03cab1db8e122fd26ebaa38377584350e4c6b016f3206f15d81e66dbf14d4553d077c7b793bbe36b528596cce19257c9987a06c6e3535b939f7cfc9a06bc9a95ae1886298880f4d77a28184b7a9e9d4ece5b88adca65d454479cc0ad4f6e89ab6003201f5e36caeff474554f9c1391d3caaf5c46f8082f165e6848824c796e622448f2d6e67d9d9cbba6a33cb6328ab7eb9f095b5479207fa59a859775dd0b7bb15dcfe630eb4e2f1141e15a34876a69463888ddd8ab538be5836d2dc925f334332139589da9f31a2472bd38942d1218e7286e397175fdea6f02fc6bd6206b34ce58ae619ada05a8f3f21fcf519f7803475b9853657fef7cfd25f963ecc0b3275d4f105e95ad2bf45f6e2cd8dbae788f3aca07198315c55c90352694e7bbcb263490f425a782dca8650585a1cd53787e4fbc076b3e862a6843da809c8bb2095dba65ea7be3a2e010c0692a17df5e43c42bf57772304bd9715aa33734fe3284582eba306ad7e8a33ad2ea8f070acd6f60953f1ff62;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h5dce15d3b490462b9e854d80247ce5528e9bcc80d53c431c5defe865e8c62347dbb3a78dd3571469e1643dc525721d6187149995985b7124530a78194132e2e79db44e0db664fd861a4c5a3b7ac03eae4d3b1e8ec673f80ef84e262905d5cb04d65c2d19d52c5ad6a3b795b4c063403d67fa585a685f3c8869dabbd5a79ff719bd58f5200a668e28e300bc667afbd7f873d27bcff7665b487995c52bae7711464df06ce54424548a45a2deca712c810a4831f14c10e1bcae5522673ee013e8e46d81ea49b99b8c07d04386e477730f52828931f585ce5a153fc5ddcddd7157bd27d4a874a787f8feb7ad30461d609d4c6f7d34a634a1ff4073634742a394861128ab910dfebd6078e6d305fc95b45f356065b59d90e794f8fd98c451fc9f294caaf7ac1a42f2e124e80dea9edfbf1f9c666ca6187015aa2aabd7eb26cde79b7074a2a4d47346b42892bf91e42b911e672ef48e8fdb324b1e4113cb3604adbd37f660e464fd40fc06fbe382a0e95f82a69ed1bc4b826766a643f5cf601932b413ec39fce2efd1dab95430998f93ab097a51766908ef931087b3d84bfd2284082447f8d658fc96ce8b860d30fc9d87e7c54900f87152895bad956ef016168b59389451dbf697f10c2ebdf556c48a4134879e371dc9ffa5dc826976687e9cfcebc9c8fb27f1ecc7fa910a45871570e361465a9a9c98afbacce6889f5dca3a58f2d4;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he109565ad66c3119ca54d8217d7a16f160913c78aec230e3cb2d295f20779173c8c458f02db06df53be7527e3f4fad1735472e99068effc5c036ccb79929e8d28400bbce8ab466e4e7d93d18624527a938e95a5311d3db21b420e7b1322d968a71a2be4caef5c0e26a8dd350fb3ec74e0a702455ccf28c87b6bfd53f1cfa04c0ab511c42b4c80cfb8c3a431da146ed286e630cafef7744dcfea93f40ef1f65c3351cdaeac2453b913374a7afb1264480fddd3e1fff7b6f4e74b8eafd989cbe18289162b82ae6756d196e2381eafb4f2aad7159d5748f48b77c431e15db656d544090bd914f0f78bc39a6a9664e01207c7573b6c795806dc310308fc73e99d145b959129448b54602afd02b4a89070a2ac80d7fd299b6045c2e33beede4eb391b75edcc557fc87a6b30fbb8254fb9885f2f3a25b61619cd77747074473fe43e13efe30ea1fbd31d5540b1a2405191ddb5700b77c52d96aaf638e45f796149a866371da241b50eb5a3b2fc26397d4e29fa99be23769e33f971ba825af8d554732301d0c9c87aac69f79e8b4ff68f099e10e268d05bb795408fb5045a252091d47dc776fb652cbb921872cd20800668bc1ea841dd1d42050a402d82bf976b2afb54563f39c256f62c774dcf45018f4755a655790e078905f173621de99369934cab67b227065ac04433f1637121a561fa7d44ec2f376b883f03700fc98b3c57fa3d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h94975b668c3f71359d5ee558a646f252e5b316c40657712d29d9fd470c54643d1ded10ca074440436ee67efeb356b616c6b3e6e164e86d394a7d6c91fb811e05759bfeda5bab92c7dd28a0075f90eb54a937afab3f51afa236cc5798594721621fde4ae53d6ca0d633e7c40f468b10925705c5b277c9398982b93d42fd28a5c4c3599c0246c36fe550eea7c467c3505f7daa87349c80fb9a3502871a55bba5b55ce768ebbdf67d97825e26088edc444599aa2c8fe2654db0e49a287e9a7a33b7cff5c1279091f81567de75d14909e2f10925778ff420665be59528f2accb2c1e507e084fef96186de5de01ee928d60bc1f705bfa4d2290acbcab5655d0a39281caad8efdd1c641cb54e9ae30b9b3fc49558b207beb6e495a65047c2716fae50d958e2fbef97716245004f6639c262ebaa64938f38dc9d33f332522881151a9138908c7d606def61f23437588799453883a40ad02bfa5ddbee3db1edb634576221bb0c2ebefb9d9b866b83019dc9928980ab464acb4c5cd7a5d81f1574676070a64563272f2e1595806ef7e0609c27a682cca181e13580f56e73ad3f46eac287375fcc128b0d5c426d48eee348d9949f9cb4a98706b44f8a6bdc26081d7e21b4b08eb3bee29b52ae4823b0a4b3b56dddb720947ade8181ee7ddbdc0c0ce54dd3780f3bf4ec5149390da7e62428063d00536aa23acec098f08f1e95e65f8be882f;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'ha73242431cd9f6dc6b40504e143e2c4e90711d3209585fa45c733be443bc054ec845a2b1cfafeebdf87d96f21ea865086112ac755d0fc5a8c9f339b92a4bfcdf079b9b94ac0f679871373865dcc100c709dae8ef022a2d6e92daccc2b652e2acefa2f9412983ba4a7d4c5a41871a46cdc3fd670d3c38648fd2e8cb29da3ca23197dcb9f79e62290482dc7e0e4cb6248f146eecd47111a22183e0561a3b74508345bbdbff7ff4ba8449492f83cebab051a42ae60edba801a3d1dc164073360237aa61df1206329bd9d2128f4dc5e53fa7f8b80735fdf1352f52b4868de8832b6c3dcc8a213d1e45d46c1f7418b5766d4ac4f771eb8cfeb5c3ebe34fbd40d3b30a06f37de01c7e3046682b26f276ec8458de67233db9346d1457561bd2f41fd50c69198cefcc4f3d3beae775f1b29a6da5b70a3ba3422c0b03f6d7fbdb4caae9a139ceb49ef0b7c68ae4a943b09376ec8a7b03ed06a8897474a36866a9807497d927e003429ed62d39e92b16d5b76d1d1636d17ca6d232d2bc1ebeb86049753bc1c10479fbdb27027fb0880269023d8a2315ca5b9e07c1b502c701fe101c2735844e1f425d3e69e33323986f1a01fcba52257c87b787a81d4915faedf93d09d39e58952a7f7cc67aabb500a24ad951df2f39eff94924c7f68da913f960027e3aa3de6b4b0c5575abef21cf4dbacdd976ad22d1bfc6db770ea8b7f5f555722e80d;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h48d5b0caed859e93ee53543d426a2833a1dbb6466037799d12f0d481b62a77dca3440c6597109f0d5172888ec501bf5b7ff11bc6e4d38e972062eb0d57f7ec6625feceb0fca094691bf3f60b8b274acd82cf4720392ebe853068dc4fb7217f48e7af84cebd3951d24574c45e8776224fa065298ed8bf7f15d6082e25be2b9697842c5d05a0b809d1e154d783dbc2ea24a55dac2db284f6d8c72143502688c46acbdcda96e31fd78e53da24b8e904c5833da5b19739b7da6b738d9425aa561166473709d8274cf2bbad75265035c5cb7a1cc0ae39699f7144a741efbed71c341ec86aa5d005d9b1008de3197fff7dfb82ca503b18f8199790c5a4a00985de0f89f426be11b7a45f8c8745b59afca2201a903c71ddd7b1f8f50c0474e0e0e48902270aeafcfefc28ddc2d368b50395f9cb13497e791085f569d92a81ca4eed37bbae5b3068de6b0700110963aaf60877998d65677a1c36003a6cb4d0aa1c3d02dda78c30484602867fe24cb1d2034cf354fe3c5df88651554fb6a7858fd276ca05c4f8d06ab438ae8e88dcd5bcf2aafda83f42f31c4b2a85ba93f66d87f2014075dbede068ebbe754b2867342165a30ca1ed7aca47ce06fa92ccc7dac7bdd01a3b7cc939756968747fcf351f13a46acb1febee3bc829be2127bd99e9c48080e87a1df6cd19327a7d4a947e3219bb601d8387c9d7554cf7f45213288e5ba1868602;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hd86c2b1b8da378ac7efdab1a8b26f202b139a532da85ed3229f365c37e1a32d22c01b3c3cf960a899e8c73a3c03d449673ff4fae5af304063946d4de87c040603daca367db1fcac4ee0a70018fae572e7595bc1a2ff82ffff6a1de9cd079118d05368b1b14e2a44c43e88d074bb22f2396201516af2ad492ebda4de9af65b03f634aec02479002139c7060e97f690618337176e7ec8e6879826c4838f7d31131bc6105d0473d3f873cc577fb2c71555fb839c7bd38cc12be466e72710d472131baa5608cafa3e8f8de98790b72c8eddd96907622b72569b1fcb66b650f4f55e10bde836f315a5524885cdf3a82a72397eaede16dabfb10aa0365961ede1798443cf53c85dc81dc2bb0ebd6e0cefecda13f5520881e2801dd52c03cc852b9983ed943a47dfcdc142de96db6463a76c25e0ef2899ffb0a8d980346a4f7631f439976092ef842b6571b666143c030e3729de81f22a670fe0367ad2e8a0cac6afc2db2324201a79a337269e13cf29d2b662e3b6cdbeff4be60c738201fe1f89a3d2ff3dc328c4b8b11d47c12c19b030a76164b3b039b44ab40c7238fdf9dbeb4cefbeffc8831f906ec3483a85baad30fcbcc15caacba88835c014f6a54c579de10bb02548d135e6b680b2c10f7bee64ea070ba6509f2b9c503303d8d2fa0c4bf94626c20e0682af16ebd6dd542da737efebf1f8762c78188fa9cd32a6c00b005a884;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h483ea95691eafa367ffc425167fc33aac198fc8123e1d50de7061a0bd12fb755866da795dc480c4af5ee9e83cc0cff35889defa006419c65f7dbf45a937eb129218429950c4f593a0101fdae087cbb910c7278dfd32cf4413e2592ac42b7566dea67ee256d28b43d28cae83a11a872b4c48b8122d9d527c7582e4c56d531a0bfe68d33d236658252fc79e6534ef83e744fe220b59a6a35eb6e793d2f4481f2b9698d1b5d5b56599b567509f26420529104420ae6f9463004618fb9eaeb74a8349927e078b061352631a0b201ca78461028ff62b951e0b8522af4e6f6247c21d7997799417d7bd4a1829ac56f87cb2aecc40c15850b8b620ec2b4ab265104adcf49643a9fc6ea2f0163b3c9c58c4c2a212e8cfef34e1800c1bce773bf149f72e5cf54baf11c0ae8861e1b94095ad0b2c9370738056d0c7f030986f7419377f4b729f9161807d73d4fe5b26e6aabed7a2aa35a83994dc0f7e6f055466402eec1ef134c997a4eba855ccddad0cab580ccfdb127f266634121e0e7ce6353086122c5b02da0a3eb08fa58d326f58eaeb9530d7558456bb3863b7562814777cadcdd501f85d0b57f9a2206a6fce1fbbe4e41319d787bffcf3c841ceb30a88f6a4e751d7bf1dfec9f91865164d4e0ab36746ec990eb0d21b5dc0d025645ccd428c77d342247eb0dd696168de162afff68334307edc22d197ac16cfa5ed4753809d5b773;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h80c7f7d3d6b3b4eec281db77c3f33a3596196b2e7993c2b330eb034e2fe5865bb825a5e1a0066791be708f99899571a6ee989a90a580708d8d44874710a4e8c56410b2ce5a0ddb14a0efd351910707dba41b406a19a8c09ca02660f31bbed2b7e120d3232852346e805a2bcb40cb70a7477c9f8d12925e2f40e1fd461264402c3fd7df02f867216b6bc4c179879ba14f03e14f65730742a45f8410a320f37f3516994a36dcda85f562a17199ad7c712f168d12da214d8d1d8fd88159fa8933905cccfb1395f321afbb9828a45b88e9fb86b22e0494a1134416ab0c0220879ab57c4ecc5ec56e1806ff2694776292bdcc1fe28cbf2773f5869541c78e6de9419c8c7c6888aa43bf0c8cd6bf95d2c996566b3fb18b5871972187d39ec5e0741f6cf4bd1bf7f4472144fbed14992410e04e7d59b72e5a2df738de66b8e95667a8a836182a860b8f2f44dfa1f4559f456acd747a09b46b8a4d62a3780f8af144b456865d2e061106445ece5a4842c0dd9a102cb763b782415276e7af5d27ed02f128a2ef382e7931f8160c1b5d200eefd2362ac44bed279992b533c2c4289fd01976ed5a606ad736968788a926debef28854613f0a6680fa28af1a7d0ebcf9f0357948039dec9547f262da6537bb475a76ebe39c2fc1bda26d8f2416d457c366e65325a9562a68c06761b840622635f51c57e22ece7f029ec57e047c8a06cca3bdda;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1af8f1941785a6df2ef1393460cef002e789de128a07f2c4f2f94fffca5703bbea86328a72eb24c0e183f8d3b3fc6b5f212c3efaeae17b903027857169e3d4eab736c682202b1efb263b77ef490f78dd39de0f51604673a141a5151c9de5ef21c127b52f78222a05e9fcb1fe6362549e996f7a0963519724182cac202962aa73fa18cc0a3c82e43f5040dff0c752c6e9a5d4caf0b31b0092a5fc8b4141cc36cc5eadbd1ae66df062748436b5a0e62baf27f38e2656fcaafabd0af01e95be61795851b75466224120edb7c25403c530b02cc673ae28fd1e21bfc6ab73b14227f041d1b8bc97d1aab74f35d19b0decff2f1197290612059f916262278c27e11b6ab7f5371e767ffe4fe35905a5c7829d16d8cc789345daebf15db1147db288c47f7bb86bd7fc41b160eeeed5f0527018dca35748430ede36e27aad7e51685df6c2a757489b3ddcd59dd95d4cd93896659df8c3bb3f482a80703fcd513ff4571e57883a6f4f4cc8753b0a5188ce6042fee5f7eeac7c8c4c11856a8d9c680e00bafe1656dd3497b555a07dbd34c8beb617b31208899be2ea8f966fba14110b6502d4fd4c20314859ca2a13a19ba86545238750e4b0ab540cf598aea8c9602e25005b1f59b2ecbfde32052e8fc285271b326ed382aafa876ca089c7695400adee22e6f2879700b3e9ddba55ef574ec4bcb555d0d0c51bc9fd4a0fdb3a71fd6885740c;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hc30f0b2e8f8ca0829f14aa2167633b479c4b26bc41e48e3595091f32d85ac964f94dc6a2513c0cda3c8b88d3cb420858f4b27a193dec1b145dde5fd98504062bb27e5316df6bb22e41019570d554bf61bf0b6165e1a6bb763e2a5e8e9ae5e20bd6372fceb5e7323343d2ae61e0f195417afcd59a80436dfb4c2bcdf1bb8cf2a9991c73b50a7be88e994bc3babeb8d5efe07258eb1380c0f97ed42640d25b8246d744eac2e39205e4564723f1b7c53b9f0606556322c12f36a0e0264892e3cbdbc440dec9158428f427164d1c884add5fa271321d6b35ec91f3913b16866b5a6fa6743a474db01ed3bfe177ea8bcc409e1704b09e9b9839d89cc8f2add861bac69daa2f4460fe0f955bec79c0acd54ab6dc58b284ed13983070f1493e7262b8aa76d0b87568bb2abf1e615416ae34a1346fcb07b845840fec6cd0b54751f9720d10f5170de2d5e49d88a6d0609b65f21f3a0e45526844deb4d5a3708884db740cf3a2366fc239ac02560dd466790e03b77fb2db05741d4fd12037c6160fb590ce115f473ad7e96f77b6223a06111b647ff0757b73ab026f480cbde17ea202b477bdfb2b7a849a86a1e8479360fda14ee88053d5c56847e852dc10055d1c731963ae30ca4801ef9a48830c08e12a1137de59d15ef874d82eb5b59f1f1bdcb43ab712d70b23c084246629035f63a0c6fcb749e468e2bbcabbbf7ad610dc088dc68a;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hacb3ec81983124435a64a0f88f11e2c7fc14c2a3c982d27d4b4b670a07f92c0e467ceb62f26385ad073f97eb825332a2b6b73460d2a37dcc5c94f171898b78e132139b6a414876cb00a5222bd4fe855ce18fa033494fb12cba97c3baaf844e05247a084bbea86b28bc164ffb52513544c62adf4eb44cbb4433fa8ab63ea7575191533d6282c5571faf8530a9345a429bbf1f1d6c85cc3701d4fa6606a6fed8b5d62f704c3f0a4cae3d8f8fbc75a511a594f2b09b225b69dba363ec4acfe005ea4b8163028b476b22d92a99c087c124a66691c75364f1bb69d035562266dd11306a2bac34942bb8503bd184ad2be310a665c84d5e4e6960cda7190ce2b27de27228be255ee5b13c159d87ba29d8e75f09d01075d91c8a03eddc95cb3b6a5a0dd3c4762fca702e4e09c1f4f55eb864e6b57fd2047b3730b6fc04e6d81b694daaac3da332606bf82c2f985d24fccb2c7a823a235875f22ac2baab21630e0b7acee62c1ffd29217a45833ee2098ef70ad8b2c9a37348d88cd440fadcb9b39bb21be4f24ac8e3fb315adcda6c3c2a3e0a08237f23b05159f93dee825a1dcdcee37cf6322287e7c29ed1f73cc2fd256490287c9a9a64a42c71bde01b6887fce57686ec544ba835de6980667149efc6fa8d7a1a057cf3b30f34194cde579b972a8105821d3690968af17583ea626a32d0724ff3235e4017b8e8b232bdd1637c8d02347;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8c15f718fd3c700d58d4da747568bb65aa0a2c597d3cf3802bf831c1aff7e3a7bece720b578109e75ee75bb72c46d38545a1f51d0d7a8831cf9b0f84a7567e5ceee2210eea46e0e4874d1361a2c15f3dc7dfa2d836896d0eff18dd6ee2eb6f552bff8d28db78960ba7d0d9bfe30ec421b0d69e9a5c4c3b5568ec6c437615db70e7e2d2098014bdc8574aef2c1aba8ab40aef4ca41a17ae6b91ee561ebcd763ef769cc774a834b23b70d3bae0685869b0499ce1ee66c4cee6d90be0fee05f0264b1c378d74472eccdae989e7a445f40ac642d6ef638614c5892910e54103def8c3957f37613b80e61754d219119376f59c873a62c7c04308bb26065c9b28bfa1be10501502d7748aa32de9967813dfb5ed9d3731aaee76623299e612a4ab72e8434c72182d808e287e830cc4374bb3b5a38a587ed80e6cc79999235f574c29b5767f7bf260c687a316493896a4cf5434b1a0780bbd598efedbbb1b755fd73c0735c320694eb44388f19d1b3641065a1deaee2a8dbfcb81a4aac676266acc71c0d533e8aa365331132da91a0be83e448322c21c5f18395a2cc00fe12dcf48260570c387b5f45cb4472b298831314d4805aaae1a53111da84eead0c30c48287ad0c49af014f47ca3fa61623f0d27cf8d97d66747f5644e6f431b25734d7aaa84fd6c192b0ee92afc1ef839eb0cc8ddad798d6718d91ce92a2b5c8b33d0e96c8dfdb;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h30fe97ac4dc6005bdfe230e052166e892e877ef43d04869d26ae456a7298807e7949ae835688c0c2427a135f0b900642342874c0178cbf4cd823cb86991c1f0b91899afb4174ef9342204da55c8018157609efd4107adbe419096094f500441b1bd62f9ac98c4b9c7d2efdf7aaafb79115cfc3b1b1bdd258e8ca4fca3813d96a809fd10f4be59e56eef7dcb7f9f7436caacafcd8517a77e9c6e47877c18d321e4b8db949db2d57eb273e420cd8f5ffbb9b9252c576fb26ddbfcf54cc95bb3dd840ba0ad9b08032203592cb9d47e9d371f43b2ac2d739bf17a58c393ea2886485ade95959711f6d41616b46b36eb28bb535e3eec5b4b59687fa6d4aef44ad5bb470d3183b09cc59bc64020f3cc366d7fc84fdbbde0102fddc281cd15dd1028db4fd1e086ec5b19b7b0320f5c05cbd417b14865162c672a31a2efc46a63fe4b88bbfa93e32ae4d9924203e5015b21a5867100cf5de73c0557907525d1fc72373e7abf26b4d61203c405d279007bdf74d34858114de362aa66f376947552523e0b8c9e974061747cb05be649ccb974803ffdbe449e8503e3fe5242ba1974b25bcd40aff669db7c30d9684cf54a0f4d7a3da63fb64a2b519ceab166008067eac19252eb9946edaf493a9119f28013f8301988b97b708abd2e57cc971ea58169ae72feebe8295ca6ccddba33312816d1ba536ee430e81dd3f68f2056530652d517051;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h76428985ab847ebeab141f9a2185b7a1ea9acf4ccb184d2de7bf9d271ceb28538ac00d34b8142516ee8bbe9c1f695de347b27854e33b53783aabd82618b50a99921e500572cab15a05980ea9c5d2684b6a570c681818db0ea89015c9fc0f40145993e6ee792290ae97d1cddcb6f50639a4dca9e7bc426bd06b4408405e81d13a0e05ae9a27a2e8a10793776f0c789cc9a274f27aaf65828567d89358a871f5b9ab881ddb41bb64e5f118c82bcf98c9bec1f1ecb20d00dc61a982ec66ded6cd08c5d54c7c51adf30840bdac25628aeb064dd1dcf5160f145244eeb66948099d19f140cb3cbc9031e4d3250ee6d280f31100e6425788d63d0cab884deb8995419f7d20d2a11afbe0d2a2969f990d68c873fc6eb181da96c7d247099cf9e83f7f63e6efe0aebc1d59aef837f9f5932cf2b8e4a2b3da876443ebf618004507941ab859ea58212d6486324ca5cf83c068c84552f28c85024916718a855374b58c2be2924bc337ec58487611b0f472dcb952fcad637552b38f1664ed359e646a77e54b698a344d21b6d1ddc0ac21d28b37b27ca95c48cb73a008bcd85bfa0aec67618f1c9787ec11677f5a29b73b4eb04aa8298b948b2d416f87e3966bec906c27dfffddf77e72cbfb140f5506ae60f524674e54b771d52e39b4ad46c27dfcbbb1d23dcf23675594b9fadddb3d86f3dbcac45040a0f62e56ab625f34d80454d74f7aac;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hb4b707a3fa4d29a620250ed92bd287ea140493c2ab39b0ca2efd895caf82feceddab55a82d9f79b03fc841f7068e0aba702ababe27a17892e311d269365b9efb802ad8dc7eb86da6adddb60e933581b6351bf1378e88cfec0b8b295605c949506ddee07d9b8ffd81199e244ea01057fe98747824dca8c3886489488dd0264b7cc450a157a310d16778226769a7e6aed97f3ac194850f5b51dea09a4726128dc01f0daa632fdcc61effd8c6af3bfc7d9d705a7a2973ceb62a56e4d29c0d0479fc8a28eb11df210dd4347256006defefbab005ed72e15f85c03bb4198cab44044ce5d16d49d4ab98cd42cb3eeecd9ef8605eed074c7fc035a6c2758e13dfd2bcfd1c289fbdfbb1b18a6bd78d1018165cdce981afecb4b6fca037f184da1362983e4ea4eb7a93d3b1066c55473fed58f9d0fc2c7ad92400db558542d6e081571b2a4663f3ed1e2127bc2e8d0c158ee10abf95a1d624f2681d0148c118c23f2cfb82f88c873b58e4052570189dc65c9f358037d440859f6b6d965b00bca1fdc10b124283fdfd95e4b0b1dd0c6f7f247688fb4252570271cd833aba7208e95ce8f21f0eed1d7abe60a02883a0fd9f12bb4aed09634421af5637c13140653b50be014753b551047d8aedb685eab4c67b50176815e6bfdb45ee6529011022b6236c76ab8b28a25f7c3bd91f7283694ce539614c3359d90e230b9a9ff1ab23fd2df70d84;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h2eac8520131c2e0ffdc7d051221521cae9c2eb8b32a6566c662dc5898cf3f676ea78a99c6ff9c60b529f805348dde3213195140ab498fd1a56b97fe7ae8875104c5690d8b0e5db4d6451946143ce647602242bf0fe93060b63908276026864e36c54edd080f006e1bbb0ec99a45109a72297b22471faea2a67d44ad3ded10c62c12cc393172fac97ade78e8a2e431744d5881971b833340952face45cfd3994376cea379fa459460ca77c8f3ab400f77ef28dc61cab8c35cda1879504530f5ada642cc9db6dd64896befc61a163a14d016e52ac45a87d776fa6068379c0d1d667cd70465e0f547d148da6e343e0c62a4f33c787d905e712215066f3b62ef2172dd5630768dd605ad00aea6783873ca90b8f2947739b6f073daf69fc2bc2732981b7d88f39d5ce26e9dbb3b882f4eb374d57e43067159ba181000bda524f5a5fa55e689b28c26bbc0ae80cb558aa99a6e5ea683d9dc377743509563f62499d7380a6322b0e5958a82af2fc2041eec52d1af92703b4349c18fdf18cea5153da3a4c71548075e462e97e9294481fca7d79322f3b443e791ce2ce79f6e6f740e450ac1bd9f61ab878deb1acb1f5c70ab2e149625126e9ed5596862a6ba71889aad9b2737cf679f41ad10ede1fa5648a7c1a2c3222a1d98f4543f6d279eb7568abef1847c9df28138f4f5f82875ad940e4714868fdfdc6cbbed7c3b6df965956834bc;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'he2c0987424bfcc29958c98be5c84d736dcd001329b3e4f8365faffe3490065a2fa2f71e025d2e669776ec1e5e8c8560a2690c57a693eca134b2cde6a0f90957197b6d734731424ac9635cc975e3cfdbf3005f608be676fed7acdab57e9847a86dec2eed29809ad5a1adee26b8d26e4f5581702d2b6324606b95d2155a1c3304e0f47900d4d0beb0855a4d412fa16299829eb0f3979e70475c7d7ea9e70cda5dfbc841a20709738fa6bfffd4dba464e1195df07afadd789b532fc27ecfb0c7263f43dc610a7f3e3d1861a571c75a233c28f418962ae7bb21dbb3ed6798b671644ba9b9388f7741075c01ae90070a3eb437c266b8534cd35ab48bad00e54de7de424ea50f11a8c2fc888306235c902dc22cdb84c6ac18a3c56e13779fb3ed0785d7881acf5b1ebe1ef02cf5c7e395f6c0d1182469ed2e3fc4e55b8fe02cb7e0247f52eb063bc08cd1bb414b013970551e7a7e3e61c66027b2702fc8de518442e0b212fa3b20cd137bac1e22e4fb6e32681aa27ecbbdd6ba82e755a30c2b58f451f811995a45e9c3e68f30aa9b34869ef557c59591ea5f0722a0d1db604ae50d295ea855297b7e853e00743eef871f63d2bbd5bc3a6cb8d98cd1e8d850dbffbdf8f98539407f4f6bbef49c31961c1a01adfffa7baf5ffdebdfdea5aa5a85337aaf6082dc977a2ad933da3fc84d9ee391b8b2f6e45d0b5ad75448ff97844313cbde8;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'hfcdbc49afcb9e6857c72fec88c37dc5e485cade65ffffef0b7431f9735d946bcaf92c80fe1964206c53d6aeeac7fa617fcdc82f899df790885c6f5129545769d7aee447bf9896656b04f4fb5d8f0e80714a59521e85bcfe69436f1f478cd2fb29fd40904cb8e903a3b24d15b101a813e886079286793d9fa6a86bd5bfe75858ecf77fab580f9effc8ae569854310f887c38a14bb2443067776220f9e95d1432051c165a7aed7655148d7dd14dd302c455902d61781939f91f4302ca178625ac7b246f10f89513e655aff21dcd865e9374c00116c95d1fb0010d6b4b1816e00f13ad2dfbf20eb19d9670942501ade84b3779ec5dce140df9ec706c698df0b165957993c9de9a83ca95532b4e71202dd0e1055266d5954bfee792d1c4a7a072709cbb49fdef530606608a145ea68b1dd6c38aa8077c5488562709f90dfbf6ffc83e1e82205a152d9a91295de05c16197adb18bfc8f87674b6a5b1e2478d74a30023fe7e80d24823e0c51e9d5365bcda666e57d865109e3420a881b1d0bb666bd8e73afb9a95bcfa2fa2af49c0b657f3997e76b21cb4f9943a163c2ae845b83fbd014d785cb0f73e7afec4a5e364f05f6335f8d080a9e83ccbe85f24b369d6b029d549d8a493ac297c9a093fd48acafde5bf01afda90d57424abc90d8e26d6efef12aaa23dec04f3e8cd530847a3913df881bc72899211fc8fea4be56d90858514b;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h531d17c303ba5509ab2e17b956b29cd1e8295490441a56736ed630dc7115a0707a8c60e9a6f0e0d90f29ca5ea88fa8794ee66d931eb87949ec6dc210a3431fbc6e3b01afcaf8766f2496ebb61c6c433c449f7699931bbc165303c0355bce2a064bd96fa07cfcc528a4bb0ef54731789147eda55bbfc7b10c0faa5b95e9e96d7d9ac12c101aab86b2d0206048e8d861fadaf3f6ec17d7874476031fa149d6c89ab4d930e0164c2506e75476a5d37c3bfe67adbe4e8678596c4a507c5db74c176b834194f906292151e953327a4e2604193d6e1bbc4ea285ab449d58479999e9cf461df7ae25e808310be62925aaa61d59001f1a67712ee893c9e136bbe183cfbce3ac2a8c8adcddf3b4f0dba0ffeb5a8fec183eb34108e7038e04b09188c91ea2d4791374d527c50102c9528b876a7a864fce0abf6abd190c0d8fc0e2934fa337bcb3b1334adb219600e99fe664a71bee8127d5b3b5126d4da4aa9d5256fe8fce821e769f1c23b0ffe790c56f0f54f268cddb59ab39fb5b9d8690bddff4aca2291ed8a7e0b5d7cc1d7fef455564e7b2626579a73df0ce0b049d9bd294cca10301ab944cddc81d55cfd1585bb0526d1b8216c1dd30c1b623b852980a3b8308a37a5dd90322253b4b7df295e1e874ad79e069d51db60f21668f80aca615db0debd3658cda18280bf23d0801f4dede36e22e444f7f1b8e4e074cf932317bf3166716;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h8e46e95d975b91bcb3439b6d51461ef8c6ca00385c7cdaff9e33365de1fd6b36d67897aa0b138a53c5597d1ac07c21d5f0f5d17d82b6cee272d8b0a9e8ae278b3107b5071a47b0d6a440ab04022c71d863738ff144f466209b077776f6b7e0f65c505e5aea6f0a5f71ed9307a339e57a24c13dcf64002dbf9abb5d947688af4fa20fb504d1c34f291e757b11ee6cba45e53fabaf80223a0c5c26114bce9299e4c6331a5506f80bfcd4e44f6be96773756864131d828ba3b147112169c0084fc17565fff6346eac4389ac747f188700f13c5b317fb1be57730b5a1e4acadf6d40166320c497d4b2823fe44ff5a4e4cda0f98b263fcc6bb506dcbe4c0e893ba16f04610c6756ad033a586ec35306faa6cdf9fc21d397f8f7a4a3cf8fe3dbdbb39a62baa6b68901502060cb1096715ceadf9d3ac67a9e1b18edb21979044d00c482325cfa87e60bf889b2e11f4119dcd998c99469f1d12d0a451b57614b546f02aac8997e7109ff72360c9e2ef244a96cf8ba6d7b3db3a68983feffd8f030bb6c878be7e814e35e70f7f6723063288565407cbf7481558b60a0fe9c0a3b4432b7721df1486f7dfb351c4183b8283611cc837bb079dba2a6ac30d569bc7840b1eee5c19519095e2e73a30382b1a134a18fc8bde9cb897fac0b3ec9207c785d7a716b16627eef424889a04fa174e99b60eab0edcc1c68d4140d1105f6a8ec4da7e3b2;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h74affeb3df16b231a95f5edb2da71bdb81e8b835356f09d77e87f0011888ca93de269292a562779d223f3551373b603bc251166d7ba9725893b350d7d54f154fdcca54cb969ba0c6c4e623174cd7733b65b2209c67817583df34d434b9b4444f7ee6f2274b7cc6e76568386afa1a5cda9db936df7f22b34ad506f3a3ec2297f2e15152c5ec9f559850573c4b610ccfda53224ebfd6bc296af9e60db68ac8fc8c0a9d3ef335b76032c55a78fcff48d0b5feba730b9f5e426842ed2000ad6f60a3d5199138eae7cf3dad594d55273357e224cfab4aab4411422c63b065fead02a9bbebaeb5708cb69c4d7910441ca62f95dc0e155556f7c7941d641c6abc83b54ce9700e1c896ed2c93389a30ef483f2f9d7a27947d74eaa5f95d62035d26878b37b9f200e23c71b9bf0cc9e791fdb041a0e6692f4c13af1fd4fbf4005d404014c00cd817040e82803de58696761c9a2226336cd7b2fc83e4c7a22d04833e6e4d537d606f93ac7c54d4d899643b57b5b6595b2b99532fc2ded09a3fc2e814dd30f514173d0d003a998f74d8cb3405fb24067513dca5ce58a663a6309ac21438e40da01f28fe1d3bc163292bc4e50f4389ca6d63a8b20250587d84facf576ad013722717af02e46f898f3bf9d2f022286d0a5c0ce91dc23e42bc8bd2955f1c6d062e10426685d033591624d9747a9b48e0bfd25a491039f4fa51c3d63423c7a42c0;
        #1
        {src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 4096'h1e682fff3302c042821be80e4d48a148517203733660842163f41e30877b3d445ce028ef2506ce7acec0e66295ced6176b67a99da3063728c9cda2b59ef63c1ccefd7dacf729ea662c68a60842187c8a864a69fdd8114dc0361ee70929c19078f2e17477440099c50f5230ea468d7c06275a3b5b473573117d1e89b375aedf74b83ede5bab44f1823d1664b45f65ae9ba8467ffd65d260c6cc5792a357afe1ff49c3a329a3699ec1129ba38ffd00ac6a8e8efdcf4ea19695b733242a1533f1d18f231d9c9c9d3ccc261428f617402ad9b15e27126889d84f57fa511a387a0bed6101725d42870a6f387d67420c6457d5ed27a4401dbcf454763573b57ddca180acd53abb2e70311b3b3e209e6ea9c982ce6795a5192bf424274d0c656285e42ae79785be697444af7e799c34c4613ea38ea4a4c88687a8a9e9245d360ac568a8042c03f79c279e1a1d3238393878230c556c275a5b4a60e4d777f14f8a9ab17cc7c5f810fa197eaa40df118465467d20ddcc1f12da2590f2473d23ef9242bce45d036bcc718ceb2e51052217b234b962e9bdbcc28341a05210d1f9cdf8e7e9039b7bda5a67e54e6db5ead084754bb3ab508f6de60f1109acf031e4717c4a48bcc70ac6bb2c49a93b05d4ec014913e6b56da789788a39466b7030175758a48d46f84ac8f62f8243fdcfd1f19ceb9510b727a4d8c8d2874b76fd7be8ff63124c26;
        #1
        $finish();
    end
endmodule
