module testbench();
    reg [8:0] src0;
    reg [8:0] src1;
    reg [8:0] src2;
    reg [8:0] src3;
    reg [8:0] src4;
    reg [8:0] src5;
    reg [8:0] src6;
    reg [8:0] src7;
    reg [8:0] src8;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [12:0] srcsum;
    wire [12:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ffffffffffffffffffff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a6e066fa05e5e8c6fe1c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h57eeaeded7991f9ec788;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdfd779fc6c7400ae27e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14bcda270d18be02af04;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h44c31f9d31ced32e95b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd52a48d3919cdc131345;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12550465bfb2ace6d36c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h62834703e73f72712081;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10d8c32d0e46e20b1610a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d038619ed7854bdcd523;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h145421ce059469e4645d2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h92e4e757f40156af6346;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h855bea12ec31774ab311;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c4d6d49c135d5bedbc2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4b0ed5ab64d0019e0c35;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h175a78471d3fb1cd6d71c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ab4d989b5cd5aac3c77;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16af6579bfb01534a0b15;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c83b17151cafe57829;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he57c1e90c27b0e98fe0b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f383637c9abc9c3ebda;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hefd282428106c3a365f4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bb2f66d083eb4fcc10c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15f9cac2eaa62ff87a598;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1760564bebcc46590fccb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h51c741db3b149ae0700f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13d446bfd9513c7503504;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc137a5758c3487777300;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1178dd9cb6ff6aceabaa0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf3794bc02ec67443c33d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc90dc6808b0934803e65;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6183eda1706ad69d674;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ba6318a987e9f4fed312;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h106adb7fbdb0b2edbc3f9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h156529c55b34bb0f55bfa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h131813bf8b68a0cc1c484;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf54189d30cb412e13df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1448bc495a2f0b192ece6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e47073f4c8fa28dd454e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb8edd44bcb294dc4da09;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h948ace8e93b7d3a0b33a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c3d7bc5343169b3a167f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1113900a0fe1daa81aff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha5b007677678a010d2d4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10ca0c85d10a901720c24;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbbb0fb1ec844e7830e3d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d8c9512457948463ccf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16e8c58edb4592a41861a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d3d3f4f0ca94386a8b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1885ce3afec7f721ee31e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h107ae392ff61b81cf4f28;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e494c3fd2eff6e620455;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b56d88c31ac0dfb985bb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h22fad8bb10aae396fa2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13318536867971358b9ec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7926af1c00d984ad017a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a701253893d32f176248;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb5aa284e58713951aa17;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1967f78bef5579e31f36c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b965aa59111823f70bdb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h87691a12bd6649b70f1d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc3577bf12ca8b2d73e4e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hba1beddab0c47a5d3f9d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f4525090fa2eeabf48d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heb82f0578426999b7ff8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fca44938a83fca334777;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd32a445b47c37943c440;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haca48e78286534f16665;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1255baae50852eb2ee378;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h721a72cb222d730259c2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c9bb26a355bc746f5bfd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1884de4c41f07a453fe7c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h257efdbd98d241780770;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be25a38482e6fab26567;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb321d6b6964b3b152e41;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e8c0f472a9b67906cfff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h132cdf621a20167020060;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1575051ff881f470b60e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb4718bd346fae2169a0c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a20745141749e0dd650d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eff8e4ece2f3d37da327;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1555f45acfc230d43ca55;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h39921e68f48b6d961fc2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb778e3756a72be001645;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h707eeb2fa64f0b0a83fd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11f2a33d2d7c7dea2bb2a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1905094e542fb8f7671d9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ab95a0f23842d1b7f92;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cc95573121077b5a5ffa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1467f3f73aec1bb701e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17e50f5575a0784955514;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9ff14b6eb5082fed7867;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d717810c39e717502620;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h116fad8e259e6a70e7bb3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h134caa1e81d3825719324;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb6ec4d3977e6096437ac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4784ce1b51fb9efb2c56;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12f33b6f7f42f1aba1836;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbb408509f078092a9c98;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h754ff018e1830a4704d5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b98331298f95985ed49c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18be9ee994aec79b8300f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hecd53db9c3945a3a1a16;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a3f3c41cee901cdf9fb5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h318e4c34fc949b5b4dee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2cfdd263c16157b9a894;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h191740c2e368a6526e14c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9762e84ea117ce66a8c7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fce0393fdf3dc9034b66;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c9035c4d8f5c22185a43;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2f9c370f6c0b488f9abf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf06985c8505e46584ed8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8c8577d7ab3fade3eee0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8e7e5ae4681065c7a2e2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5242a47dcdaae0e61361;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6c95156b141daa2caa73;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bbb71ca418e5ad521e41;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5a61ae6b4c3ee24ce250;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h128dbf7898570901ae20;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h179c70d95ce67701f4e43;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a4cc07832cf1740ae15e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14d5fa40ccc987296da4e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cdae4a8f0b4f7ea6a7b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13b6aaa33511a36a2193b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c21c9b832c67ff8d3e56;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1868236928d4ebbd4991b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fb4e1e97cd9e0e5f68b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12bb5d73f5347be122dac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3849f933afd454be0451;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13fefb6e709b7e0cb868c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15840f6333cf180b3558;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he78d414a514df56fb7b4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h56f7e25a98f549cdb09c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd35cda8406b40662c1fe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h147bd444149aa19561f79;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a3d5235c60580081d223;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heee9d84d0325adb3e530;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h70b6be80ecb8d81c5cdc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17a9c292ffd0a66f00b12;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb426d927f1460c58c91f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ea4f883e49b882ba83e4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15eadbad2b0cfa667d6e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hab7c29356079e21bdd7c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3f568d815ce9c7742a47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfc42aff210958a6308e9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c5062cac3fc271c1982;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f92498c746072c5a74d4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h76b0de8b05849060cd15;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ff3aa51bad4a8679fdfc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c857ceaeaf403aad7ed7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc684fe12099af9d2b090;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5dd4b30b1dbd71d7a3b2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13bda84d74478f63929a4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf0ae9405b7ab8c5c71ab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h27663a3443c2c380fdab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18d5c748f3f8be49014bb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7d7e09e8f5e9946920d5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19e2820c3a69ecfc6b919;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h186c5bc321f2e70d8e85f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h117031bea019d707a8a5a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h197ad9d1403a2f14ead54;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h51dcfe05af5175452292;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf5a53f2a713d23d374f4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb02d5464970a34431355;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he74e9fec4107bf7303e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2459f650126ea249b2ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h20258647f12b0e5e19dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h116b64120d53463a20425;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdebf47c3b17140caabd8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c1a50050131f5919e8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18ae11e9e07e9bf2e7ea6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb2617f16322518e5a858;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10a4096b28647a3063cf0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a59122c6adc4999c71ac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd925367d8ac97294f13f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1735f0c346fe59f23259;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13b82735a37b8916c302c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h743a6a9cc903e640329;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b87a5751188f50f89717;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d7ec7feea6fa3cd53a6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h491474c54d75f243733a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd2c4686937af7e692df8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf2787be66cb723535353;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16b2d364d827e7d23d96e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb3a9698e672911c5daf3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d3686d0034c7d891023c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eaa64f0c034b95de6574;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h598698671c2b8c92b00b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b5d9bb7426450320a7e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h60cd1e166d331f30a5c1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e5cb360b4064556754cb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3af59cd1467be78f6938;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d0aace4335774d5270b4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7d36d993a1b283abb38d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c2685e248d724a874751;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h61184cec2fec0983a061;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d566e53fce3a9f21fe0d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8fff88bd35e48bf81a55;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbd36acb36d7b4d1081ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18a676bd3c1eb2509e8dd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a0965884978791ca6a4e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h42d4386ca7f317df865f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5455ec0ef4e857766fee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc88d06e85379a6a8161d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18b51309c76bbf5dcbc68;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5739585af407d17a36b3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h198375fe20549056c60aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18cd75154fb15d3b16854;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a0420277f9ec71d8d008;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d21fa9ce837f73e1c32;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10a268e8a117907c250f3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcaf47df372d615a0d99f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h38bfbec146b17c1427ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h866a50611120dc9c0bfd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h182522794fa5b79e787a1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15517136e0d5d0cf2e089;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h32f97b2cdd42d5bd48e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h159067ece271b00217686;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he2c77f241520b0a8d7d4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1237af1f1e74844e42a12;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h67a555f32c6ebe60d18a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12ba3860dd26ca2e09a45;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14d0989dc56ca099daa28;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h313a7b93d825cf2e38e3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3d5fbaa42b6007b5dd69;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdf8b93b6a395df9d7ba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h546ea181b4602c8f7cc0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cbfd77e4f2422d4cfcfc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1feb00a742ffb3bf64a2f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd37927809bd3ad685460;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h60a603dc7fddc8a4dd54;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h255c1728eec1a102a6cb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdedbf7c8eec432feb2bc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1896077438a525ece183;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h875ad8860b3a5d9631d2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c72df98a25773201ad93;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10bef3c0e2f837c717da5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3b09e07fda47fe8eb8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10d88880fecefb622b013;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d5ed0f99d27a473e1f20;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18e9d33bcc583c27c1e09;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9e5c6dd2129e98325d8f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16666945fdb1d76ea89ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e6e77daa47e556856afe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14d8affc75984ab761caa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be0d4cca9a769a4ceae8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ad52c2bb24dd7ee193b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h141ffd4288fe6ad99b6bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcb0f57e6b0b49feec106;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a0fe385dba577bb5b216;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h185d94b2eae3222689b4d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h196d888446c1d6775fe18;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h225b0be5a841e9039c2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11577d8b2ed4688ed6aaf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h110431c9ca4660f0e6658;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h116d277b7f8733a9895a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bdab94767ea55cb5e543;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h37ea967aee447b13fe6d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h137eff6906ffa26dd4ca1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hadb58ea13d0f800897fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b014339e2a6de5e9de26;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aa8a2af89df1a7be3211;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb2fda988e933da1a5802;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb5de480224372b35050a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be902ce045ce03b62b49;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h151a14d710563b6ffe81e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1529e0d60a88bfe2c655d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aba078c58bb930779554;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13d6f667f3ffe97411a4f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb1eee622e8609761c043;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4cfc3a007506bd88f48;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1347cdbc789515131f3d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19dc0991bc3a1237cdc4c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11f0780ba918141619283;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c40957eabadb07db609c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h89efc0bdf9a4624a8bf6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18c19b069a160a47f2402;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13dd825c25d787b1e4d4c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1951aa6872e96c7044051;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h168475631e93b4595cbe4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1109064cdc25f79629519;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc959b4b82b9741d002a1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h117e75e6475f2f2a2fea9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6932b45aae58735a72a6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h50120d6b653e7c53c087;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h118a10a13acf1a290ac6f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4a2158ed46d013a99848;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15d437248ad443de0f15a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h48c5f5f03f4cc2dce289;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h181ca307a7dec62e24355;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e9643d0d31fa214e9089;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h43e8c22b2bf21cfbd3d3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9b368117b89a748ead87;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf86c9428c24e129a4510;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4ba28b5bcdeb4bdb5da6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9a97b4f3843971d489f3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2c8b21739a8744c6899b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc96d860a1ee04b7d3169;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12103d4e759d02d1b8bac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he98538a237188bff9e19;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h177682c90082802e43c07;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h123888ca107aab116126a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdd557797128f06ab850a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16544e4f3744c3d10f149;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c40d0df0925f1433e138;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf41226f16d9e6486458;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h32d987292e88f50683f4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3a09e8fcd207d31b9c03;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h110e52db1ce5047d37287;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aee892a775245be15a79;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12c8e7c6dba37745e1f57;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e55b6e2302cf55eb46e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18bc8df6b4ffe9e7ccee7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9ef4142805377a31dc1b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c1e17548cd9be3773e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h123959aca1e33993e7dd0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15164d2a2fd1346615e45;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h92ecc3c3f5c166330b58;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e297ffe49f579667b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c4eb6be1ca5a4c1e27cd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f8eae466e42583d75c86;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11705d782e3ca9780027e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h677bc0d6a0c65d810fba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h59b3ee78e652fb024536;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h607c2b68da69a4f071c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h89ccd9920e58f36871c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he208051bbe3bd2adc03a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h54aaa50feeee65e7447f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc9cdbd9d6486fd47174f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h163493cda7e6ef1822878;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf579968b2cba79214f64;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h178481a4dd7ffa989f3f1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1701d7fd91aa524221351;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ea4c6d17d176b639e114;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h152d01807d3578a13db58;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf87838dd990da6b549c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hac1e870ff92b12268aa0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1361bcaae040feedf96e9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha60373fe1a3f30e981a0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h964c366271cd752e0b5d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6d24b0a130db4047f9a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6f66164d799f839765ca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10541e15c2ffc5e33f4b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14993a17a5c7100ca65c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5155b3e3ef704782cdd9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11af4de76b0608c11673a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bb38d5c3d893d16abf61;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3f4a47917a787a81bb2f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h129eddaa4fd67f9f79d65;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h990d084f4b8a1cd80b17;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f6258cad1d3d313b351f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e18543d64afd23b117b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hff66e5c3a52ed8cae9a3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc22da0d6348659da080f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18b76ea1918b6db4e9628;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a2bc5605808b58c0f5a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15f4d214b62f6fc9e16e0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he81fcb2227b7c93a25c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8a20435073e6c273d10f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h32ce55954758fb26bb39;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14c5af14e5e615fe17eba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9e83e7dd240c1a0c95e3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd2050dfa6dd72ff6a26e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h176af4f3eb03268450c1a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8b68d38287c5d94475c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h95ee88493acf6c9989ec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5ba6065275cd929464d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18df9ab72a87efdeadfc8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e5615369dbd918396dee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1454c50b1c5dc180074bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha77004880393b76d4d2c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e4bd4c879ed9bea0518e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bbd765d08f8c8a6bab8e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c7f7f7b1da5ef6bbdf45;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10a647e11d1098a43a613;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h603e94def737e3042a5e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfa85a18410ffc5b1662f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc53400b2f1bfbc612902;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf5881a0b98548abdef84;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12ec29fe46f923b5dd93a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha43fb956d3141bb76e56;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he30323692c50b2a4b326;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h152cd2987ad170927113b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e498aad9d473ad7c608a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b5862c8099e8d83e34c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb14585c3cd9d7ae9a16e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h190554c80ba2ec6b2ffc1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h578af908f051abeb8069;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d9d38d22ba9db5144504;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h96e4b879f752bcefb9e2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c668c4bc955ebb0d405f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10eac55e093bc7966fa81;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e641f5f39278b8f97663;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13a9ff4dbfa0951c53869;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8dfbba8d177011f88ede;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbb508e9e6f0c2c9dcbc4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ba6e850673f6006ae1d3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1058fa16093752cb3986e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h208095b9577785869d46;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d958d7438841f31942a0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14c2255fef1ff5c4ab044;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hae8ba71303af52906dd7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f19acc5a4fe6418fbb99;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h790e1da814a177b6d847;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h368ea2cfd328e12b129a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h35bfcaa027a67609f82a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h89c793a7cb288de77034;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4a12e9d02b4eefa7aa6e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18bd46a6bdf93932d85c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h189497266cb6ed7396929;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1114744330a11fd287df4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he698e81625ea8c3d0f65;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1afc17618d274f7c97fc5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd8f4ac5b220782ecea12;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h824f4dc95161294ca117;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5c76612014b53ffca2b4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hea3772012db6d30c2c0c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h26c2c7a15552bf0648cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h157ee8d508a0189474c63;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he1c0ceba53d7614bfe98;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ae7cb8458672f801d9f5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11306b6f0f552eb8d970f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18665a1823cad6b8cd012;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17a4ae587e93f89a9300e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8843d052a0d8fb42d7bb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h93afb84d3a1c7ede995f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf13c5aa1c730cde5b6ac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h154db8fb5629a1684b04e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h103cfc9e202698ae2fd52;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1603c2b74550b098e52a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h132f2194d0a64a51373fe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcdb6db348ee50319cae7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h137254a972ac61047ce1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11fc73226bc6ea4cb07c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c733f2b41aeb8f2dd0b7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6622acfd74d1043f73e1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cd2fad7e137d59d78095;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1569955b0ecc709293eeb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1881ebf790f3163afc064;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha883a4ed17542e61fd95;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1583f593f868dbd638289;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h94a5516b8fb6a2106f94;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb0ab691fb9e0a757cfdb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e2c70bffca74ee535ec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h98dc747cc85c3b13388f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13ec76d7b11d9caccfc39;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h113d1d1f7154e162b3115;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc3e6105c946b57de1d2d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4bf6da5b00430118219c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16e323a7f4291bb829707;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d7584a040f09f4f2f19;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4b4c0c04374ff6d9ab5e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19c462eb0862c53fea345;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h32fd3bb03434c9e9716a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha9a7369aa27b48883cef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14b37d1b02fb797aee64e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h58909e90711fc68800e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19e7f95d4aec1460e53f2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3173af5549cbfd30045b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15278bb1b05a75061c6a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h302c528fc7285ed3a364;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heafa3ea58b72f2e1f031;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13538b7f8c28386bd539c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h160cd69e08e6b46cede13;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d938ccf1840b6a5556ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5876dc63b0511e543b34;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc69896eca65eea3cc7df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1daf4fca1503e82d7b6e0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hef411f8daf9673fc04df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h158065c19f238071261f7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7c941f1ebcb3eb5495c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h149b2dc6ffa00451f6978;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf69061a15ab72fe711e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h847b5a74fbe453dc922f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf16cbb74e5ebd23f65ec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h108fd5725bef1d4ebd1f6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha40fde33404840a114a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1131a307b894cec3ccf74;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h83aaaa3be0e9e53cc193;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h20b8937202e4577d25df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19783794c72c2a3fde1a6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h90eb0b32138a9f02fc34;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1de7e50c90e2c67c45616;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd9a09ebad520721d81a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf262a4c668d8be2906d3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a2bb888575c5a8f06804;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d8e429ac8b21becaaae0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9c5ca75309ef2ad73318;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10b015604886226f728cb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd100b8453a502f475f3a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h21af2281777a0497c628;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1955725d64ff425748140;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he9aac380e420cc4bcd4a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he9f81d0340db122d528a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf7c0a4559b5245cae59f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb82fbbb19091737209ae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dd6102c5e259467a8e54;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d0bc54eef726b0603654;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd50ef4d79c16a5825240;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4a35f1b2788ee9f8fd52;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1239f1b597ec280f84244;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3541a46e71453e633ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19ed1189f097e2b9e7c2d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h156946299ea5c91f9bbcb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3644476e34bf9518703d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11089ea85a5d615d926d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1584ae1dbb94d15bcf9b2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16f6843cf66836a9a04de;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'habd275e0d5945b947203;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c611e83ec6dabfedb65;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h167a953f651ab8e05af1a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c46b57cfd251f16d7542;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1011c9b2a3c10470d6777;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e4a19ce9a1a04b65553f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h102cac4df7c3f0f36fd91;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc54f8f08309876cf7d12;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h56b50caf43a8e4b329b1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h177a9c5b89bfec4af76eb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10fa82429808a21343e1c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12f214a09ced9df96d5ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fbaacc1f3372fc0cb761;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10741a7f30a8541e98485;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha5906391b81c8723b50;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14ddbdace2a210bc92d7f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15bbf7c04c9f0b038aa07;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h97b99c9f6fbbf3ce2949;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h105256d7599f78eaa9fd1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cbbf88ad9d77f0bbe2a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1085ac550ef0f660c0606;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd20412075a997c44038c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16fbcb2f6cef123ff1a9e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h143dde63846d03d207c17;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13ac8a32b224e0cc4a0b1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h175d413ad85ffe744a099;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h106ef113915afe5a3ef61;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc5a6a8a40e499f57dd6b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h908198b67b2316932713;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha6f2e827de72cfc9f6be;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h85df1e60294d95399142;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c45d806861860f2623a0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9e8629bd33975eba6556;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1511fa690423169d54b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h182452a179391a2ee433c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb9295351ab3d006cec65;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc9d9ede3796160b6fd5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4289267560e7957a7350;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e707066ea500a6608ac3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18402b1ac80f0140b292;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13bf4c0152a23bd8ff5a0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15e798228d8d21a048912;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hafd1a068bc5bbdcd1d7e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6c2371b2c07fcfa2f542;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d1ac439cf33a5836727d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbfab88f3385079674bb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b20d3581bde0b94c97bc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h54578f0f0abfe6edcc6f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ef661c8d245e2b856ff4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6cece99d90d058bc1b02;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h70c815d6347295f53602;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2f8d74b23f5956684bf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he34e78461fb57cca486b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h88321d60858fffb5322a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h176f9a71160b37afd744b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h408439bec4de778687ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b7315b4ed55da3d7d924;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hed679b22dc15ffbf60a4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7de77afa75ef7f9fdb1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6f820587218246013fd4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12bcd0085217f4c896196;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c907ecfd547c1e1c4d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d0ae23fbdeffa381f6e9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f2bff82a61f63e53c9b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1789aa4dde46f17a64dc7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h146b787e48a3e206a2dd3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hae2634b355928073bf3b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d2e973eb56c18657bc2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cd722cf2d6a001d2ab20;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12dddbc398c8b61d8e1ba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13593c77959bf6ad915ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1259b811b9aa3efac6816;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18e6f33897999623bf2ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e1907ee0e126359c086c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eef19a13174cfff3d624;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2b17b997470e96cb0b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a7752b303bbf9f79e46;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdb01363481b3ae50ae24;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1201baec5278a4e539256;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h100680681a7a8ab263974;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13955f907beb4877c6b88;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h94572fd5281ad0aec96a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h144c75f34cdc17f418357;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb3cca5ca6f402eafd48c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b0edd1b426b26298731;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1de5eb024c564bcc252bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7990ee1bdd36c3e7b971;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h33d7f5a52332a7cdc703;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f080b8017537a2bd55a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e94b60cc1ccac211551;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h174abec52dc9527db7c6d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10099fdb4a05f8f1e3b10;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h53b130765b938849c080;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h196b56becab40b4c5a24e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf77fb30bd6f5bbf4438d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18afde94d97d00fd9e335;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1066664bb6c324598ab4a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1102f388041578b0352e2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3172ca2a355efc58c108;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ddd263cc024e7ca6b074;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd3974d0fb088f23008ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haccd2222a55b4b815df5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e7a7fd88c835ddb274d0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19bc6a2aa2bc2d7f6c01f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16d96b7abce991e576a10;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfea5d7b4e9c4ff72eb9b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8f52fcfadb012176d2e0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6e18caebd2eb39fb7dda;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16de21157e92cf7d00f93;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hae13be6567e80de52f7b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b313d2488187e7d3ae00;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a337ffbf0a56b7c67937;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h100a572ecf0506d67b328;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfb92dd38709366161e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19eb8c9b33fe4854aeb5c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12174438fdd466a7a391c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14363ce082db6549bed6d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f9b08db579c9ebb0104;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15be833400254176ea6d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ed0588bfc3cf8484faf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1864032c8b6c39c79d6dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17dde13dd1aabc95f2434;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc997ca6c4f1c8a559084;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha9eec4d4ff062cd95d3a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3dac9b363d5d4ac38cbc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8c3ac0743215dfbbee20;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8e7da0b35f6678e45929;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hec8fd13feea6f0162483;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h505768ffdcbbb6a632f1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5226277782585b7a4332;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6bbe0c40cacf3bd05520;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h545bc28c1dd68aa3ff56;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd4f04c73ab86a0345b2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13b62b07151b306e6a5c9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h84ff721b2667e0663f7c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h459852c1d23b44f1534c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8880f46c9f249c031d5d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18219151e41270cdc8452;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hffefa9c7dde69c1e35bc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h689f474b4f55bf8f9f49;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc221e32066925692be8b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c5929e2552d311a7541;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h69b2f892768747fb0b67;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc91b67f6a890a4798a67;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb6ad47eb3b36514538f6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha0040da28ebe4541f1fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18c90598c78e008bd8551;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7189a9f9fc345b29f426;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c12d86031dd943e0233d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11418ac6ef419bd38d359;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd7cba183d6dbed530b9a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f629f2e371f9b1ece3de;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ed8e37f6c4abbf9b5f87;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d7ca6e3921afb453606f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e73643273daf26a6e99c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f09debe862f4ab0a6a0f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha66d637597b3b4fd1031;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h82a2df1621c2aedcbb32;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ef476110ab4b5aa99b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f600a75e5b18cd27869d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a3bc243a0ff1ecb5a2b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be6e35e24c83c280e5bc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h49e3183a28e2aabc565d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h393ae9b81853b5fd948e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15d28e821659a8956263b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he9a9476bfe2530a3cca0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd030600273338cea753c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5e1fe23676c4d72ce1b6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1adde7ed5c2d5c6cbbb89;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h198659258b4e9b6a411af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b30d3dcdbbb115605564;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h28806ed399bc1af6784e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hda05d1e3e166028c7f37;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f917c5b5814fcf50362e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbd9bf2c768f83e3febcb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f73b78f1fbad38bfa73;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c600a41e16589c9c26d4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c33c690f5f6153cde9c2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h31784a2e2e6f628be106;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h418415fb7392d549a927;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14e958865ee8b70db5eb4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13a6fa49071b91bbfa100;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4272c11676df0167f6f5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1619fe72d445ae301cb90;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha5cbfa85d389f6b25198;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10e0e4471460c0b63e0c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a083e37f76e58d42daff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h32ef86cc24c37dbafba0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h26884a966a3b393d7ad8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8660034e30d56a7bf23;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd176f85fc8fd0320aab5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e9a29afcec8a2090280d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e014c317206aaf0dbe64;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f61a9cc92b99d708b372;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cdec944230d33a09143e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he0b69222f96106efde8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd285e897c66f9988a79c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e1afc29eea70dbb736b7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18f255bd1b7103ef6076b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c81e41fa3ae73edc4473;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h83effa9ec479cec62b84;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e1b470fa6e47f4dd7d89;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1603c7436daf4fde32aa1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf497829a8ba66c88e9af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hde47793b7d9d12b2ef1b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha8934043e5a947f14e7e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e93bce95a7c4950f0355;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h101359bb8d81776289107;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18d312461409c664cf701;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfea494e56a5c72eb7083;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c4a3d57f435bb4ae2112;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1461704d34226e7128c55;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h135de30ae93718d97544f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfd6ccab7ad04a6866d2a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2baecc832d303bb80c15;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf6db34439b6e3d0f9408;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbe998d2ae65b92a95280;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ce529e71ec37db8c470f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cbcfee9eec26e6857d6a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha37e3a7e5c04787af9d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h60a1445ebbae98e0063e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b076620ce08355b271d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h609109dcbaeaf8a8fbda;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha7c2b3e6589a7faaf735;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc212af1271fd172bdcfa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he373c2ed480e0dad27ba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h143795875e4ef6d7a9757;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb0583361e9665b8b3bbf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he77272144276d481b6fe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h150ea7e50fc5613ff7b68;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a0548f221f58861d513;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h46569181a973311feb97;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9188db22d86d69c3f266;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h354675b8abde7e77723a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13e134d91fec539b3d532;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf087cbf42a8fa1722411;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h112d3e9ff51124aa3f820;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1096b1dc2b665cdf9eefd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ab547d6a6641e8710e78;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h146534223b9f12a130343;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd5b3b11e51163aaee472;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19312665a34d0cb78f10c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf211fedb4cbca92592a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he7fe7fdca6ea53f4b3ab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h181e40c2cd29518506dff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd56fadac6f37a0edf5c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1035c721c54063d658145;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6b0537c199afe8beb1c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd787a8d92fc9f8038ce5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h137c92ab982d45295c871;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf52b551b39f8f115c197;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15b2d9330bfc1a9c3f490;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1050246751f7e1211b55b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a08d37d6e2a3443cc9a3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h24fb5a0d67688439b808;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1945ad2b8739bcf135250;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcdcc6a91cb761d5b525;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h28f6297d205978dcfdb7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h35ae86c7e13bee9a8e70;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb5f838f8feb573d01eee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ec590d96afed5c03d0cd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he450cda28c7ad0a90cdb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1370fc8776b8411d3b0cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha348c5e829284e2ba697;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1626b3fd1d5e0c8a9d07a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18cf58766bb0bc66ed984;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16da46e55582690db3a2f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1616338eb0cfd252109d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb202a4aef4d6adadb3f6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bcff62c47e7122685737;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f40e5c0fc997eb493484;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c59ee82f27476d80f9c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h128a1e56e2c06cc12016d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h131efb2230a77d0c3a2a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h39c6181ff6b217af27f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdef549c2dade54e5757a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fb0f7be3b769c11fa76d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h81a5d2e58a1d12ae8f57;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc91b9bcf02d1031ae8a6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h179541d3d2aae4ad8807;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h953a1cb72c5fa7058f61;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f823176109733659d3bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c0b260cd87893c3885a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbb1b0dc942b22621bc0a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16d44fe71d7a39e668da6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h137e243a0ceed85c13e86;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c81eb54a6785ec816e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha2547268550647a021f6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h178705ddd30bb0163cb1c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc53884aa1ca02896cd83;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ac497151efee04a5b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h35de5ad5191c99a437a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd5102ea1dbe5bec95c47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h94e4b8578631e15f18f0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfcd27c0f19674fbd6d70;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a1203778d0c9f4f9da68;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h144c2347f4ff21f1669ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h668fb23bebfca0f7092c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f7cb27f349cc89f0107;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e2415f2047c794dd2e6b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8b10319506bf21122bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdd1ddf1180b3fea01d58;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h197346f86f7303516d8d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1580bf2106bba4a76ac6b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14404fe92f211a37c3e54;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb1acd744721be52c06c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d9e11d9e1b66570150ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h66046587b5ee380df983;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h81674b4219518ccfadd7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h187f0bba3d10f094bc39b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1639924bda554e8509f73;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b8a9d53d236a71e64ad6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h96f62edb2dd84da792ba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hda858a53906885e7544a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h35a966b777d897bb354;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19f3e43672e6d62ed1f88;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e7beaad17c8d317bc391;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d92d91a139f049dfd2a0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12e95abb9fd016a43ba30;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ce3494b9193c9407ab0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h846ef3807176f73e6339;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h83415784b50cfa701f2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19621c5b12cacd1dacb96;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h384fcbd243a52b5e19c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17938b4b831ca930420fa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13123dd7433dcc1ba2f9e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb5d5cd6cfe8f6cedde81;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13b57481689771bedd395;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfc3050b56b15a24cef69;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf5a331de8bebf557fc41;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8e6d18368c0f75b453b9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2644424286741418ad9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cdb60d62d2a0dcae6ac7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c1366caedeffd8c6496f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d19465c9f71311c1037b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1779d1b8e581f10d62066;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a2bed934fee7638e1c0d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ac7a4d402fa2636490b9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h158b91bbb806e50ec7059;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13fe741e29f15c1324396;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cd8a63b67efdb4cb6482;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h38c27f777ffeb37d1c90;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heaf0ac4468f51069a64f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a43aba55f9b68e1c66ce;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7839dcdd0576a94da0ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9af33a754357dcf4ed07;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1048a75ee79c89deb422d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9e8be76fb011d09bb37b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d66044afdeda8c2a3a4d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h70cdbbef2214202c55cd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c25080c01a649a06d492;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd788580a670d663f24bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b19bec97c9835661e2b2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1458a1351a6d646298c67;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e997f687951e46bd2115;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h177e2a2019186ea477a65;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c701e65fbf198a776ee1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c7cb8d10008b90fa671d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f20a7891a0623cc3b168;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hab75aff8cb18ddd95679;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18b3ae3389514ab8c4308;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b36e066c1dc8c2c1cf99;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ed2e5ba1abe13fa35202;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h161de6c5be1135ee7c663;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1716d04c6c790534658e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9affe53baf6ce501e052;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbb6553ea999f0c29879b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha79a504acd2da00a8892;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc34c0c63df4622fb8972;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf4af285f8ebd2b155399;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h124825c7bf5e0537ac49d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1305a8906372c5f7c14ce;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f4eee52c31ec36ddc4d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16776331404e766dced0e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6d022b5a06a51447af7c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d0a3a8d2c174ccd71d04;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h23d029c44452ebbcfee7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h51a123ec6690357651f1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdd2ac09aa01879b58975;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbaef4e35298daabd2df0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h106f728fe1a5af75a56d9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ff55c8cb5a2ad86cf9c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15ee6bd62801b63144d3c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h150cab39ba33eca294586;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h89e512aa3c5b09083480;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb658eb0eec26de5dfc5e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h175e6e89424f37e32b8e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he3d3216db7a42250a51d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bcac3d3fcbf1f8107a3d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a269d33fde731b8e4607;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17cfb42df24a198f8def5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcdc4a6b7112978ef0047;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb340f558f218475cfed4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4209547b4c5566cb66c1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16800b2ed9a7777229242;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fe22bca37837a97017a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hba7b870111e3be0e24b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1703e8fb91ab6b78b6746;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h155c7c0a8cf89db40d335;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h59ee352710120269b439;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10c37aa0cc0bc14bb5a89;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cafaa652715a877f2b0c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11d4994ee77d5ad5e727d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3da57031a3bbae1d0d0c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd09561f3f0ad635aab98;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h107eaa2f439128acb2414;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13a18af993fe5016f766f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7b2888e74569be6f7d5c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb09c7997c056d3003e59;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf896b157c3a3a82a0887;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12e883c49730cb66f5b46;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7ee39ca38380452617e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf512e859aa8ceeb72e44;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4aff70a03d01e3d31635;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h41b58124f86377175067;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hea55d7debf0cadf98fdd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cd52eb582333069f2a7e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h234e7e79ef17e6f07eda;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1455ed76fab41b24eb6a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11de7cc345aa246e61fc0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h68a348d901f0c39db824;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19ef8decf6e1e60804983;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf3e03034909e342bb4e1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h28c3a44b399b48b700e4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h104d7268f37d01eccff41;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e2be0c078a09d5fb1068;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3fdac4d7409b87fe3bc2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h156a5f2909f9681094249;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h109e730f5578b704111fa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c97b300c8127320a6d1d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ea630862363642a7065f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc9dceb7e2dfd54c26306;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18bc026345fd170759dfc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e12d682d6f7289f1c7e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbfa7aab8af51ac6a500c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ec22004e67387438bf8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1373359b6fa6a91793bfd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a71a0f7101ca754dde7b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10438afebc696e750e4cb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbfa3def51c1553ad9a31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c1782e1f9149311fb5f7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1188d65617289be39cc72;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18afa2242d109226af4c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ec4678adc6d53d2ffe4a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1930660c7ed7c0d942a82;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2e4b133fddefe4abec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b644a4e182d0db2193b2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbd4dc1c482cf06133689;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a72ec8782973dc8c760;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11866cf06d0008570f08f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1142cba11ed3f7ea36b49;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8139b0eebefa358de95a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15be8a375c99a41e0f355;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd337a3bdb97976eb3f5b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d1cbe0f46f71c735fea7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f409aa0557e0786a470;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h132892104d5360e8b6141;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h109303e0894d404714fa9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7354bf03c8fb3d90dcc8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b1acd9e3cda5fbcdc767;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdad94166c8a353dd916e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1020a2543f353012c55e3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7fcf11ca5b36a8f287cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h85a33378f3f2d3487dd2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d45f94afa3bae230c7d9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hee795c9f9566a1076773;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c372e4da7ecea5eb6eb0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6a086cfa0b9a66fcfdbd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc4cd832d8b26429dfa4a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcfceea7fdb147b9df341;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6d355c53249201c837a2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h140c69af7a87e65cdbe52;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdde9ebee3a413ef6a245;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h93491c50d6aa74b7a80a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h180265a12b92fb9f0ed77;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb319a171ecbbb1f9af0a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he90754d00044d41b64e9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3bac1a5ab972bb4ce1a9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16b752d6504e15d7e5040;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18426ecfecdb80bbab471;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1be6af4e71c0dbc98bd1a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a1e9dbc606ae84ea3035;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf1a49fa5daeb43eb0c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a9f03b773d386e42699b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ea7d53f20e3f90c78d89;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1955ef94fa25ad9c0ea5e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h83186851f3e28026c3e9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15638048dd17a9bb90e85;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h52feda2f1f653287ae72;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11c16b2bb497994c10e39;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb96a625f2bb5425fc331;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1677258aa8041650e2116;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11f97da5c9799b86fdca9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he52c5f3ffbadd8c4ac14;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19e8112919a418e2b789d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h179709d8f741b4ce4a67;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h28968f87a08eb18c236b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bfb395f5dd2656088d31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1005610abc5450d0ed161;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd74247d43970b663b03;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h162f1dda4905dc6f0ac9a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1539794ae5503640db5a3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h53ed0d52c848334d0831;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1045fe10cf3b63899fe2e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h56a32ea2a4e89ac8a5bc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1833e9d49358f490df826;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18adbe422c2d61709c044;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h95c776efc3485710c7d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9ec838230e64010d174;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h117225a5f7c603e539eea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1efb6981596ab818008a6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1821f2144b0925eaa1fe8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h584d0ee1517ec4840509;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3c086b3fc404f98eee48;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c7bf6e6fb9cd3b14878c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc626a8c4a4006e1aa073;
        #1
        $finish();
    end
endmodule
