module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68,
        output wire [0:0] dst69,
        output wire [0:0] dst70);
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    reg [127:0] src12;
    reg [127:0] src13;
    reg [127:0] src14;
    reg [127:0] src15;
    reg [127:0] src16;
    reg [127:0] src17;
    reg [127:0] src18;
    reg [127:0] src19;
    reg [127:0] src20;
    reg [127:0] src21;
    reg [127:0] src22;
    reg [127:0] src23;
    reg [127:0] src24;
    reg [127:0] src25;
    reg [127:0] src26;
    reg [127:0] src27;
    reg [127:0] src28;
    reg [127:0] src29;
    reg [127:0] src30;
    reg [127:0] src31;
    reg [127:0] src32;
    reg [127:0] src33;
    reg [127:0] src34;
    reg [127:0] src35;
    reg [127:0] src36;
    reg [127:0] src37;
    reg [127:0] src38;
    reg [127:0] src39;
    reg [127:0] src40;
    reg [127:0] src41;
    reg [127:0] src42;
    reg [127:0] src43;
    reg [127:0] src44;
    reg [127:0] src45;
    reg [127:0] src46;
    reg [127:0] src47;
    reg [127:0] src48;
    reg [127:0] src49;
    reg [127:0] src50;
    reg [127:0] src51;
    reg [127:0] src52;
    reg [127:0] src53;
    reg [127:0] src54;
    reg [127:0] src55;
    reg [127:0] src56;
    reg [127:0] src57;
    reg [127:0] src58;
    reg [127:0] src59;
    reg [127:0] src60;
    reg [127:0] src61;
    reg [127:0] src62;
    reg [127:0] src63;
    compressor_CLA128_64 compressor_CLA128_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68),
            .dst69(dst69),
            .dst70(dst70));
    initial begin
        src0 <= 128'h0;
        src1 <= 128'h0;
        src2 <= 128'h0;
        src3 <= 128'h0;
        src4 <= 128'h0;
        src5 <= 128'h0;
        src6 <= 128'h0;
        src7 <= 128'h0;
        src8 <= 128'h0;
        src9 <= 128'h0;
        src10 <= 128'h0;
        src11 <= 128'h0;
        src12 <= 128'h0;
        src13 <= 128'h0;
        src14 <= 128'h0;
        src15 <= 128'h0;
        src16 <= 128'h0;
        src17 <= 128'h0;
        src18 <= 128'h0;
        src19 <= 128'h0;
        src20 <= 128'h0;
        src21 <= 128'h0;
        src22 <= 128'h0;
        src23 <= 128'h0;
        src24 <= 128'h0;
        src25 <= 128'h0;
        src26 <= 128'h0;
        src27 <= 128'h0;
        src28 <= 128'h0;
        src29 <= 128'h0;
        src30 <= 128'h0;
        src31 <= 128'h0;
        src32 <= 128'h0;
        src33 <= 128'h0;
        src34 <= 128'h0;
        src35 <= 128'h0;
        src36 <= 128'h0;
        src37 <= 128'h0;
        src38 <= 128'h0;
        src39 <= 128'h0;
        src40 <= 128'h0;
        src41 <= 128'h0;
        src42 <= 128'h0;
        src43 <= 128'h0;
        src44 <= 128'h0;
        src45 <= 128'h0;
        src46 <= 128'h0;
        src47 <= 128'h0;
        src48 <= 128'h0;
        src49 <= 128'h0;
        src50 <= 128'h0;
        src51 <= 128'h0;
        src52 <= 128'h0;
        src53 <= 128'h0;
        src54 <= 128'h0;
        src55 <= 128'h0;
        src56 <= 128'h0;
        src57 <= 128'h0;
        src58 <= 128'h0;
        src59 <= 128'h0;
        src60 <= 128'h0;
        src61 <= 128'h0;
        src62 <= 128'h0;
        src63 <= 128'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor_CLA128_64(
    input [127:0]src0,
    input [127:0]src1,
    input [127:0]src2,
    input [127:0]src3,
    input [127:0]src4,
    input [127:0]src5,
    input [127:0]src6,
    input [127:0]src7,
    input [127:0]src8,
    input [127:0]src9,
    input [127:0]src10,
    input [127:0]src11,
    input [127:0]src12,
    input [127:0]src13,
    input [127:0]src14,
    input [127:0]src15,
    input [127:0]src16,
    input [127:0]src17,
    input [127:0]src18,
    input [127:0]src19,
    input [127:0]src20,
    input [127:0]src21,
    input [127:0]src22,
    input [127:0]src23,
    input [127:0]src24,
    input [127:0]src25,
    input [127:0]src26,
    input [127:0]src27,
    input [127:0]src28,
    input [127:0]src29,
    input [127:0]src30,
    input [127:0]src31,
    input [127:0]src32,
    input [127:0]src33,
    input [127:0]src34,
    input [127:0]src35,
    input [127:0]src36,
    input [127:0]src37,
    input [127:0]src38,
    input [127:0]src39,
    input [127:0]src40,
    input [127:0]src41,
    input [127:0]src42,
    input [127:0]src43,
    input [127:0]src44,
    input [127:0]src45,
    input [127:0]src46,
    input [127:0]src47,
    input [127:0]src48,
    input [127:0]src49,
    input [127:0]src50,
    input [127:0]src51,
    input [127:0]src52,
    input [127:0]src53,
    input [127:0]src54,
    input [127:0]src55,
    input [127:0]src56,
    input [127:0]src57,
    input [127:0]src58,
    input [127:0]src59,
    input [127:0]src60,
    input [127:0]src61,
    input [127:0]src62,
    input [127:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68,
    output dst69,
    output dst70);

    wire [0:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [0:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [1:0] comp_out62;
    wire [0:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [1:0] comp_out67;
    wire [1:0] comp_out68;
    wire [0:0] comp_out69;
    wire [1:0] comp_out70;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68),
        .dst69(comp_out69),
        .dst70(comp_out70)
    );
    LookAheadCarryUnit256 LCU256(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out70[0], comp_out69[0], comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out70[1], 1'h0, comp_out68[1], comp_out67[1], comp_out66[1], comp_out65[1], comp_out64[1], 1'h0, comp_out62[1], comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], 1'h0, comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], 1'h0}),
        .dst({dst70, dst69, dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [127:0] src0,
      input wire [127:0] src1,
      input wire [127:0] src2,
      input wire [127:0] src3,
      input wire [127:0] src4,
      input wire [127:0] src5,
      input wire [127:0] src6,
      input wire [127:0] src7,
      input wire [127:0] src8,
      input wire [127:0] src9,
      input wire [127:0] src10,
      input wire [127:0] src11,
      input wire [127:0] src12,
      input wire [127:0] src13,
      input wire [127:0] src14,
      input wire [127:0] src15,
      input wire [127:0] src16,
      input wire [127:0] src17,
      input wire [127:0] src18,
      input wire [127:0] src19,
      input wire [127:0] src20,
      input wire [127:0] src21,
      input wire [127:0] src22,
      input wire [127:0] src23,
      input wire [127:0] src24,
      input wire [127:0] src25,
      input wire [127:0] src26,
      input wire [127:0] src27,
      input wire [127:0] src28,
      input wire [127:0] src29,
      input wire [127:0] src30,
      input wire [127:0] src31,
      input wire [127:0] src32,
      input wire [127:0] src33,
      input wire [127:0] src34,
      input wire [127:0] src35,
      input wire [127:0] src36,
      input wire [127:0] src37,
      input wire [127:0] src38,
      input wire [127:0] src39,
      input wire [127:0] src40,
      input wire [127:0] src41,
      input wire [127:0] src42,
      input wire [127:0] src43,
      input wire [127:0] src44,
      input wire [127:0] src45,
      input wire [127:0] src46,
      input wire [127:0] src47,
      input wire [127:0] src48,
      input wire [127:0] src49,
      input wire [127:0] src50,
      input wire [127:0] src51,
      input wire [127:0] src52,
      input wire [127:0] src53,
      input wire [127:0] src54,
      input wire [127:0] src55,
      input wire [127:0] src56,
      input wire [127:0] src57,
      input wire [127:0] src58,
      input wire [127:0] src59,
      input wire [127:0] src60,
      input wire [127:0] src61,
      input wire [127:0] src62,
      input wire [127:0] src63,
      output wire [0:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [0:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [1:0] dst62,
      output wire [0:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [1:0] dst68,
      output wire [0:0] dst69,
      output wire [1:0] dst70);

   wire [127:0] stage0_0;
   wire [127:0] stage0_1;
   wire [127:0] stage0_2;
   wire [127:0] stage0_3;
   wire [127:0] stage0_4;
   wire [127:0] stage0_5;
   wire [127:0] stage0_6;
   wire [127:0] stage0_7;
   wire [127:0] stage0_8;
   wire [127:0] stage0_9;
   wire [127:0] stage0_10;
   wire [127:0] stage0_11;
   wire [127:0] stage0_12;
   wire [127:0] stage0_13;
   wire [127:0] stage0_14;
   wire [127:0] stage0_15;
   wire [127:0] stage0_16;
   wire [127:0] stage0_17;
   wire [127:0] stage0_18;
   wire [127:0] stage0_19;
   wire [127:0] stage0_20;
   wire [127:0] stage0_21;
   wire [127:0] stage0_22;
   wire [127:0] stage0_23;
   wire [127:0] stage0_24;
   wire [127:0] stage0_25;
   wire [127:0] stage0_26;
   wire [127:0] stage0_27;
   wire [127:0] stage0_28;
   wire [127:0] stage0_29;
   wire [127:0] stage0_30;
   wire [127:0] stage0_31;
   wire [127:0] stage0_32;
   wire [127:0] stage0_33;
   wire [127:0] stage0_34;
   wire [127:0] stage0_35;
   wire [127:0] stage0_36;
   wire [127:0] stage0_37;
   wire [127:0] stage0_38;
   wire [127:0] stage0_39;
   wire [127:0] stage0_40;
   wire [127:0] stage0_41;
   wire [127:0] stage0_42;
   wire [127:0] stage0_43;
   wire [127:0] stage0_44;
   wire [127:0] stage0_45;
   wire [127:0] stage0_46;
   wire [127:0] stage0_47;
   wire [127:0] stage0_48;
   wire [127:0] stage0_49;
   wire [127:0] stage0_50;
   wire [127:0] stage0_51;
   wire [127:0] stage0_52;
   wire [127:0] stage0_53;
   wire [127:0] stage0_54;
   wire [127:0] stage0_55;
   wire [127:0] stage0_56;
   wire [127:0] stage0_57;
   wire [127:0] stage0_58;
   wire [127:0] stage0_59;
   wire [127:0] stage0_60;
   wire [127:0] stage0_61;
   wire [127:0] stage0_62;
   wire [127:0] stage0_63;
   wire [29:0] stage1_0;
   wire [32:0] stage1_1;
   wire [46:0] stage1_2;
   wire [66:0] stage1_3;
   wire [65:0] stage1_4;
   wire [51:0] stage1_5;
   wire [88:0] stage1_6;
   wire [70:0] stage1_7;
   wire [65:0] stage1_8;
   wire [60:0] stage1_9;
   wire [40:0] stage1_10;
   wire [63:0] stage1_11;
   wire [55:0] stage1_12;
   wire [53:0] stage1_13;
   wire [65:0] stage1_14;
   wire [67:0] stage1_15;
   wire [88:0] stage1_16;
   wire [66:0] stage1_17;
   wire [41:0] stage1_18;
   wire [54:0] stage1_19;
   wire [71:0] stage1_20;
   wire [54:0] stage1_21;
   wire [70:0] stage1_22;
   wire [53:0] stage1_23;
   wire [61:0] stage1_24;
   wire [60:0] stage1_25;
   wire [83:0] stage1_26;
   wire [55:0] stage1_27;
   wire [47:0] stage1_28;
   wire [79:0] stage1_29;
   wire [71:0] stage1_30;
   wire [59:0] stage1_31;
   wire [82:0] stage1_32;
   wire [62:0] stage1_33;
   wire [67:0] stage1_34;
   wire [47:0] stage1_35;
   wire [60:0] stage1_36;
   wire [96:0] stage1_37;
   wire [43:0] stage1_38;
   wire [92:0] stage1_39;
   wire [62:0] stage1_40;
   wire [39:0] stage1_41;
   wire [50:0] stage1_42;
   wire [78:0] stage1_43;
   wire [49:0] stage1_44;
   wire [57:0] stage1_45;
   wire [79:0] stage1_46;
   wire [69:0] stage1_47;
   wire [45:0] stage1_48;
   wire [50:0] stage1_49;
   wire [70:0] stage1_50;
   wire [47:0] stage1_51;
   wire [60:0] stage1_52;
   wire [61:0] stage1_53;
   wire [51:0] stage1_54;
   wire [67:0] stage1_55;
   wire [56:0] stage1_56;
   wire [57:0] stage1_57;
   wire [59:0] stage1_58;
   wire [55:0] stage1_59;
   wire [52:0] stage1_60;
   wire [58:0] stage1_61;
   wire [97:0] stage1_62;
   wire [52:0] stage1_63;
   wire [29:0] stage1_64;
   wire [17:0] stage1_65;
   wire [19:0] stage2_0;
   wire [12:0] stage2_1;
   wire [24:0] stage2_2;
   wire [27:0] stage2_3;
   wire [25:0] stage2_4;
   wire [28:0] stage2_5;
   wire [25:0] stage2_6;
   wire [38:0] stage2_7;
   wire [31:0] stage2_8;
   wire [41:0] stage2_9;
   wire [30:0] stage2_10;
   wire [21:0] stage2_11;
   wire [27:0] stage2_12;
   wire [16:0] stage2_13;
   wire [38:0] stage2_14;
   wire [30:0] stage2_15;
   wire [23:0] stage2_16;
   wire [33:0] stage2_17;
   wire [30:0] stage2_18;
   wire [26:0] stage2_19;
   wire [33:0] stage2_20;
   wire [21:0] stage2_21;
   wire [34:0] stage2_22;
   wire [27:0] stage2_23;
   wire [27:0] stage2_24;
   wire [31:0] stage2_25;
   wire [26:0] stage2_26;
   wire [32:0] stage2_27;
   wire [26:0] stage2_28;
   wire [20:0] stage2_29;
   wire [51:0] stage2_30;
   wire [27:0] stage2_31;
   wire [24:0] stage2_32;
   wire [28:0] stage2_33;
   wire [31:0] stage2_34;
   wire [29:0] stage2_35;
   wire [32:0] stage2_36;
   wire [36:0] stage2_37;
   wire [35:0] stage2_38;
   wire [21:0] stage2_39;
   wire [34:0] stage2_40;
   wire [31:0] stage2_41;
   wire [17:0] stage2_42;
   wire [20:0] stage2_43;
   wire [29:0] stage2_44;
   wire [34:0] stage2_45;
   wire [22:0] stage2_46;
   wire [35:0] stage2_47;
   wire [30:0] stage2_48;
   wire [15:0] stage2_49;
   wire [32:0] stage2_50;
   wire [30:0] stage2_51;
   wire [17:0] stage2_52;
   wire [38:0] stage2_53;
   wire [28:0] stage2_54;
   wire [19:0] stage2_55;
   wire [26:0] stage2_56;
   wire [32:0] stage2_57;
   wire [23:0] stage2_58;
   wire [34:0] stage2_59;
   wire [21:0] stage2_60;
   wire [28:0] stage2_61;
   wire [37:0] stage2_62;
   wire [37:0] stage2_63;
   wire [25:0] stage2_64;
   wire [17:0] stage2_65;
   wire [5:0] stage2_66;
   wire [1:0] stage2_67;
   wire [4:0] stage3_0;
   wire [7:0] stage3_1;
   wire [5:0] stage3_2;
   wire [21:0] stage3_3;
   wire [11:0] stage3_4;
   wire [23:0] stage3_5;
   wire [9:0] stage3_6;
   wire [11:0] stage3_7;
   wire [15:0] stage3_8;
   wire [19:0] stage3_9;
   wire [11:0] stage3_10;
   wire [12:0] stage3_11;
   wire [13:0] stage3_12;
   wire [11:0] stage3_13;
   wire [9:0] stage3_14;
   wire [25:0] stage3_15;
   wire [11:0] stage3_16;
   wire [11:0] stage3_17;
   wire [12:0] stage3_18;
   wire [15:0] stage3_19;
   wire [13:0] stage3_20;
   wire [17:0] stage3_21;
   wire [8:0] stage3_22;
   wire [12:0] stage3_23;
   wire [15:0] stage3_24;
   wire [19:0] stage3_25;
   wire [12:0] stage3_26;
   wire [13:0] stage3_27;
   wire [16:0] stage3_28;
   wire [7:0] stage3_29;
   wire [14:0] stage3_30;
   wire [19:0] stage3_31;
   wire [11:0] stage3_32;
   wire [11:0] stage3_33;
   wire [17:0] stage3_34;
   wire [9:0] stage3_35;
   wire [14:0] stage3_36;
   wire [14:0] stage3_37;
   wire [12:0] stage3_38;
   wire [13:0] stage3_39;
   wire [17:0] stage3_40;
   wire [11:0] stage3_41;
   wire [19:0] stage3_42;
   wire [9:0] stage3_43;
   wire [7:0] stage3_44;
   wire [14:0] stage3_45;
   wire [11:0] stage3_46;
   wire [10:0] stage3_47;
   wire [18:0] stage3_48;
   wire [11:0] stage3_49;
   wire [6:0] stage3_50;
   wire [12:0] stage3_51;
   wire [19:0] stage3_52;
   wire [8:0] stage3_53;
   wire [23:0] stage3_54;
   wire [11:0] stage3_55;
   wire [7:0] stage3_56;
   wire [11:0] stage3_57;
   wire [11:0] stage3_58;
   wire [13:0] stage3_59;
   wire [13:0] stage3_60;
   wire [20:0] stage3_61;
   wire [15:0] stage3_62;
   wire [17:0] stage3_63;
   wire [12:0] stage3_64;
   wire [11:0] stage3_65;
   wire [6:0] stage3_66;
   wire [6:0] stage3_67;
   wire [0:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [9:0] stage4_3;
   wire [13:0] stage4_4;
   wire [8:0] stage4_5;
   wire [8:0] stage4_6;
   wire [6:0] stage4_7;
   wire [5:0] stage4_8;
   wire [6:0] stage4_9;
   wire [10:0] stage4_10;
   wire [5:0] stage4_11;
   wire [5:0] stage4_12;
   wire [4:0] stage4_13;
   wire [5:0] stage4_14;
   wire [7:0] stage4_15;
   wire [6:0] stage4_16;
   wire [7:0] stage4_17;
   wire [5:0] stage4_18;
   wire [6:0] stage4_19;
   wire [10:0] stage4_20;
   wire [3:0] stage4_21;
   wire [4:0] stage4_22;
   wire [5:0] stage4_23;
   wire [10:0] stage4_24;
   wire [7:0] stage4_25;
   wire [10:0] stage4_26;
   wire [5:0] stage4_27;
   wire [5:0] stage4_28;
   wire [9:0] stage4_29;
   wire [3:0] stage4_30;
   wire [6:0] stage4_31;
   wire [6:0] stage4_32;
   wire [5:0] stage4_33;
   wire [5:0] stage4_34;
   wire [5:0] stage4_35;
   wire [6:0] stage4_36;
   wire [6:0] stage4_37;
   wire [5:0] stage4_38;
   wire [7:0] stage4_39;
   wire [11:0] stage4_40;
   wire [10:0] stage4_41;
   wire [5:0] stage4_42;
   wire [4:0] stage4_43;
   wire [5:0] stage4_44;
   wire [5:0] stage4_45;
   wire [5:0] stage4_46;
   wire [6:0] stage4_47;
   wire [4:0] stage4_48;
   wire [5:0] stage4_49;
   wire [6:0] stage4_50;
   wire [2:0] stage4_51;
   wire [16:0] stage4_52;
   wire [5:0] stage4_53;
   wire [11:0] stage4_54;
   wire [3:0] stage4_55;
   wire [7:0] stage4_56;
   wire [5:0] stage4_57;
   wire [3:0] stage4_58;
   wire [5:0] stage4_59;
   wire [5:0] stage4_60;
   wire [9:0] stage4_61;
   wire [5:0] stage4_62;
   wire [8:0] stage4_63;
   wire [8:0] stage4_64;
   wire [4:0] stage4_65;
   wire [4:0] stage4_66;
   wire [3:0] stage4_67;
   wire [1:0] stage4_68;
   wire [0:0] stage4_69;
   wire [0:0] stage5_0;
   wire [1:0] stage5_1;
   wire [1:0] stage5_2;
   wire [3:0] stage5_3;
   wire [4:0] stage5_4;
   wire [3:0] stage5_5;
   wire [3:0] stage5_6;
   wire [2:0] stage5_7;
   wire [3:0] stage5_8;
   wire [3:0] stage5_9;
   wire [6:0] stage5_10;
   wire [1:0] stage5_11;
   wire [5:0] stage5_12;
   wire [4:0] stage5_13;
   wire [0:0] stage5_14;
   wire [8:0] stage5_15;
   wire [3:0] stage5_16;
   wire [2:0] stage5_17;
   wire [1:0] stage5_18;
   wire [2:0] stage5_19;
   wire [8:0] stage5_20;
   wire [4:0] stage5_21;
   wire [3:0] stage5_22;
   wire [0:0] stage5_23;
   wire [5:0] stage5_24;
   wire [2:0] stage5_25;
   wire [3:0] stage5_26;
   wire [7:0] stage5_27;
   wire [1:0] stage5_28;
   wire [5:0] stage5_29;
   wire [3:0] stage5_30;
   wire [1:0] stage5_31;
   wire [2:0] stage5_32;
   wire [2:0] stage5_33;
   wire [7:0] stage5_34;
   wire [0:0] stage5_35;
   wire [1:0] stage5_36;
   wire [2:0] stage5_37;
   wire [3:0] stage5_38;
   wire [4:0] stage5_39;
   wire [2:0] stage5_40;
   wire [3:0] stage5_41;
   wire [3:0] stage5_42;
   wire [3:0] stage5_43;
   wire [3:0] stage5_44;
   wire [1:0] stage5_45;
   wire [1:0] stage5_46;
   wire [4:0] stage5_47;
   wire [5:0] stage5_48;
   wire [0:0] stage5_49;
   wire [1:0] stage5_50;
   wire [2:0] stage5_51;
   wire [6:0] stage5_52;
   wire [3:0] stage5_53;
   wire [2:0] stage5_54;
   wire [3:0] stage5_55;
   wire [5:0] stage5_56;
   wire [1:0] stage5_57;
   wire [3:0] stage5_58;
   wire [2:0] stage5_59;
   wire [1:0] stage5_60;
   wire [2:0] stage5_61;
   wire [2:0] stage5_62;
   wire [3:0] stage5_63;
   wire [5:0] stage5_64;
   wire [2:0] stage5_65;
   wire [1:0] stage5_66;
   wire [2:0] stage5_67;
   wire [1:0] stage5_68;
   wire [0:0] stage5_69;
   wire [0:0] stage5_70;
   wire [0:0] stage6_0;
   wire [1:0] stage6_1;
   wire [1:0] stage6_2;
   wire [1:0] stage6_3;
   wire [1:0] stage6_4;
   wire [1:0] stage6_5;
   wire [1:0] stage6_6;
   wire [1:0] stage6_7;
   wire [1:0] stage6_8;
   wire [1:0] stage6_9;
   wire [1:0] stage6_10;
   wire [1:0] stage6_11;
   wire [1:0] stage6_12;
   wire [1:0] stage6_13;
   wire [1:0] stage6_14;
   wire [1:0] stage6_15;
   wire [1:0] stage6_16;
   wire [1:0] stage6_17;
   wire [1:0] stage6_18;
   wire [1:0] stage6_19;
   wire [1:0] stage6_20;
   wire [1:0] stage6_21;
   wire [1:0] stage6_22;
   wire [1:0] stage6_23;
   wire [1:0] stage6_24;
   wire [1:0] stage6_25;
   wire [1:0] stage6_26;
   wire [1:0] stage6_27;
   wire [1:0] stage6_28;
   wire [1:0] stage6_29;
   wire [1:0] stage6_30;
   wire [1:0] stage6_31;
   wire [1:0] stage6_32;
   wire [1:0] stage6_33;
   wire [1:0] stage6_34;
   wire [1:0] stage6_35;
   wire [1:0] stage6_36;
   wire [1:0] stage6_37;
   wire [0:0] stage6_38;
   wire [1:0] stage6_39;
   wire [1:0] stage6_40;
   wire [1:0] stage6_41;
   wire [1:0] stage6_42;
   wire [1:0] stage6_43;
   wire [1:0] stage6_44;
   wire [1:0] stage6_45;
   wire [1:0] stage6_46;
   wire [1:0] stage6_47;
   wire [1:0] stage6_48;
   wire [1:0] stage6_49;
   wire [1:0] stage6_50;
   wire [1:0] stage6_51;
   wire [1:0] stage6_52;
   wire [1:0] stage6_53;
   wire [1:0] stage6_54;
   wire [1:0] stage6_55;
   wire [1:0] stage6_56;
   wire [1:0] stage6_57;
   wire [1:0] stage6_58;
   wire [1:0] stage6_59;
   wire [1:0] stage6_60;
   wire [1:0] stage6_61;
   wire [1:0] stage6_62;
   wire [0:0] stage6_63;
   wire [1:0] stage6_64;
   wire [1:0] stage6_65;
   wire [1:0] stage6_66;
   wire [1:0] stage6_67;
   wire [1:0] stage6_68;
   wire [0:0] stage6_69;
   wire [1:0] stage6_70;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage6_0;
   assign dst1 = stage6_1;
   assign dst2 = stage6_2;
   assign dst3 = stage6_3;
   assign dst4 = stage6_4;
   assign dst5 = stage6_5;
   assign dst6 = stage6_6;
   assign dst7 = stage6_7;
   assign dst8 = stage6_8;
   assign dst9 = stage6_9;
   assign dst10 = stage6_10;
   assign dst11 = stage6_11;
   assign dst12 = stage6_12;
   assign dst13 = stage6_13;
   assign dst14 = stage6_14;
   assign dst15 = stage6_15;
   assign dst16 = stage6_16;
   assign dst17 = stage6_17;
   assign dst18 = stage6_18;
   assign dst19 = stage6_19;
   assign dst20 = stage6_20;
   assign dst21 = stage6_21;
   assign dst22 = stage6_22;
   assign dst23 = stage6_23;
   assign dst24 = stage6_24;
   assign dst25 = stage6_25;
   assign dst26 = stage6_26;
   assign dst27 = stage6_27;
   assign dst28 = stage6_28;
   assign dst29 = stage6_29;
   assign dst30 = stage6_30;
   assign dst31 = stage6_31;
   assign dst32 = stage6_32;
   assign dst33 = stage6_33;
   assign dst34 = stage6_34;
   assign dst35 = stage6_35;
   assign dst36 = stage6_36;
   assign dst37 = stage6_37;
   assign dst38 = stage6_38;
   assign dst39 = stage6_39;
   assign dst40 = stage6_40;
   assign dst41 = stage6_41;
   assign dst42 = stage6_42;
   assign dst43 = stage6_43;
   assign dst44 = stage6_44;
   assign dst45 = stage6_45;
   assign dst46 = stage6_46;
   assign dst47 = stage6_47;
   assign dst48 = stage6_48;
   assign dst49 = stage6_49;
   assign dst50 = stage6_50;
   assign dst51 = stage6_51;
   assign dst52 = stage6_52;
   assign dst53 = stage6_53;
   assign dst54 = stage6_54;
   assign dst55 = stage6_55;
   assign dst56 = stage6_56;
   assign dst57 = stage6_57;
   assign dst58 = stage6_58;
   assign dst59 = stage6_59;
   assign dst60 = stage6_60;
   assign dst61 = stage6_61;
   assign dst62 = stage6_62;
   assign dst63 = stage6_63;
   assign dst64 = stage6_64;
   assign dst65 = stage6_65;
   assign dst66 = stage6_66;
   assign dst67 = stage6_67;
   assign dst68 = stage6_68;
   assign dst69 = stage6_69;
   assign dst70 = stage6_70;

   gpc117_4 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5], stage0_0[6]},
      {stage0_1[0]},
      {stage0_2[0]},
      {stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc117_4 gpc1 (
      {stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11], stage0_0[12], stage0_0[13]},
      {stage0_1[1]},
      {stage0_2[1]},
      {stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[14], stage0_0[15], stage0_0[16]},
      {stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7]},
      {stage0_2[2]},
      {stage0_3[0]},
      {stage1_4[0],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1163_5 gpc3 (
      {stage0_0[17], stage0_0[18], stage0_0[19]},
      {stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13]},
      {stage0_2[3]},
      {stage0_3[1]},
      {stage1_4[1],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc1163_5 gpc4 (
      {stage0_0[20], stage0_0[21], stage0_0[22]},
      {stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19]},
      {stage0_2[4]},
      {stage0_3[2]},
      {stage1_4[2],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc1163_5 gpc5 (
      {stage0_0[23], stage0_0[24], stage0_0[25]},
      {stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25]},
      {stage0_2[5]},
      {stage0_3[3]},
      {stage1_4[3],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc1163_5 gpc6 (
      {stage0_0[26], stage0_0[27], stage0_0[28]},
      {stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31]},
      {stage0_2[6]},
      {stage0_3[4]},
      {stage1_4[4],stage1_3[6],stage1_2[6],stage1_1[6],stage1_0[6]}
   );
   gpc1163_5 gpc7 (
      {stage0_0[29], stage0_0[30], stage0_0[31]},
      {stage0_1[32], stage0_1[33], stage0_1[34], stage0_1[35], stage0_1[36], stage0_1[37]},
      {stage0_2[7]},
      {stage0_3[5]},
      {stage1_4[5],stage1_3[7],stage1_2[7],stage1_1[7],stage1_0[7]}
   );
   gpc1163_5 gpc8 (
      {stage0_0[32], stage0_0[33], stage0_0[34]},
      {stage0_1[38], stage0_1[39], stage0_1[40], stage0_1[41], stage0_1[42], stage0_1[43]},
      {stage0_2[8]},
      {stage0_3[6]},
      {stage1_4[6],stage1_3[8],stage1_2[8],stage1_1[8],stage1_0[8]}
   );
   gpc1163_5 gpc9 (
      {stage0_0[35], stage0_0[36], stage0_0[37]},
      {stage0_1[44], stage0_1[45], stage0_1[46], stage0_1[47], stage0_1[48], stage0_1[49]},
      {stage0_2[9]},
      {stage0_3[7]},
      {stage1_4[7],stage1_3[9],stage1_2[9],stage1_1[9],stage1_0[9]}
   );
   gpc1163_5 gpc10 (
      {stage0_0[38], stage0_0[39], stage0_0[40]},
      {stage0_1[50], stage0_1[51], stage0_1[52], stage0_1[53], stage0_1[54], stage0_1[55]},
      {stage0_2[10]},
      {stage0_3[8]},
      {stage1_4[8],stage1_3[10],stage1_2[10],stage1_1[10],stage1_0[10]}
   );
   gpc1163_5 gpc11 (
      {stage0_0[41], stage0_0[42], stage0_0[43]},
      {stage0_1[56], stage0_1[57], stage0_1[58], stage0_1[59], stage0_1[60], stage0_1[61]},
      {stage0_2[11]},
      {stage0_3[9]},
      {stage1_4[9],stage1_3[11],stage1_2[11],stage1_1[11],stage1_0[11]}
   );
   gpc1163_5 gpc12 (
      {stage0_0[44], stage0_0[45], stage0_0[46]},
      {stage0_1[62], stage0_1[63], stage0_1[64], stage0_1[65], stage0_1[66], stage0_1[67]},
      {stage0_2[12]},
      {stage0_3[10]},
      {stage1_4[10],stage1_3[12],stage1_2[12],stage1_1[12],stage1_0[12]}
   );
   gpc1163_5 gpc13 (
      {stage0_0[47], stage0_0[48], stage0_0[49]},
      {stage0_1[68], stage0_1[69], stage0_1[70], stage0_1[71], stage0_1[72], stage0_1[73]},
      {stage0_2[13]},
      {stage0_3[11]},
      {stage1_4[11],stage1_3[13],stage1_2[13],stage1_1[13],stage1_0[13]}
   );
   gpc1163_5 gpc14 (
      {stage0_0[50], stage0_0[51], stage0_0[52]},
      {stage0_1[74], stage0_1[75], stage0_1[76], stage0_1[77], stage0_1[78], stage0_1[79]},
      {stage0_2[14]},
      {stage0_3[12]},
      {stage1_4[12],stage1_3[14],stage1_2[14],stage1_1[14],stage1_0[14]}
   );
   gpc1163_5 gpc15 (
      {stage0_0[53], stage0_0[54], stage0_0[55]},
      {stage0_1[80], stage0_1[81], stage0_1[82], stage0_1[83], stage0_1[84], stage0_1[85]},
      {stage0_2[15]},
      {stage0_3[13]},
      {stage1_4[13],stage1_3[15],stage1_2[15],stage1_1[15],stage1_0[15]}
   );
   gpc1163_5 gpc16 (
      {stage0_0[56], stage0_0[57], stage0_0[58]},
      {stage0_1[86], stage0_1[87], stage0_1[88], stage0_1[89], stage0_1[90], stage0_1[91]},
      {stage0_2[16]},
      {stage0_3[14]},
      {stage1_4[14],stage1_3[16],stage1_2[16],stage1_1[16],stage1_0[16]}
   );
   gpc1163_5 gpc17 (
      {stage0_0[59], stage0_0[60], stage0_0[61]},
      {stage0_1[92], stage0_1[93], stage0_1[94], stage0_1[95], stage0_1[96], stage0_1[97]},
      {stage0_2[17]},
      {stage0_3[15]},
      {stage1_4[15],stage1_3[17],stage1_2[17],stage1_1[17],stage1_0[17]}
   );
   gpc1163_5 gpc18 (
      {stage0_0[62], stage0_0[63], stage0_0[64]},
      {stage0_1[98], stage0_1[99], stage0_1[100], stage0_1[101], stage0_1[102], stage0_1[103]},
      {stage0_2[18]},
      {stage0_3[16]},
      {stage1_4[16],stage1_3[18],stage1_2[18],stage1_1[18],stage1_0[18]}
   );
   gpc1163_5 gpc19 (
      {stage0_0[65], stage0_0[66], stage0_0[67]},
      {stage0_1[104], stage0_1[105], stage0_1[106], stage0_1[107], stage0_1[108], stage0_1[109]},
      {stage0_2[19]},
      {stage0_3[17]},
      {stage1_4[17],stage1_3[19],stage1_2[19],stage1_1[19],stage1_0[19]}
   );
   gpc606_5 gpc20 (
      {stage0_0[68], stage0_0[69], stage0_0[70], stage0_0[71], stage0_0[72], stage0_0[73]},
      {stage0_2[20], stage0_2[21], stage0_2[22], stage0_2[23], stage0_2[24], stage0_2[25]},
      {stage1_4[18],stage1_3[20],stage1_2[20],stage1_1[20],stage1_0[20]}
   );
   gpc606_5 gpc21 (
      {stage0_0[74], stage0_0[75], stage0_0[76], stage0_0[77], stage0_0[78], stage0_0[79]},
      {stage0_2[26], stage0_2[27], stage0_2[28], stage0_2[29], stage0_2[30], stage0_2[31]},
      {stage1_4[19],stage1_3[21],stage1_2[21],stage1_1[21],stage1_0[21]}
   );
   gpc606_5 gpc22 (
      {stage0_0[80], stage0_0[81], stage0_0[82], stage0_0[83], stage0_0[84], stage0_0[85]},
      {stage0_2[32], stage0_2[33], stage0_2[34], stage0_2[35], stage0_2[36], stage0_2[37]},
      {stage1_4[20],stage1_3[22],stage1_2[22],stage1_1[22],stage1_0[22]}
   );
   gpc606_5 gpc23 (
      {stage0_0[86], stage0_0[87], stage0_0[88], stage0_0[89], stage0_0[90], stage0_0[91]},
      {stage0_2[38], stage0_2[39], stage0_2[40], stage0_2[41], stage0_2[42], stage0_2[43]},
      {stage1_4[21],stage1_3[23],stage1_2[23],stage1_1[23],stage1_0[23]}
   );
   gpc606_5 gpc24 (
      {stage0_0[92], stage0_0[93], stage0_0[94], stage0_0[95], stage0_0[96], stage0_0[97]},
      {stage0_2[44], stage0_2[45], stage0_2[46], stage0_2[47], stage0_2[48], stage0_2[49]},
      {stage1_4[22],stage1_3[24],stage1_2[24],stage1_1[24],stage1_0[24]}
   );
   gpc606_5 gpc25 (
      {stage0_0[98], stage0_0[99], stage0_0[100], stage0_0[101], stage0_0[102], stage0_0[103]},
      {stage0_2[50], stage0_2[51], stage0_2[52], stage0_2[53], stage0_2[54], stage0_2[55]},
      {stage1_4[23],stage1_3[25],stage1_2[25],stage1_1[25],stage1_0[25]}
   );
   gpc606_5 gpc26 (
      {stage0_0[104], stage0_0[105], stage0_0[106], stage0_0[107], stage0_0[108], stage0_0[109]},
      {stage0_2[56], stage0_2[57], stage0_2[58], stage0_2[59], stage0_2[60], stage0_2[61]},
      {stage1_4[24],stage1_3[26],stage1_2[26],stage1_1[26],stage1_0[26]}
   );
   gpc606_5 gpc27 (
      {stage0_0[110], stage0_0[111], stage0_0[112], stage0_0[113], stage0_0[114], stage0_0[115]},
      {stage0_2[62], stage0_2[63], stage0_2[64], stage0_2[65], stage0_2[66], stage0_2[67]},
      {stage1_4[25],stage1_3[27],stage1_2[27],stage1_1[27],stage1_0[27]}
   );
   gpc606_5 gpc28 (
      {stage0_0[116], stage0_0[117], stage0_0[118], stage0_0[119], stage0_0[120], stage0_0[121]},
      {stage0_2[68], stage0_2[69], stage0_2[70], stage0_2[71], stage0_2[72], stage0_2[73]},
      {stage1_4[26],stage1_3[28],stage1_2[28],stage1_1[28],stage1_0[28]}
   );
   gpc606_5 gpc29 (
      {stage0_0[122], stage0_0[123], stage0_0[124], stage0_0[125], stage0_0[126], stage0_0[127]},
      {stage0_2[74], stage0_2[75], stage0_2[76], stage0_2[77], stage0_2[78], stage0_2[79]},
      {stage1_4[27],stage1_3[29],stage1_2[29],stage1_1[29],stage1_0[29]}
   );
   gpc606_5 gpc30 (
      {stage0_1[110], stage0_1[111], stage0_1[112], stage0_1[113], stage0_1[114], stage0_1[115]},
      {stage0_3[18], stage0_3[19], stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23]},
      {stage1_5[0],stage1_4[28],stage1_3[30],stage1_2[30],stage1_1[30]}
   );
   gpc606_5 gpc31 (
      {stage0_1[116], stage0_1[117], stage0_1[118], stage0_1[119], stage0_1[120], stage0_1[121]},
      {stage0_3[24], stage0_3[25], stage0_3[26], stage0_3[27], stage0_3[28], stage0_3[29]},
      {stage1_5[1],stage1_4[29],stage1_3[31],stage1_2[31],stage1_1[31]}
   );
   gpc606_5 gpc32 (
      {stage0_1[122], stage0_1[123], stage0_1[124], stage0_1[125], stage0_1[126], stage0_1[127]},
      {stage0_3[30], stage0_3[31], stage0_3[32], stage0_3[33], stage0_3[34], stage0_3[35]},
      {stage1_5[2],stage1_4[30],stage1_3[32],stage1_2[32],stage1_1[32]}
   );
   gpc606_5 gpc33 (
      {stage0_2[80], stage0_2[81], stage0_2[82], stage0_2[83], stage0_2[84], stage0_2[85]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[3],stage1_4[31],stage1_3[33],stage1_2[33]}
   );
   gpc606_5 gpc34 (
      {stage0_2[86], stage0_2[87], stage0_2[88], stage0_2[89], stage0_2[90], stage0_2[91]},
      {stage0_4[6], stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11]},
      {stage1_6[1],stage1_5[4],stage1_4[32],stage1_3[34],stage1_2[34]}
   );
   gpc606_5 gpc35 (
      {stage0_2[92], stage0_2[93], stage0_2[94], stage0_2[95], stage0_2[96], stage0_2[97]},
      {stage0_4[12], stage0_4[13], stage0_4[14], stage0_4[15], stage0_4[16], stage0_4[17]},
      {stage1_6[2],stage1_5[5],stage1_4[33],stage1_3[35],stage1_2[35]}
   );
   gpc606_5 gpc36 (
      {stage0_2[98], stage0_2[99], stage0_2[100], stage0_2[101], stage0_2[102], stage0_2[103]},
      {stage0_4[18], stage0_4[19], stage0_4[20], stage0_4[21], stage0_4[22], stage0_4[23]},
      {stage1_6[3],stage1_5[6],stage1_4[34],stage1_3[36],stage1_2[36]}
   );
   gpc606_5 gpc37 (
      {stage0_2[104], stage0_2[105], stage0_2[106], stage0_2[107], stage0_2[108], stage0_2[109]},
      {stage0_4[24], stage0_4[25], stage0_4[26], stage0_4[27], stage0_4[28], stage0_4[29]},
      {stage1_6[4],stage1_5[7],stage1_4[35],stage1_3[37],stage1_2[37]}
   );
   gpc606_5 gpc38 (
      {stage0_2[110], stage0_2[111], stage0_2[112], stage0_2[113], stage0_2[114], stage0_2[115]},
      {stage0_4[30], stage0_4[31], stage0_4[32], stage0_4[33], stage0_4[34], stage0_4[35]},
      {stage1_6[5],stage1_5[8],stage1_4[36],stage1_3[38],stage1_2[38]}
   );
   gpc615_5 gpc39 (
      {stage0_2[116], stage0_2[117], stage0_2[118], stage0_2[119], stage0_2[120]},
      {stage0_3[36]},
      {stage0_4[36], stage0_4[37], stage0_4[38], stage0_4[39], stage0_4[40], stage0_4[41]},
      {stage1_6[6],stage1_5[9],stage1_4[37],stage1_3[39],stage1_2[39]}
   );
   gpc615_5 gpc40 (
      {stage0_3[37], stage0_3[38], stage0_3[39], stage0_3[40], stage0_3[41]},
      {stage0_4[42]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[7],stage1_5[10],stage1_4[38],stage1_3[40]}
   );
   gpc615_5 gpc41 (
      {stage0_3[42], stage0_3[43], stage0_3[44], stage0_3[45], stage0_3[46]},
      {stage0_4[43]},
      {stage0_5[6], stage0_5[7], stage0_5[8], stage0_5[9], stage0_5[10], stage0_5[11]},
      {stage1_7[1],stage1_6[8],stage1_5[11],stage1_4[39],stage1_3[41]}
   );
   gpc615_5 gpc42 (
      {stage0_3[47], stage0_3[48], stage0_3[49], stage0_3[50], stage0_3[51]},
      {stage0_4[44]},
      {stage0_5[12], stage0_5[13], stage0_5[14], stage0_5[15], stage0_5[16], stage0_5[17]},
      {stage1_7[2],stage1_6[9],stage1_5[12],stage1_4[40],stage1_3[42]}
   );
   gpc615_5 gpc43 (
      {stage0_3[52], stage0_3[53], stage0_3[54], stage0_3[55], stage0_3[56]},
      {stage0_4[45]},
      {stage0_5[18], stage0_5[19], stage0_5[20], stage0_5[21], stage0_5[22], stage0_5[23]},
      {stage1_7[3],stage1_6[10],stage1_5[13],stage1_4[41],stage1_3[43]}
   );
   gpc615_5 gpc44 (
      {stage0_3[57], stage0_3[58], stage0_3[59], stage0_3[60], stage0_3[61]},
      {stage0_4[46]},
      {stage0_5[24], stage0_5[25], stage0_5[26], stage0_5[27], stage0_5[28], stage0_5[29]},
      {stage1_7[4],stage1_6[11],stage1_5[14],stage1_4[42],stage1_3[44]}
   );
   gpc615_5 gpc45 (
      {stage0_3[62], stage0_3[63], stage0_3[64], stage0_3[65], stage0_3[66]},
      {stage0_4[47]},
      {stage0_5[30], stage0_5[31], stage0_5[32], stage0_5[33], stage0_5[34], stage0_5[35]},
      {stage1_7[5],stage1_6[12],stage1_5[15],stage1_4[43],stage1_3[45]}
   );
   gpc615_5 gpc46 (
      {stage0_3[67], stage0_3[68], stage0_3[69], stage0_3[70], stage0_3[71]},
      {stage0_4[48]},
      {stage0_5[36], stage0_5[37], stage0_5[38], stage0_5[39], stage0_5[40], stage0_5[41]},
      {stage1_7[6],stage1_6[13],stage1_5[16],stage1_4[44],stage1_3[46]}
   );
   gpc615_5 gpc47 (
      {stage0_3[72], stage0_3[73], stage0_3[74], stage0_3[75], stage0_3[76]},
      {stage0_4[49]},
      {stage0_5[42], stage0_5[43], stage0_5[44], stage0_5[45], stage0_5[46], stage0_5[47]},
      {stage1_7[7],stage1_6[14],stage1_5[17],stage1_4[45],stage1_3[47]}
   );
   gpc615_5 gpc48 (
      {stage0_3[77], stage0_3[78], stage0_3[79], stage0_3[80], stage0_3[81]},
      {stage0_4[50]},
      {stage0_5[48], stage0_5[49], stage0_5[50], stage0_5[51], stage0_5[52], stage0_5[53]},
      {stage1_7[8],stage1_6[15],stage1_5[18],stage1_4[46],stage1_3[48]}
   );
   gpc615_5 gpc49 (
      {stage0_3[82], stage0_3[83], stage0_3[84], stage0_3[85], stage0_3[86]},
      {stage0_4[51]},
      {stage0_5[54], stage0_5[55], stage0_5[56], stage0_5[57], stage0_5[58], stage0_5[59]},
      {stage1_7[9],stage1_6[16],stage1_5[19],stage1_4[47],stage1_3[49]}
   );
   gpc615_5 gpc50 (
      {stage0_3[87], stage0_3[88], stage0_3[89], stage0_3[90], stage0_3[91]},
      {stage0_4[52]},
      {stage0_5[60], stage0_5[61], stage0_5[62], stage0_5[63], stage0_5[64], stage0_5[65]},
      {stage1_7[10],stage1_6[17],stage1_5[20],stage1_4[48],stage1_3[50]}
   );
   gpc615_5 gpc51 (
      {stage0_3[92], stage0_3[93], stage0_3[94], stage0_3[95], stage0_3[96]},
      {stage0_4[53]},
      {stage0_5[66], stage0_5[67], stage0_5[68], stage0_5[69], stage0_5[70], stage0_5[71]},
      {stage1_7[11],stage1_6[18],stage1_5[21],stage1_4[49],stage1_3[51]}
   );
   gpc615_5 gpc52 (
      {stage0_3[97], stage0_3[98], stage0_3[99], stage0_3[100], stage0_3[101]},
      {stage0_4[54]},
      {stage0_5[72], stage0_5[73], stage0_5[74], stage0_5[75], stage0_5[76], stage0_5[77]},
      {stage1_7[12],stage1_6[19],stage1_5[22],stage1_4[50],stage1_3[52]}
   );
   gpc615_5 gpc53 (
      {stage0_3[102], stage0_3[103], stage0_3[104], stage0_3[105], stage0_3[106]},
      {stage0_4[55]},
      {stage0_5[78], stage0_5[79], stage0_5[80], stage0_5[81], stage0_5[82], stage0_5[83]},
      {stage1_7[13],stage1_6[20],stage1_5[23],stage1_4[51],stage1_3[53]}
   );
   gpc615_5 gpc54 (
      {stage0_3[107], stage0_3[108], stage0_3[109], stage0_3[110], stage0_3[111]},
      {stage0_4[56]},
      {stage0_5[84], stage0_5[85], stage0_5[86], stage0_5[87], stage0_5[88], stage0_5[89]},
      {stage1_7[14],stage1_6[21],stage1_5[24],stage1_4[52],stage1_3[54]}
   );
   gpc615_5 gpc55 (
      {stage0_3[112], stage0_3[113], stage0_3[114], stage0_3[115], stage0_3[116]},
      {stage0_4[57]},
      {stage0_5[90], stage0_5[91], stage0_5[92], stage0_5[93], stage0_5[94], stage0_5[95]},
      {stage1_7[15],stage1_6[22],stage1_5[25],stage1_4[53],stage1_3[55]}
   );
   gpc606_5 gpc56 (
      {stage0_4[58], stage0_4[59], stage0_4[60], stage0_4[61], stage0_4[62], stage0_4[63]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[16],stage1_6[23],stage1_5[26],stage1_4[54]}
   );
   gpc606_5 gpc57 (
      {stage0_4[64], stage0_4[65], stage0_4[66], stage0_4[67], stage0_4[68], stage0_4[69]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9], stage0_6[10], stage0_6[11]},
      {stage1_8[1],stage1_7[17],stage1_6[24],stage1_5[27],stage1_4[55]}
   );
   gpc606_5 gpc58 (
      {stage0_4[70], stage0_4[71], stage0_4[72], stage0_4[73], stage0_4[74], stage0_4[75]},
      {stage0_6[12], stage0_6[13], stage0_6[14], stage0_6[15], stage0_6[16], stage0_6[17]},
      {stage1_8[2],stage1_7[18],stage1_6[25],stage1_5[28],stage1_4[56]}
   );
   gpc606_5 gpc59 (
      {stage0_4[76], stage0_4[77], stage0_4[78], stage0_4[79], stage0_4[80], stage0_4[81]},
      {stage0_6[18], stage0_6[19], stage0_6[20], stage0_6[21], stage0_6[22], stage0_6[23]},
      {stage1_8[3],stage1_7[19],stage1_6[26],stage1_5[29],stage1_4[57]}
   );
   gpc606_5 gpc60 (
      {stage0_4[82], stage0_4[83], stage0_4[84], stage0_4[85], stage0_4[86], stage0_4[87]},
      {stage0_6[24], stage0_6[25], stage0_6[26], stage0_6[27], stage0_6[28], stage0_6[29]},
      {stage1_8[4],stage1_7[20],stage1_6[27],stage1_5[30],stage1_4[58]}
   );
   gpc606_5 gpc61 (
      {stage0_4[88], stage0_4[89], stage0_4[90], stage0_4[91], stage0_4[92], stage0_4[93]},
      {stage0_6[30], stage0_6[31], stage0_6[32], stage0_6[33], stage0_6[34], stage0_6[35]},
      {stage1_8[5],stage1_7[21],stage1_6[28],stage1_5[31],stage1_4[59]}
   );
   gpc606_5 gpc62 (
      {stage0_4[94], stage0_4[95], stage0_4[96], stage0_4[97], stage0_4[98], stage0_4[99]},
      {stage0_6[36], stage0_6[37], stage0_6[38], stage0_6[39], stage0_6[40], stage0_6[41]},
      {stage1_8[6],stage1_7[22],stage1_6[29],stage1_5[32],stage1_4[60]}
   );
   gpc606_5 gpc63 (
      {stage0_4[100], stage0_4[101], stage0_4[102], stage0_4[103], stage0_4[104], stage0_4[105]},
      {stage0_6[42], stage0_6[43], stage0_6[44], stage0_6[45], stage0_6[46], stage0_6[47]},
      {stage1_8[7],stage1_7[23],stage1_6[30],stage1_5[33],stage1_4[61]}
   );
   gpc606_5 gpc64 (
      {stage0_4[106], stage0_4[107], stage0_4[108], stage0_4[109], stage0_4[110], stage0_4[111]},
      {stage0_6[48], stage0_6[49], stage0_6[50], stage0_6[51], stage0_6[52], stage0_6[53]},
      {stage1_8[8],stage1_7[24],stage1_6[31],stage1_5[34],stage1_4[62]}
   );
   gpc606_5 gpc65 (
      {stage0_4[112], stage0_4[113], stage0_4[114], stage0_4[115], stage0_4[116], stage0_4[117]},
      {stage0_6[54], stage0_6[55], stage0_6[56], stage0_6[57], stage0_6[58], stage0_6[59]},
      {stage1_8[9],stage1_7[25],stage1_6[32],stage1_5[35],stage1_4[63]}
   );
   gpc615_5 gpc66 (
      {stage0_4[118], stage0_4[119], stage0_4[120], stage0_4[121], stage0_4[122]},
      {stage0_5[96]},
      {stage0_6[60], stage0_6[61], stage0_6[62], stage0_6[63], stage0_6[64], stage0_6[65]},
      {stage1_8[10],stage1_7[26],stage1_6[33],stage1_5[36],stage1_4[64]}
   );
   gpc615_5 gpc67 (
      {stage0_4[123], stage0_4[124], stage0_4[125], stage0_4[126], stage0_4[127]},
      {stage0_5[97]},
      {stage0_6[66], stage0_6[67], stage0_6[68], stage0_6[69], stage0_6[70], stage0_6[71]},
      {stage1_8[11],stage1_7[27],stage1_6[34],stage1_5[37],stage1_4[65]}
   );
   gpc615_5 gpc68 (
      {stage0_5[98], stage0_5[99], stage0_5[100], stage0_5[101], stage0_5[102]},
      {stage0_6[72]},
      {stage0_7[0], stage0_7[1], stage0_7[2], stage0_7[3], stage0_7[4], stage0_7[5]},
      {stage1_9[0],stage1_8[12],stage1_7[28],stage1_6[35],stage1_5[38]}
   );
   gpc615_5 gpc69 (
      {stage0_5[103], stage0_5[104], stage0_5[105], stage0_5[106], stage0_5[107]},
      {stage0_6[73]},
      {stage0_7[6], stage0_7[7], stage0_7[8], stage0_7[9], stage0_7[10], stage0_7[11]},
      {stage1_9[1],stage1_8[13],stage1_7[29],stage1_6[36],stage1_5[39]}
   );
   gpc615_5 gpc70 (
      {stage0_5[108], stage0_5[109], stage0_5[110], stage0_5[111], stage0_5[112]},
      {stage0_6[74]},
      {stage0_7[12], stage0_7[13], stage0_7[14], stage0_7[15], stage0_7[16], stage0_7[17]},
      {stage1_9[2],stage1_8[14],stage1_7[30],stage1_6[37],stage1_5[40]}
   );
   gpc615_5 gpc71 (
      {stage0_5[113], stage0_5[114], stage0_5[115], stage0_5[116], stage0_5[117]},
      {stage0_6[75]},
      {stage0_7[18], stage0_7[19], stage0_7[20], stage0_7[21], stage0_7[22], stage0_7[23]},
      {stage1_9[3],stage1_8[15],stage1_7[31],stage1_6[38],stage1_5[41]}
   );
   gpc623_5 gpc72 (
      {stage0_6[76], stage0_6[77], stage0_6[78]},
      {stage0_7[24], stage0_7[25]},
      {stage0_8[0], stage0_8[1], stage0_8[2], stage0_8[3], stage0_8[4], stage0_8[5]},
      {stage1_10[0],stage1_9[4],stage1_8[16],stage1_7[32],stage1_6[39]}
   );
   gpc606_5 gpc73 (
      {stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29], stage0_7[30], stage0_7[31]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[1],stage1_9[5],stage1_8[17],stage1_7[33]}
   );
   gpc606_5 gpc74 (
      {stage0_7[32], stage0_7[33], stage0_7[34], stage0_7[35], stage0_7[36], stage0_7[37]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[2],stage1_9[6],stage1_8[18],stage1_7[34]}
   );
   gpc606_5 gpc75 (
      {stage0_7[38], stage0_7[39], stage0_7[40], stage0_7[41], stage0_7[42], stage0_7[43]},
      {stage0_9[12], stage0_9[13], stage0_9[14], stage0_9[15], stage0_9[16], stage0_9[17]},
      {stage1_11[2],stage1_10[3],stage1_9[7],stage1_8[19],stage1_7[35]}
   );
   gpc606_5 gpc76 (
      {stage0_7[44], stage0_7[45], stage0_7[46], stage0_7[47], stage0_7[48], stage0_7[49]},
      {stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22], stage0_9[23]},
      {stage1_11[3],stage1_10[4],stage1_9[8],stage1_8[20],stage1_7[36]}
   );
   gpc606_5 gpc77 (
      {stage0_7[50], stage0_7[51], stage0_7[52], stage0_7[53], stage0_7[54], stage0_7[55]},
      {stage0_9[24], stage0_9[25], stage0_9[26], stage0_9[27], stage0_9[28], stage0_9[29]},
      {stage1_11[4],stage1_10[5],stage1_9[9],stage1_8[21],stage1_7[37]}
   );
   gpc606_5 gpc78 (
      {stage0_7[56], stage0_7[57], stage0_7[58], stage0_7[59], stage0_7[60], stage0_7[61]},
      {stage0_9[30], stage0_9[31], stage0_9[32], stage0_9[33], stage0_9[34], stage0_9[35]},
      {stage1_11[5],stage1_10[6],stage1_9[10],stage1_8[22],stage1_7[38]}
   );
   gpc606_5 gpc79 (
      {stage0_7[62], stage0_7[63], stage0_7[64], stage0_7[65], stage0_7[66], stage0_7[67]},
      {stage0_9[36], stage0_9[37], stage0_9[38], stage0_9[39], stage0_9[40], stage0_9[41]},
      {stage1_11[6],stage1_10[7],stage1_9[11],stage1_8[23],stage1_7[39]}
   );
   gpc606_5 gpc80 (
      {stage0_7[68], stage0_7[69], stage0_7[70], stage0_7[71], stage0_7[72], stage0_7[73]},
      {stage0_9[42], stage0_9[43], stage0_9[44], stage0_9[45], stage0_9[46], stage0_9[47]},
      {stage1_11[7],stage1_10[8],stage1_9[12],stage1_8[24],stage1_7[40]}
   );
   gpc606_5 gpc81 (
      {stage0_7[74], stage0_7[75], stage0_7[76], stage0_7[77], stage0_7[78], stage0_7[79]},
      {stage0_9[48], stage0_9[49], stage0_9[50], stage0_9[51], stage0_9[52], stage0_9[53]},
      {stage1_11[8],stage1_10[9],stage1_9[13],stage1_8[25],stage1_7[41]}
   );
   gpc606_5 gpc82 (
      {stage0_7[80], stage0_7[81], stage0_7[82], stage0_7[83], stage0_7[84], stage0_7[85]},
      {stage0_9[54], stage0_9[55], stage0_9[56], stage0_9[57], stage0_9[58], stage0_9[59]},
      {stage1_11[9],stage1_10[10],stage1_9[14],stage1_8[26],stage1_7[42]}
   );
   gpc606_5 gpc83 (
      {stage0_7[86], stage0_7[87], stage0_7[88], stage0_7[89], stage0_7[90], stage0_7[91]},
      {stage0_9[60], stage0_9[61], stage0_9[62], stage0_9[63], stage0_9[64], stage0_9[65]},
      {stage1_11[10],stage1_10[11],stage1_9[15],stage1_8[27],stage1_7[43]}
   );
   gpc606_5 gpc84 (
      {stage0_7[92], stage0_7[93], stage0_7[94], stage0_7[95], stage0_7[96], stage0_7[97]},
      {stage0_9[66], stage0_9[67], stage0_9[68], stage0_9[69], stage0_9[70], stage0_9[71]},
      {stage1_11[11],stage1_10[12],stage1_9[16],stage1_8[28],stage1_7[44]}
   );
   gpc615_5 gpc85 (
      {stage0_7[98], stage0_7[99], stage0_7[100], stage0_7[101], stage0_7[102]},
      {stage0_8[6]},
      {stage0_9[72], stage0_9[73], stage0_9[74], stage0_9[75], stage0_9[76], stage0_9[77]},
      {stage1_11[12],stage1_10[13],stage1_9[17],stage1_8[29],stage1_7[45]}
   );
   gpc606_5 gpc86 (
      {stage0_8[7], stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11], stage0_8[12]},
      {stage0_10[0], stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5]},
      {stage1_12[0],stage1_11[13],stage1_10[14],stage1_9[18],stage1_8[30]}
   );
   gpc606_5 gpc87 (
      {stage0_8[13], stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17], stage0_8[18]},
      {stage0_10[6], stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11]},
      {stage1_12[1],stage1_11[14],stage1_10[15],stage1_9[19],stage1_8[31]}
   );
   gpc606_5 gpc88 (
      {stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23], stage0_8[24]},
      {stage0_10[12], stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17]},
      {stage1_12[2],stage1_11[15],stage1_10[16],stage1_9[20],stage1_8[32]}
   );
   gpc606_5 gpc89 (
      {stage0_8[25], stage0_8[26], stage0_8[27], stage0_8[28], stage0_8[29], stage0_8[30]},
      {stage0_10[18], stage0_10[19], stage0_10[20], stage0_10[21], stage0_10[22], stage0_10[23]},
      {stage1_12[3],stage1_11[16],stage1_10[17],stage1_9[21],stage1_8[33]}
   );
   gpc606_5 gpc90 (
      {stage0_8[31], stage0_8[32], stage0_8[33], stage0_8[34], stage0_8[35], stage0_8[36]},
      {stage0_10[24], stage0_10[25], stage0_10[26], stage0_10[27], stage0_10[28], stage0_10[29]},
      {stage1_12[4],stage1_11[17],stage1_10[18],stage1_9[22],stage1_8[34]}
   );
   gpc606_5 gpc91 (
      {stage0_8[37], stage0_8[38], stage0_8[39], stage0_8[40], stage0_8[41], stage0_8[42]},
      {stage0_10[30], stage0_10[31], stage0_10[32], stage0_10[33], stage0_10[34], stage0_10[35]},
      {stage1_12[5],stage1_11[18],stage1_10[19],stage1_9[23],stage1_8[35]}
   );
   gpc606_5 gpc92 (
      {stage0_8[43], stage0_8[44], stage0_8[45], stage0_8[46], stage0_8[47], stage0_8[48]},
      {stage0_10[36], stage0_10[37], stage0_10[38], stage0_10[39], stage0_10[40], stage0_10[41]},
      {stage1_12[6],stage1_11[19],stage1_10[20],stage1_9[24],stage1_8[36]}
   );
   gpc606_5 gpc93 (
      {stage0_8[49], stage0_8[50], stage0_8[51], stage0_8[52], stage0_8[53], stage0_8[54]},
      {stage0_10[42], stage0_10[43], stage0_10[44], stage0_10[45], stage0_10[46], stage0_10[47]},
      {stage1_12[7],stage1_11[20],stage1_10[21],stage1_9[25],stage1_8[37]}
   );
   gpc606_5 gpc94 (
      {stage0_8[55], stage0_8[56], stage0_8[57], stage0_8[58], stage0_8[59], stage0_8[60]},
      {stage0_10[48], stage0_10[49], stage0_10[50], stage0_10[51], stage0_10[52], stage0_10[53]},
      {stage1_12[8],stage1_11[21],stage1_10[22],stage1_9[26],stage1_8[38]}
   );
   gpc606_5 gpc95 (
      {stage0_8[61], stage0_8[62], stage0_8[63], stage0_8[64], stage0_8[65], stage0_8[66]},
      {stage0_10[54], stage0_10[55], stage0_10[56], stage0_10[57], stage0_10[58], stage0_10[59]},
      {stage1_12[9],stage1_11[22],stage1_10[23],stage1_9[27],stage1_8[39]}
   );
   gpc606_5 gpc96 (
      {stage0_8[67], stage0_8[68], stage0_8[69], stage0_8[70], stage0_8[71], stage0_8[72]},
      {stage0_10[60], stage0_10[61], stage0_10[62], stage0_10[63], stage0_10[64], stage0_10[65]},
      {stage1_12[10],stage1_11[23],stage1_10[24],stage1_9[28],stage1_8[40]}
   );
   gpc606_5 gpc97 (
      {stage0_8[73], stage0_8[74], stage0_8[75], stage0_8[76], stage0_8[77], stage0_8[78]},
      {stage0_10[66], stage0_10[67], stage0_10[68], stage0_10[69], stage0_10[70], stage0_10[71]},
      {stage1_12[11],stage1_11[24],stage1_10[25],stage1_9[29],stage1_8[41]}
   );
   gpc606_5 gpc98 (
      {stage0_8[79], stage0_8[80], stage0_8[81], stage0_8[82], stage0_8[83], stage0_8[84]},
      {stage0_10[72], stage0_10[73], stage0_10[74], stage0_10[75], stage0_10[76], stage0_10[77]},
      {stage1_12[12],stage1_11[25],stage1_10[26],stage1_9[30],stage1_8[42]}
   );
   gpc606_5 gpc99 (
      {stage0_8[85], stage0_8[86], stage0_8[87], stage0_8[88], stage0_8[89], stage0_8[90]},
      {stage0_10[78], stage0_10[79], stage0_10[80], stage0_10[81], stage0_10[82], stage0_10[83]},
      {stage1_12[13],stage1_11[26],stage1_10[27],stage1_9[31],stage1_8[43]}
   );
   gpc606_5 gpc100 (
      {stage0_8[91], stage0_8[92], stage0_8[93], stage0_8[94], stage0_8[95], stage0_8[96]},
      {stage0_10[84], stage0_10[85], stage0_10[86], stage0_10[87], stage0_10[88], stage0_10[89]},
      {stage1_12[14],stage1_11[27],stage1_10[28],stage1_9[32],stage1_8[44]}
   );
   gpc606_5 gpc101 (
      {stage0_8[97], stage0_8[98], stage0_8[99], stage0_8[100], stage0_8[101], stage0_8[102]},
      {stage0_10[90], stage0_10[91], stage0_10[92], stage0_10[93], stage0_10[94], stage0_10[95]},
      {stage1_12[15],stage1_11[28],stage1_10[29],stage1_9[33],stage1_8[45]}
   );
   gpc606_5 gpc102 (
      {stage0_8[103], stage0_8[104], stage0_8[105], stage0_8[106], stage0_8[107], stage0_8[108]},
      {stage0_10[96], stage0_10[97], stage0_10[98], stage0_10[99], stage0_10[100], stage0_10[101]},
      {stage1_12[16],stage1_11[29],stage1_10[30],stage1_9[34],stage1_8[46]}
   );
   gpc615_5 gpc103 (
      {stage0_9[78], stage0_9[79], stage0_9[80], stage0_9[81], stage0_9[82]},
      {stage0_10[102]},
      {stage0_11[0], stage0_11[1], stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5]},
      {stage1_13[0],stage1_12[17],stage1_11[30],stage1_10[31],stage1_9[35]}
   );
   gpc615_5 gpc104 (
      {stage0_9[83], stage0_9[84], stage0_9[85], stage0_9[86], stage0_9[87]},
      {stage0_10[103]},
      {stage0_11[6], stage0_11[7], stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11]},
      {stage1_13[1],stage1_12[18],stage1_11[31],stage1_10[32],stage1_9[36]}
   );
   gpc615_5 gpc105 (
      {stage0_9[88], stage0_9[89], stage0_9[90], stage0_9[91], stage0_9[92]},
      {stage0_10[104]},
      {stage0_11[12], stage0_11[13], stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17]},
      {stage1_13[2],stage1_12[19],stage1_11[32],stage1_10[33],stage1_9[37]}
   );
   gpc615_5 gpc106 (
      {stage0_9[93], stage0_9[94], stage0_9[95], stage0_9[96], stage0_9[97]},
      {stage0_10[105]},
      {stage0_11[18], stage0_11[19], stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23]},
      {stage1_13[3],stage1_12[20],stage1_11[33],stage1_10[34],stage1_9[38]}
   );
   gpc615_5 gpc107 (
      {stage0_9[98], stage0_9[99], stage0_9[100], stage0_9[101], stage0_9[102]},
      {stage0_10[106]},
      {stage0_11[24], stage0_11[25], stage0_11[26], stage0_11[27], stage0_11[28], stage0_11[29]},
      {stage1_13[4],stage1_12[21],stage1_11[34],stage1_10[35],stage1_9[39]}
   );
   gpc615_5 gpc108 (
      {stage0_9[103], stage0_9[104], stage0_9[105], stage0_9[106], stage0_9[107]},
      {stage0_10[107]},
      {stage0_11[30], stage0_11[31], stage0_11[32], stage0_11[33], stage0_11[34], stage0_11[35]},
      {stage1_13[5],stage1_12[22],stage1_11[35],stage1_10[36],stage1_9[40]}
   );
   gpc615_5 gpc109 (
      {stage0_10[108], stage0_10[109], stage0_10[110], stage0_10[111], stage0_10[112]},
      {stage0_11[36]},
      {stage0_12[0], stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5]},
      {stage1_14[0],stage1_13[6],stage1_12[23],stage1_11[36],stage1_10[37]}
   );
   gpc615_5 gpc110 (
      {stage0_10[113], stage0_10[114], stage0_10[115], stage0_10[116], stage0_10[117]},
      {stage0_11[37]},
      {stage0_12[6], stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11]},
      {stage1_14[1],stage1_13[7],stage1_12[24],stage1_11[37],stage1_10[38]}
   );
   gpc615_5 gpc111 (
      {stage0_10[118], stage0_10[119], stage0_10[120], stage0_10[121], stage0_10[122]},
      {stage0_11[38]},
      {stage0_12[12], stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17]},
      {stage1_14[2],stage1_13[8],stage1_12[25],stage1_11[38],stage1_10[39]}
   );
   gpc615_5 gpc112 (
      {stage0_10[123], stage0_10[124], stage0_10[125], stage0_10[126], stage0_10[127]},
      {stage0_11[39]},
      {stage0_12[18], stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23]},
      {stage1_14[3],stage1_13[9],stage1_12[26],stage1_11[39],stage1_10[40]}
   );
   gpc117_4 gpc113 (
      {stage0_11[40], stage0_11[41], stage0_11[42], stage0_11[43], stage0_11[44], stage0_11[45], stage0_11[46]},
      {stage0_12[24]},
      {stage0_13[0]},
      {stage1_14[4],stage1_13[10],stage1_12[27],stage1_11[40]}
   );
   gpc117_4 gpc114 (
      {stage0_11[47], stage0_11[48], stage0_11[49], stage0_11[50], stage0_11[51], stage0_11[52], stage0_11[53]},
      {stage0_12[25]},
      {stage0_13[1]},
      {stage1_14[5],stage1_13[11],stage1_12[28],stage1_11[41]}
   );
   gpc117_4 gpc115 (
      {stage0_11[54], stage0_11[55], stage0_11[56], stage0_11[57], stage0_11[58], stage0_11[59], stage0_11[60]},
      {stage0_12[26]},
      {stage0_13[2]},
      {stage1_14[6],stage1_13[12],stage1_12[29],stage1_11[42]}
   );
   gpc117_4 gpc116 (
      {stage0_11[61], stage0_11[62], stage0_11[63], stage0_11[64], stage0_11[65], stage0_11[66], stage0_11[67]},
      {stage0_12[27]},
      {stage0_13[3]},
      {stage1_14[7],stage1_13[13],stage1_12[30],stage1_11[43]}
   );
   gpc615_5 gpc117 (
      {stage0_11[68], stage0_11[69], stage0_11[70], stage0_11[71], stage0_11[72]},
      {stage0_12[28]},
      {stage0_13[4], stage0_13[5], stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9]},
      {stage1_15[0],stage1_14[8],stage1_13[14],stage1_12[31],stage1_11[44]}
   );
   gpc615_5 gpc118 (
      {stage0_11[73], stage0_11[74], stage0_11[75], stage0_11[76], stage0_11[77]},
      {stage0_12[29]},
      {stage0_13[10], stage0_13[11], stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15]},
      {stage1_15[1],stage1_14[9],stage1_13[15],stage1_12[32],stage1_11[45]}
   );
   gpc615_5 gpc119 (
      {stage0_11[78], stage0_11[79], stage0_11[80], stage0_11[81], stage0_11[82]},
      {stage0_12[30]},
      {stage0_13[16], stage0_13[17], stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21]},
      {stage1_15[2],stage1_14[10],stage1_13[16],stage1_12[33],stage1_11[46]}
   );
   gpc615_5 gpc120 (
      {stage0_11[83], stage0_11[84], stage0_11[85], stage0_11[86], stage0_11[87]},
      {stage0_12[31]},
      {stage0_13[22], stage0_13[23], stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27]},
      {stage1_15[3],stage1_14[11],stage1_13[17],stage1_12[34],stage1_11[47]}
   );
   gpc615_5 gpc121 (
      {stage0_11[88], stage0_11[89], stage0_11[90], stage0_11[91], stage0_11[92]},
      {stage0_12[32]},
      {stage0_13[28], stage0_13[29], stage0_13[30], stage0_13[31], stage0_13[32], stage0_13[33]},
      {stage1_15[4],stage1_14[12],stage1_13[18],stage1_12[35],stage1_11[48]}
   );
   gpc615_5 gpc122 (
      {stage0_11[93], stage0_11[94], stage0_11[95], stage0_11[96], stage0_11[97]},
      {stage0_12[33]},
      {stage0_13[34], stage0_13[35], stage0_13[36], stage0_13[37], stage0_13[38], stage0_13[39]},
      {stage1_15[5],stage1_14[13],stage1_13[19],stage1_12[36],stage1_11[49]}
   );
   gpc615_5 gpc123 (
      {stage0_11[98], stage0_11[99], stage0_11[100], stage0_11[101], stage0_11[102]},
      {stage0_12[34]},
      {stage0_13[40], stage0_13[41], stage0_13[42], stage0_13[43], stage0_13[44], stage0_13[45]},
      {stage1_15[6],stage1_14[14],stage1_13[20],stage1_12[37],stage1_11[50]}
   );
   gpc615_5 gpc124 (
      {stage0_11[103], stage0_11[104], stage0_11[105], stage0_11[106], stage0_11[107]},
      {stage0_12[35]},
      {stage0_13[46], stage0_13[47], stage0_13[48], stage0_13[49], stage0_13[50], stage0_13[51]},
      {stage1_15[7],stage1_14[15],stage1_13[21],stage1_12[38],stage1_11[51]}
   );
   gpc615_5 gpc125 (
      {stage0_11[108], stage0_11[109], stage0_11[110], stage0_11[111], stage0_11[112]},
      {stage0_12[36]},
      {stage0_13[52], stage0_13[53], stage0_13[54], stage0_13[55], stage0_13[56], stage0_13[57]},
      {stage1_15[8],stage1_14[16],stage1_13[22],stage1_12[39],stage1_11[52]}
   );
   gpc615_5 gpc126 (
      {stage0_11[113], stage0_11[114], stage0_11[115], stage0_11[116], stage0_11[117]},
      {stage0_12[37]},
      {stage0_13[58], stage0_13[59], stage0_13[60], stage0_13[61], stage0_13[62], stage0_13[63]},
      {stage1_15[9],stage1_14[17],stage1_13[23],stage1_12[40],stage1_11[53]}
   );
   gpc1406_5 gpc127 (
      {stage0_12[38], stage0_12[39], stage0_12[40], stage0_12[41], stage0_12[42], stage0_12[43]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3]},
      {stage0_15[0]},
      {stage1_16[0],stage1_15[10],stage1_14[18],stage1_13[24],stage1_12[41]}
   );
   gpc606_5 gpc128 (
      {stage0_12[44], stage0_12[45], stage0_12[46], stage0_12[47], stage0_12[48], stage0_12[49]},
      {stage0_14[4], stage0_14[5], stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9]},
      {stage1_16[1],stage1_15[11],stage1_14[19],stage1_13[25],stage1_12[42]}
   );
   gpc606_5 gpc129 (
      {stage0_12[50], stage0_12[51], stage0_12[52], stage0_12[53], stage0_12[54], stage0_12[55]},
      {stage0_14[10], stage0_14[11], stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15]},
      {stage1_16[2],stage1_15[12],stage1_14[20],stage1_13[26],stage1_12[43]}
   );
   gpc606_5 gpc130 (
      {stage0_12[56], stage0_12[57], stage0_12[58], stage0_12[59], stage0_12[60], stage0_12[61]},
      {stage0_14[16], stage0_14[17], stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21]},
      {stage1_16[3],stage1_15[13],stage1_14[21],stage1_13[27],stage1_12[44]}
   );
   gpc606_5 gpc131 (
      {stage0_12[62], stage0_12[63], stage0_12[64], stage0_12[65], stage0_12[66], stage0_12[67]},
      {stage0_14[22], stage0_14[23], stage0_14[24], stage0_14[25], stage0_14[26], stage0_14[27]},
      {stage1_16[4],stage1_15[14],stage1_14[22],stage1_13[28],stage1_12[45]}
   );
   gpc606_5 gpc132 (
      {stage0_12[68], stage0_12[69], stage0_12[70], stage0_12[71], stage0_12[72], stage0_12[73]},
      {stage0_14[28], stage0_14[29], stage0_14[30], stage0_14[31], stage0_14[32], stage0_14[33]},
      {stage1_16[5],stage1_15[15],stage1_14[23],stage1_13[29],stage1_12[46]}
   );
   gpc606_5 gpc133 (
      {stage0_12[74], stage0_12[75], stage0_12[76], stage0_12[77], stage0_12[78], stage0_12[79]},
      {stage0_14[34], stage0_14[35], stage0_14[36], stage0_14[37], stage0_14[38], stage0_14[39]},
      {stage1_16[6],stage1_15[16],stage1_14[24],stage1_13[30],stage1_12[47]}
   );
   gpc606_5 gpc134 (
      {stage0_12[80], stage0_12[81], stage0_12[82], stage0_12[83], stage0_12[84], stage0_12[85]},
      {stage0_14[40], stage0_14[41], stage0_14[42], stage0_14[43], stage0_14[44], stage0_14[45]},
      {stage1_16[7],stage1_15[17],stage1_14[25],stage1_13[31],stage1_12[48]}
   );
   gpc606_5 gpc135 (
      {stage0_12[86], stage0_12[87], stage0_12[88], stage0_12[89], stage0_12[90], stage0_12[91]},
      {stage0_14[46], stage0_14[47], stage0_14[48], stage0_14[49], stage0_14[50], stage0_14[51]},
      {stage1_16[8],stage1_15[18],stage1_14[26],stage1_13[32],stage1_12[49]}
   );
   gpc606_5 gpc136 (
      {stage0_12[92], stage0_12[93], stage0_12[94], stage0_12[95], stage0_12[96], stage0_12[97]},
      {stage0_14[52], stage0_14[53], stage0_14[54], stage0_14[55], stage0_14[56], stage0_14[57]},
      {stage1_16[9],stage1_15[19],stage1_14[27],stage1_13[33],stage1_12[50]}
   );
   gpc606_5 gpc137 (
      {stage0_12[98], stage0_12[99], stage0_12[100], stage0_12[101], stage0_12[102], stage0_12[103]},
      {stage0_14[58], stage0_14[59], stage0_14[60], stage0_14[61], stage0_14[62], stage0_14[63]},
      {stage1_16[10],stage1_15[20],stage1_14[28],stage1_13[34],stage1_12[51]}
   );
   gpc606_5 gpc138 (
      {stage0_12[104], stage0_12[105], stage0_12[106], stage0_12[107], stage0_12[108], stage0_12[109]},
      {stage0_14[64], stage0_14[65], stage0_14[66], stage0_14[67], stage0_14[68], stage0_14[69]},
      {stage1_16[11],stage1_15[21],stage1_14[29],stage1_13[35],stage1_12[52]}
   );
   gpc606_5 gpc139 (
      {stage0_12[110], stage0_12[111], stage0_12[112], stage0_12[113], stage0_12[114], stage0_12[115]},
      {stage0_14[70], stage0_14[71], stage0_14[72], stage0_14[73], stage0_14[74], stage0_14[75]},
      {stage1_16[12],stage1_15[22],stage1_14[30],stage1_13[36],stage1_12[53]}
   );
   gpc606_5 gpc140 (
      {stage0_12[116], stage0_12[117], stage0_12[118], stage0_12[119], stage0_12[120], stage0_12[121]},
      {stage0_14[76], stage0_14[77], stage0_14[78], stage0_14[79], stage0_14[80], stage0_14[81]},
      {stage1_16[13],stage1_15[23],stage1_14[31],stage1_13[37],stage1_12[54]}
   );
   gpc606_5 gpc141 (
      {stage0_12[122], stage0_12[123], stage0_12[124], stage0_12[125], stage0_12[126], stage0_12[127]},
      {stage0_14[82], stage0_14[83], stage0_14[84], stage0_14[85], stage0_14[86], stage0_14[87]},
      {stage1_16[14],stage1_15[24],stage1_14[32],stage1_13[38],stage1_12[55]}
   );
   gpc606_5 gpc142 (
      {stage0_13[64], stage0_13[65], stage0_13[66], stage0_13[67], stage0_13[68], stage0_13[69]},
      {stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5], stage0_15[6]},
      {stage1_17[0],stage1_16[15],stage1_15[25],stage1_14[33],stage1_13[39]}
   );
   gpc606_5 gpc143 (
      {stage0_13[70], stage0_13[71], stage0_13[72], stage0_13[73], stage0_13[74], stage0_13[75]},
      {stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11], stage0_15[12]},
      {stage1_17[1],stage1_16[16],stage1_15[26],stage1_14[34],stage1_13[40]}
   );
   gpc606_5 gpc144 (
      {stage0_13[76], stage0_13[77], stage0_13[78], stage0_13[79], stage0_13[80], stage0_13[81]},
      {stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17], stage0_15[18]},
      {stage1_17[2],stage1_16[17],stage1_15[27],stage1_14[35],stage1_13[41]}
   );
   gpc606_5 gpc145 (
      {stage0_13[82], stage0_13[83], stage0_13[84], stage0_13[85], stage0_13[86], stage0_13[87]},
      {stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23], stage0_15[24]},
      {stage1_17[3],stage1_16[18],stage1_15[28],stage1_14[36],stage1_13[42]}
   );
   gpc606_5 gpc146 (
      {stage0_13[88], stage0_13[89], stage0_13[90], stage0_13[91], stage0_13[92], stage0_13[93]},
      {stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28], stage0_15[29], stage0_15[30]},
      {stage1_17[4],stage1_16[19],stage1_15[29],stage1_14[37],stage1_13[43]}
   );
   gpc615_5 gpc147 (
      {stage0_13[94], stage0_13[95], stage0_13[96], stage0_13[97], stage0_13[98]},
      {stage0_14[88]},
      {stage0_15[31], stage0_15[32], stage0_15[33], stage0_15[34], stage0_15[35], stage0_15[36]},
      {stage1_17[5],stage1_16[20],stage1_15[30],stage1_14[38],stage1_13[44]}
   );
   gpc615_5 gpc148 (
      {stage0_13[99], stage0_13[100], stage0_13[101], stage0_13[102], stage0_13[103]},
      {stage0_14[89]},
      {stage0_15[37], stage0_15[38], stage0_15[39], stage0_15[40], stage0_15[41], stage0_15[42]},
      {stage1_17[6],stage1_16[21],stage1_15[31],stage1_14[39],stage1_13[45]}
   );
   gpc615_5 gpc149 (
      {stage0_13[104], stage0_13[105], stage0_13[106], stage0_13[107], stage0_13[108]},
      {stage0_14[90]},
      {stage0_15[43], stage0_15[44], stage0_15[45], stage0_15[46], stage0_15[47], stage0_15[48]},
      {stage1_17[7],stage1_16[22],stage1_15[32],stage1_14[40],stage1_13[46]}
   );
   gpc615_5 gpc150 (
      {stage0_13[109], stage0_13[110], stage0_13[111], stage0_13[112], stage0_13[113]},
      {stage0_14[91]},
      {stage0_15[49], stage0_15[50], stage0_15[51], stage0_15[52], stage0_15[53], stage0_15[54]},
      {stage1_17[8],stage1_16[23],stage1_15[33],stage1_14[41],stage1_13[47]}
   );
   gpc615_5 gpc151 (
      {stage0_13[114], stage0_13[115], stage0_13[116], stage0_13[117], stage0_13[118]},
      {stage0_14[92]},
      {stage0_15[55], stage0_15[56], stage0_15[57], stage0_15[58], stage0_15[59], stage0_15[60]},
      {stage1_17[9],stage1_16[24],stage1_15[34],stage1_14[42],stage1_13[48]}
   );
   gpc615_5 gpc152 (
      {stage0_13[119], stage0_13[120], stage0_13[121], stage0_13[122], stage0_13[123]},
      {stage0_14[93]},
      {stage0_15[61], stage0_15[62], stage0_15[63], stage0_15[64], stage0_15[65], stage0_15[66]},
      {stage1_17[10],stage1_16[25],stage1_15[35],stage1_14[43],stage1_13[49]}
   );
   gpc615_5 gpc153 (
      {stage0_14[94], stage0_14[95], stage0_14[96], stage0_14[97], stage0_14[98]},
      {stage0_15[67]},
      {stage0_16[0], stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5]},
      {stage1_18[0],stage1_17[11],stage1_16[26],stage1_15[36],stage1_14[44]}
   );
   gpc615_5 gpc154 (
      {stage0_14[99], stage0_14[100], stage0_14[101], stage0_14[102], stage0_14[103]},
      {stage0_15[68]},
      {stage0_16[6], stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage1_18[1],stage1_17[12],stage1_16[27],stage1_15[37],stage1_14[45]}
   );
   gpc615_5 gpc155 (
      {stage0_14[104], stage0_14[105], stage0_14[106], stage0_14[107], stage0_14[108]},
      {stage0_15[69]},
      {stage0_16[12], stage0_16[13], stage0_16[14], stage0_16[15], stage0_16[16], stage0_16[17]},
      {stage1_18[2],stage1_17[13],stage1_16[28],stage1_15[38],stage1_14[46]}
   );
   gpc1343_5 gpc156 (
      {stage0_15[70], stage0_15[71], stage0_15[72]},
      {stage0_16[18], stage0_16[19], stage0_16[20], stage0_16[21]},
      {stage0_17[0], stage0_17[1], stage0_17[2]},
      {stage0_18[0]},
      {stage1_19[0],stage1_18[3],stage1_17[14],stage1_16[29],stage1_15[39]}
   );
   gpc606_5 gpc157 (
      {stage0_15[73], stage0_15[74], stage0_15[75], stage0_15[76], stage0_15[77], stage0_15[78]},
      {stage0_17[3], stage0_17[4], stage0_17[5], stage0_17[6], stage0_17[7], stage0_17[8]},
      {stage1_19[1],stage1_18[4],stage1_17[15],stage1_16[30],stage1_15[40]}
   );
   gpc606_5 gpc158 (
      {stage0_15[79], stage0_15[80], stage0_15[81], stage0_15[82], stage0_15[83], stage0_15[84]},
      {stage0_17[9], stage0_17[10], stage0_17[11], stage0_17[12], stage0_17[13], stage0_17[14]},
      {stage1_19[2],stage1_18[5],stage1_17[16],stage1_16[31],stage1_15[41]}
   );
   gpc606_5 gpc159 (
      {stage0_15[85], stage0_15[86], stage0_15[87], stage0_15[88], stage0_15[89], stage0_15[90]},
      {stage0_17[15], stage0_17[16], stage0_17[17], stage0_17[18], stage0_17[19], stage0_17[20]},
      {stage1_19[3],stage1_18[6],stage1_17[17],stage1_16[32],stage1_15[42]}
   );
   gpc615_5 gpc160 (
      {stage0_15[91], stage0_15[92], stage0_15[93], stage0_15[94], stage0_15[95]},
      {stage0_16[22]},
      {stage0_17[21], stage0_17[22], stage0_17[23], stage0_17[24], stage0_17[25], stage0_17[26]},
      {stage1_19[4],stage1_18[7],stage1_17[18],stage1_16[33],stage1_15[43]}
   );
   gpc615_5 gpc161 (
      {stage0_15[96], stage0_15[97], stage0_15[98], stage0_15[99], stage0_15[100]},
      {stage0_16[23]},
      {stage0_17[27], stage0_17[28], stage0_17[29], stage0_17[30], stage0_17[31], stage0_17[32]},
      {stage1_19[5],stage1_18[8],stage1_17[19],stage1_16[34],stage1_15[44]}
   );
   gpc615_5 gpc162 (
      {stage0_15[101], stage0_15[102], stage0_15[103], stage0_15[104], stage0_15[105]},
      {stage0_16[24]},
      {stage0_17[33], stage0_17[34], stage0_17[35], stage0_17[36], stage0_17[37], stage0_17[38]},
      {stage1_19[6],stage1_18[9],stage1_17[20],stage1_16[35],stage1_15[45]}
   );
   gpc606_5 gpc163 (
      {stage0_16[25], stage0_16[26], stage0_16[27], stage0_16[28], stage0_16[29], stage0_16[30]},
      {stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5], stage0_18[6]},
      {stage1_20[0],stage1_19[7],stage1_18[10],stage1_17[21],stage1_16[36]}
   );
   gpc606_5 gpc164 (
      {stage0_16[31], stage0_16[32], stage0_16[33], stage0_16[34], stage0_16[35], stage0_16[36]},
      {stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11], stage0_18[12]},
      {stage1_20[1],stage1_19[8],stage1_18[11],stage1_17[22],stage1_16[37]}
   );
   gpc606_5 gpc165 (
      {stage0_16[37], stage0_16[38], stage0_16[39], stage0_16[40], stage0_16[41], stage0_16[42]},
      {stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17], stage0_18[18]},
      {stage1_20[2],stage1_19[9],stage1_18[12],stage1_17[23],stage1_16[38]}
   );
   gpc606_5 gpc166 (
      {stage0_16[43], stage0_16[44], stage0_16[45], stage0_16[46], stage0_16[47], stage0_16[48]},
      {stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23], stage0_18[24]},
      {stage1_20[3],stage1_19[10],stage1_18[13],stage1_17[24],stage1_16[39]}
   );
   gpc606_5 gpc167 (
      {stage0_16[49], stage0_16[50], stage0_16[51], stage0_16[52], stage0_16[53], stage0_16[54]},
      {stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28], stage0_18[29], stage0_18[30]},
      {stage1_20[4],stage1_19[11],stage1_18[14],stage1_17[25],stage1_16[40]}
   );
   gpc606_5 gpc168 (
      {stage0_16[55], stage0_16[56], stage0_16[57], stage0_16[58], stage0_16[59], stage0_16[60]},
      {stage0_18[31], stage0_18[32], stage0_18[33], stage0_18[34], stage0_18[35], stage0_18[36]},
      {stage1_20[5],stage1_19[12],stage1_18[15],stage1_17[26],stage1_16[41]}
   );
   gpc606_5 gpc169 (
      {stage0_16[61], stage0_16[62], stage0_16[63], stage0_16[64], stage0_16[65], stage0_16[66]},
      {stage0_18[37], stage0_18[38], stage0_18[39], stage0_18[40], stage0_18[41], stage0_18[42]},
      {stage1_20[6],stage1_19[13],stage1_18[16],stage1_17[27],stage1_16[42]}
   );
   gpc606_5 gpc170 (
      {stage0_16[67], stage0_16[68], stage0_16[69], stage0_16[70], stage0_16[71], stage0_16[72]},
      {stage0_18[43], stage0_18[44], stage0_18[45], stage0_18[46], stage0_18[47], stage0_18[48]},
      {stage1_20[7],stage1_19[14],stage1_18[17],stage1_17[28],stage1_16[43]}
   );
   gpc606_5 gpc171 (
      {stage0_16[73], stage0_16[74], stage0_16[75], stage0_16[76], stage0_16[77], stage0_16[78]},
      {stage0_18[49], stage0_18[50], stage0_18[51], stage0_18[52], stage0_18[53], stage0_18[54]},
      {stage1_20[8],stage1_19[15],stage1_18[18],stage1_17[29],stage1_16[44]}
   );
   gpc606_5 gpc172 (
      {stage0_16[79], stage0_16[80], stage0_16[81], stage0_16[82], stage0_16[83], stage0_16[84]},
      {stage0_18[55], stage0_18[56], stage0_18[57], stage0_18[58], stage0_18[59], stage0_18[60]},
      {stage1_20[9],stage1_19[16],stage1_18[19],stage1_17[30],stage1_16[45]}
   );
   gpc606_5 gpc173 (
      {stage0_17[39], stage0_17[40], stage0_17[41], stage0_17[42], stage0_17[43], stage0_17[44]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[10],stage1_19[17],stage1_18[20],stage1_17[31]}
   );
   gpc606_5 gpc174 (
      {stage0_17[45], stage0_17[46], stage0_17[47], stage0_17[48], stage0_17[49], stage0_17[50]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[11],stage1_19[18],stage1_18[21],stage1_17[32]}
   );
   gpc606_5 gpc175 (
      {stage0_17[51], stage0_17[52], stage0_17[53], stage0_17[54], stage0_17[55], stage0_17[56]},
      {stage0_19[12], stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage1_21[2],stage1_20[12],stage1_19[19],stage1_18[22],stage1_17[33]}
   );
   gpc606_5 gpc176 (
      {stage0_17[57], stage0_17[58], stage0_17[59], stage0_17[60], stage0_17[61], stage0_17[62]},
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22], stage0_19[23]},
      {stage1_21[3],stage1_20[13],stage1_19[20],stage1_18[23],stage1_17[34]}
   );
   gpc606_5 gpc177 (
      {stage0_17[63], stage0_17[64], stage0_17[65], stage0_17[66], stage0_17[67], stage0_17[68]},
      {stage0_19[24], stage0_19[25], stage0_19[26], stage0_19[27], stage0_19[28], stage0_19[29]},
      {stage1_21[4],stage1_20[14],stage1_19[21],stage1_18[24],stage1_17[35]}
   );
   gpc606_5 gpc178 (
      {stage0_17[69], stage0_17[70], stage0_17[71], stage0_17[72], stage0_17[73], stage0_17[74]},
      {stage0_19[30], stage0_19[31], stage0_19[32], stage0_19[33], stage0_19[34], stage0_19[35]},
      {stage1_21[5],stage1_20[15],stage1_19[22],stage1_18[25],stage1_17[36]}
   );
   gpc606_5 gpc179 (
      {stage0_17[75], stage0_17[76], stage0_17[77], stage0_17[78], stage0_17[79], stage0_17[80]},
      {stage0_19[36], stage0_19[37], stage0_19[38], stage0_19[39], stage0_19[40], stage0_19[41]},
      {stage1_21[6],stage1_20[16],stage1_19[23],stage1_18[26],stage1_17[37]}
   );
   gpc606_5 gpc180 (
      {stage0_17[81], stage0_17[82], stage0_17[83], stage0_17[84], stage0_17[85], stage0_17[86]},
      {stage0_19[42], stage0_19[43], stage0_19[44], stage0_19[45], stage0_19[46], stage0_19[47]},
      {stage1_21[7],stage1_20[17],stage1_19[24],stage1_18[27],stage1_17[38]}
   );
   gpc606_5 gpc181 (
      {stage0_17[87], stage0_17[88], stage0_17[89], stage0_17[90], stage0_17[91], stage0_17[92]},
      {stage0_19[48], stage0_19[49], stage0_19[50], stage0_19[51], stage0_19[52], stage0_19[53]},
      {stage1_21[8],stage1_20[18],stage1_19[25],stage1_18[28],stage1_17[39]}
   );
   gpc615_5 gpc182 (
      {stage0_17[93], stage0_17[94], stage0_17[95], stage0_17[96], stage0_17[97]},
      {stage0_18[61]},
      {stage0_19[54], stage0_19[55], stage0_19[56], stage0_19[57], stage0_19[58], stage0_19[59]},
      {stage1_21[9],stage1_20[19],stage1_19[26],stage1_18[29],stage1_17[40]}
   );
   gpc615_5 gpc183 (
      {stage0_17[98], stage0_17[99], stage0_17[100], stage0_17[101], stage0_17[102]},
      {stage0_18[62]},
      {stage0_19[60], stage0_19[61], stage0_19[62], stage0_19[63], stage0_19[64], stage0_19[65]},
      {stage1_21[10],stage1_20[20],stage1_19[27],stage1_18[30],stage1_17[41]}
   );
   gpc606_5 gpc184 (
      {stage0_18[63], stage0_18[64], stage0_18[65], stage0_18[66], stage0_18[67], stage0_18[68]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3], stage0_20[4], stage0_20[5]},
      {stage1_22[0],stage1_21[11],stage1_20[21],stage1_19[28],stage1_18[31]}
   );
   gpc606_5 gpc185 (
      {stage0_18[69], stage0_18[70], stage0_18[71], stage0_18[72], stage0_18[73], stage0_18[74]},
      {stage0_20[6], stage0_20[7], stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11]},
      {stage1_22[1],stage1_21[12],stage1_20[22],stage1_19[29],stage1_18[32]}
   );
   gpc606_5 gpc186 (
      {stage0_18[75], stage0_18[76], stage0_18[77], stage0_18[78], stage0_18[79], stage0_18[80]},
      {stage0_20[12], stage0_20[13], stage0_20[14], stage0_20[15], stage0_20[16], stage0_20[17]},
      {stage1_22[2],stage1_21[13],stage1_20[23],stage1_19[30],stage1_18[33]}
   );
   gpc606_5 gpc187 (
      {stage0_18[81], stage0_18[82], stage0_18[83], stage0_18[84], stage0_18[85], stage0_18[86]},
      {stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21], stage0_20[22], stage0_20[23]},
      {stage1_22[3],stage1_21[14],stage1_20[24],stage1_19[31],stage1_18[34]}
   );
   gpc606_5 gpc188 (
      {stage0_18[87], stage0_18[88], stage0_18[89], stage0_18[90], stage0_18[91], stage0_18[92]},
      {stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27], stage0_20[28], stage0_20[29]},
      {stage1_22[4],stage1_21[15],stage1_20[25],stage1_19[32],stage1_18[35]}
   );
   gpc606_5 gpc189 (
      {stage0_18[93], stage0_18[94], stage0_18[95], stage0_18[96], stage0_18[97], stage0_18[98]},
      {stage0_20[30], stage0_20[31], stage0_20[32], stage0_20[33], stage0_20[34], stage0_20[35]},
      {stage1_22[5],stage1_21[16],stage1_20[26],stage1_19[33],stage1_18[36]}
   );
   gpc606_5 gpc190 (
      {stage0_18[99], stage0_18[100], stage0_18[101], stage0_18[102], stage0_18[103], stage0_18[104]},
      {stage0_20[36], stage0_20[37], stage0_20[38], stage0_20[39], stage0_20[40], stage0_20[41]},
      {stage1_22[6],stage1_21[17],stage1_20[27],stage1_19[34],stage1_18[37]}
   );
   gpc606_5 gpc191 (
      {stage0_18[105], stage0_18[106], stage0_18[107], stage0_18[108], stage0_18[109], stage0_18[110]},
      {stage0_20[42], stage0_20[43], stage0_20[44], stage0_20[45], stage0_20[46], stage0_20[47]},
      {stage1_22[7],stage1_21[18],stage1_20[28],stage1_19[35],stage1_18[38]}
   );
   gpc606_5 gpc192 (
      {stage0_18[111], stage0_18[112], stage0_18[113], stage0_18[114], stage0_18[115], stage0_18[116]},
      {stage0_20[48], stage0_20[49], stage0_20[50], stage0_20[51], stage0_20[52], stage0_20[53]},
      {stage1_22[8],stage1_21[19],stage1_20[29],stage1_19[36],stage1_18[39]}
   );
   gpc606_5 gpc193 (
      {stage0_18[117], stage0_18[118], stage0_18[119], stage0_18[120], stage0_18[121], stage0_18[122]},
      {stage0_20[54], stage0_20[55], stage0_20[56], stage0_20[57], stage0_20[58], stage0_20[59]},
      {stage1_22[9],stage1_21[20],stage1_20[30],stage1_19[37],stage1_18[40]}
   );
   gpc615_5 gpc194 (
      {stage0_18[123], stage0_18[124], stage0_18[125], stage0_18[126], stage0_18[127]},
      {stage0_19[66]},
      {stage0_20[60], stage0_20[61], stage0_20[62], stage0_20[63], stage0_20[64], stage0_20[65]},
      {stage1_22[10],stage1_21[21],stage1_20[31],stage1_19[38],stage1_18[41]}
   );
   gpc606_5 gpc195 (
      {stage0_19[67], stage0_19[68], stage0_19[69], stage0_19[70], stage0_19[71], stage0_19[72]},
      {stage0_21[0], stage0_21[1], stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5]},
      {stage1_23[0],stage1_22[11],stage1_21[22],stage1_20[32],stage1_19[39]}
   );
   gpc615_5 gpc196 (
      {stage0_19[73], stage0_19[74], stage0_19[75], stage0_19[76], stage0_19[77]},
      {stage0_20[66]},
      {stage0_21[6], stage0_21[7], stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11]},
      {stage1_23[1],stage1_22[12],stage1_21[23],stage1_20[33],stage1_19[40]}
   );
   gpc615_5 gpc197 (
      {stage0_19[78], stage0_19[79], stage0_19[80], stage0_19[81], stage0_19[82]},
      {stage0_20[67]},
      {stage0_21[12], stage0_21[13], stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17]},
      {stage1_23[2],stage1_22[13],stage1_21[24],stage1_20[34],stage1_19[41]}
   );
   gpc615_5 gpc198 (
      {stage0_19[83], stage0_19[84], stage0_19[85], stage0_19[86], stage0_19[87]},
      {stage0_20[68]},
      {stage0_21[18], stage0_21[19], stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23]},
      {stage1_23[3],stage1_22[14],stage1_21[25],stage1_20[35],stage1_19[42]}
   );
   gpc615_5 gpc199 (
      {stage0_19[88], stage0_19[89], stage0_19[90], stage0_19[91], stage0_19[92]},
      {stage0_20[69]},
      {stage0_21[24], stage0_21[25], stage0_21[26], stage0_21[27], stage0_21[28], stage0_21[29]},
      {stage1_23[4],stage1_22[15],stage1_21[26],stage1_20[36],stage1_19[43]}
   );
   gpc615_5 gpc200 (
      {stage0_19[93], stage0_19[94], stage0_19[95], stage0_19[96], stage0_19[97]},
      {stage0_20[70]},
      {stage0_21[30], stage0_21[31], stage0_21[32], stage0_21[33], stage0_21[34], stage0_21[35]},
      {stage1_23[5],stage1_22[16],stage1_21[27],stage1_20[37],stage1_19[44]}
   );
   gpc615_5 gpc201 (
      {stage0_19[98], stage0_19[99], stage0_19[100], stage0_19[101], stage0_19[102]},
      {stage0_20[71]},
      {stage0_21[36], stage0_21[37], stage0_21[38], stage0_21[39], stage0_21[40], stage0_21[41]},
      {stage1_23[6],stage1_22[17],stage1_21[28],stage1_20[38],stage1_19[45]}
   );
   gpc615_5 gpc202 (
      {stage0_19[103], stage0_19[104], stage0_19[105], stage0_19[106], stage0_19[107]},
      {stage0_20[72]},
      {stage0_21[42], stage0_21[43], stage0_21[44], stage0_21[45], stage0_21[46], stage0_21[47]},
      {stage1_23[7],stage1_22[18],stage1_21[29],stage1_20[39],stage1_19[46]}
   );
   gpc615_5 gpc203 (
      {stage0_19[108], stage0_19[109], stage0_19[110], stage0_19[111], stage0_19[112]},
      {stage0_20[73]},
      {stage0_21[48], stage0_21[49], stage0_21[50], stage0_21[51], stage0_21[52], stage0_21[53]},
      {stage1_23[8],stage1_22[19],stage1_21[30],stage1_20[40],stage1_19[47]}
   );
   gpc615_5 gpc204 (
      {stage0_19[113], stage0_19[114], stage0_19[115], stage0_19[116], stage0_19[117]},
      {stage0_20[74]},
      {stage0_21[54], stage0_21[55], stage0_21[56], stage0_21[57], stage0_21[58], stage0_21[59]},
      {stage1_23[9],stage1_22[20],stage1_21[31],stage1_20[41],stage1_19[48]}
   );
   gpc615_5 gpc205 (
      {stage0_19[118], stage0_19[119], stage0_19[120], stage0_19[121], stage0_19[122]},
      {stage0_20[75]},
      {stage0_21[60], stage0_21[61], stage0_21[62], stage0_21[63], stage0_21[64], stage0_21[65]},
      {stage1_23[10],stage1_22[21],stage1_21[32],stage1_20[42],stage1_19[49]}
   );
   gpc606_5 gpc206 (
      {stage0_20[76], stage0_20[77], stage0_20[78], stage0_20[79], stage0_20[80], stage0_20[81]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[11],stage1_22[22],stage1_21[33],stage1_20[43]}
   );
   gpc606_5 gpc207 (
      {stage0_20[82], stage0_20[83], stage0_20[84], stage0_20[85], stage0_20[86], stage0_20[87]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[12],stage1_22[23],stage1_21[34],stage1_20[44]}
   );
   gpc606_5 gpc208 (
      {stage0_20[88], stage0_20[89], stage0_20[90], stage0_20[91], stage0_20[92], stage0_20[93]},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[13],stage1_22[24],stage1_21[35],stage1_20[45]}
   );
   gpc615_5 gpc209 (
      {stage0_20[94], stage0_20[95], stage0_20[96], stage0_20[97], stage0_20[98]},
      {stage0_21[66]},
      {stage0_22[18], stage0_22[19], stage0_22[20], stage0_22[21], stage0_22[22], stage0_22[23]},
      {stage1_24[3],stage1_23[14],stage1_22[25],stage1_21[36],stage1_20[46]}
   );
   gpc615_5 gpc210 (
      {stage0_20[99], stage0_20[100], stage0_20[101], stage0_20[102], stage0_20[103]},
      {stage0_21[67]},
      {stage0_22[24], stage0_22[25], stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29]},
      {stage1_24[4],stage1_23[15],stage1_22[26],stage1_21[37],stage1_20[47]}
   );
   gpc606_5 gpc211 (
      {stage0_21[68], stage0_21[69], stage0_21[70], stage0_21[71], stage0_21[72], stage0_21[73]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[5],stage1_23[16],stage1_22[27],stage1_21[38]}
   );
   gpc606_5 gpc212 (
      {stage0_21[74], stage0_21[75], stage0_21[76], stage0_21[77], stage0_21[78], stage0_21[79]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[6],stage1_23[17],stage1_22[28],stage1_21[39]}
   );
   gpc606_5 gpc213 (
      {stage0_21[80], stage0_21[81], stage0_21[82], stage0_21[83], stage0_21[84], stage0_21[85]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage1_25[2],stage1_24[7],stage1_23[18],stage1_22[29],stage1_21[40]}
   );
   gpc615_5 gpc214 (
      {stage0_21[86], stage0_21[87], stage0_21[88], stage0_21[89], stage0_21[90]},
      {stage0_22[30]},
      {stage0_23[18], stage0_23[19], stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23]},
      {stage1_25[3],stage1_24[8],stage1_23[19],stage1_22[30],stage1_21[41]}
   );
   gpc615_5 gpc215 (
      {stage0_21[91], stage0_21[92], stage0_21[93], stage0_21[94], stage0_21[95]},
      {stage0_22[31]},
      {stage0_23[24], stage0_23[25], stage0_23[26], stage0_23[27], stage0_23[28], stage0_23[29]},
      {stage1_25[4],stage1_24[9],stage1_23[20],stage1_22[31],stage1_21[42]}
   );
   gpc615_5 gpc216 (
      {stage0_21[96], stage0_21[97], stage0_21[98], stage0_21[99], stage0_21[100]},
      {stage0_22[32]},
      {stage0_23[30], stage0_23[31], stage0_23[32], stage0_23[33], stage0_23[34], stage0_23[35]},
      {stage1_25[5],stage1_24[10],stage1_23[21],stage1_22[32],stage1_21[43]}
   );
   gpc615_5 gpc217 (
      {stage0_21[101], stage0_21[102], stage0_21[103], stage0_21[104], stage0_21[105]},
      {stage0_22[33]},
      {stage0_23[36], stage0_23[37], stage0_23[38], stage0_23[39], stage0_23[40], stage0_23[41]},
      {stage1_25[6],stage1_24[11],stage1_23[22],stage1_22[33],stage1_21[44]}
   );
   gpc615_5 gpc218 (
      {stage0_21[106], stage0_21[107], stage0_21[108], stage0_21[109], stage0_21[110]},
      {stage0_22[34]},
      {stage0_23[42], stage0_23[43], stage0_23[44], stage0_23[45], stage0_23[46], stage0_23[47]},
      {stage1_25[7],stage1_24[12],stage1_23[23],stage1_22[34],stage1_21[45]}
   );
   gpc615_5 gpc219 (
      {stage0_21[111], stage0_21[112], stage0_21[113], stage0_21[114], stage0_21[115]},
      {stage0_22[35]},
      {stage0_23[48], stage0_23[49], stage0_23[50], stage0_23[51], stage0_23[52], stage0_23[53]},
      {stage1_25[8],stage1_24[13],stage1_23[24],stage1_22[35],stage1_21[46]}
   );
   gpc615_5 gpc220 (
      {stage0_21[116], stage0_21[117], stage0_21[118], stage0_21[119], stage0_21[120]},
      {stage0_22[36]},
      {stage0_23[54], stage0_23[55], stage0_23[56], stage0_23[57], stage0_23[58], stage0_23[59]},
      {stage1_25[9],stage1_24[14],stage1_23[25],stage1_22[36],stage1_21[47]}
   );
   gpc606_5 gpc221 (
      {stage0_22[37], stage0_22[38], stage0_22[39], stage0_22[40], stage0_22[41], stage0_22[42]},
      {stage0_24[0], stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5]},
      {stage1_26[0],stage1_25[10],stage1_24[15],stage1_23[26],stage1_22[37]}
   );
   gpc606_5 gpc222 (
      {stage0_22[43], stage0_22[44], stage0_22[45], stage0_22[46], stage0_22[47], stage0_22[48]},
      {stage0_24[6], stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11]},
      {stage1_26[1],stage1_25[11],stage1_24[16],stage1_23[27],stage1_22[38]}
   );
   gpc606_5 gpc223 (
      {stage0_22[49], stage0_22[50], stage0_22[51], stage0_22[52], stage0_22[53], stage0_22[54]},
      {stage0_24[12], stage0_24[13], stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17]},
      {stage1_26[2],stage1_25[12],stage1_24[17],stage1_23[28],stage1_22[39]}
   );
   gpc606_5 gpc224 (
      {stage0_22[55], stage0_22[56], stage0_22[57], stage0_22[58], stage0_22[59], stage0_22[60]},
      {stage0_24[18], stage0_24[19], stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23]},
      {stage1_26[3],stage1_25[13],stage1_24[18],stage1_23[29],stage1_22[40]}
   );
   gpc606_5 gpc225 (
      {stage0_22[61], stage0_22[62], stage0_22[63], stage0_22[64], stage0_22[65], stage0_22[66]},
      {stage0_24[24], stage0_24[25], stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29]},
      {stage1_26[4],stage1_25[14],stage1_24[19],stage1_23[30],stage1_22[41]}
   );
   gpc606_5 gpc226 (
      {stage0_22[67], stage0_22[68], stage0_22[69], stage0_22[70], stage0_22[71], stage0_22[72]},
      {stage0_24[30], stage0_24[31], stage0_24[32], stage0_24[33], stage0_24[34], stage0_24[35]},
      {stage1_26[5],stage1_25[15],stage1_24[20],stage1_23[31],stage1_22[42]}
   );
   gpc606_5 gpc227 (
      {stage0_22[73], stage0_22[74], stage0_22[75], stage0_22[76], stage0_22[77], stage0_22[78]},
      {stage0_24[36], stage0_24[37], stage0_24[38], stage0_24[39], stage0_24[40], stage0_24[41]},
      {stage1_26[6],stage1_25[16],stage1_24[21],stage1_23[32],stage1_22[43]}
   );
   gpc606_5 gpc228 (
      {stage0_22[79], stage0_22[80], stage0_22[81], stage0_22[82], stage0_22[83], stage0_22[84]},
      {stage0_24[42], stage0_24[43], stage0_24[44], stage0_24[45], stage0_24[46], stage0_24[47]},
      {stage1_26[7],stage1_25[17],stage1_24[22],stage1_23[33],stage1_22[44]}
   );
   gpc606_5 gpc229 (
      {stage0_22[85], stage0_22[86], stage0_22[87], stage0_22[88], stage0_22[89], stage0_22[90]},
      {stage0_24[48], stage0_24[49], stage0_24[50], stage0_24[51], stage0_24[52], stage0_24[53]},
      {stage1_26[8],stage1_25[18],stage1_24[23],stage1_23[34],stage1_22[45]}
   );
   gpc615_5 gpc230 (
      {stage0_22[91], stage0_22[92], stage0_22[93], stage0_22[94], stage0_22[95]},
      {stage0_23[60]},
      {stage0_24[54], stage0_24[55], stage0_24[56], stage0_24[57], stage0_24[58], stage0_24[59]},
      {stage1_26[9],stage1_25[19],stage1_24[24],stage1_23[35],stage1_22[46]}
   );
   gpc615_5 gpc231 (
      {stage0_22[96], stage0_22[97], stage0_22[98], stage0_22[99], stage0_22[100]},
      {stage0_23[61]},
      {stage0_24[60], stage0_24[61], stage0_24[62], stage0_24[63], stage0_24[64], stage0_24[65]},
      {stage1_26[10],stage1_25[20],stage1_24[25],stage1_23[36],stage1_22[47]}
   );
   gpc615_5 gpc232 (
      {stage0_22[101], stage0_22[102], stage0_22[103], stage0_22[104], stage0_22[105]},
      {stage0_23[62]},
      {stage0_24[66], stage0_24[67], stage0_24[68], stage0_24[69], stage0_24[70], stage0_24[71]},
      {stage1_26[11],stage1_25[21],stage1_24[26],stage1_23[37],stage1_22[48]}
   );
   gpc606_5 gpc233 (
      {stage0_23[63], stage0_23[64], stage0_23[65], stage0_23[66], stage0_23[67], stage0_23[68]},
      {stage0_25[0], stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5]},
      {stage1_27[0],stage1_26[12],stage1_25[22],stage1_24[27],stage1_23[38]}
   );
   gpc606_5 gpc234 (
      {stage0_23[69], stage0_23[70], stage0_23[71], stage0_23[72], stage0_23[73], stage0_23[74]},
      {stage0_25[6], stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage1_27[1],stage1_26[13],stage1_25[23],stage1_24[28],stage1_23[39]}
   );
   gpc606_5 gpc235 (
      {stage0_23[75], stage0_23[76], stage0_23[77], stage0_23[78], stage0_23[79], stage0_23[80]},
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16], stage0_25[17]},
      {stage1_27[2],stage1_26[14],stage1_25[24],stage1_24[29],stage1_23[40]}
   );
   gpc606_5 gpc236 (
      {stage0_23[81], stage0_23[82], stage0_23[83], stage0_23[84], stage0_23[85], stage0_23[86]},
      {stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21], stage0_25[22], stage0_25[23]},
      {stage1_27[3],stage1_26[15],stage1_25[25],stage1_24[30],stage1_23[41]}
   );
   gpc606_5 gpc237 (
      {stage0_23[87], stage0_23[88], stage0_23[89], stage0_23[90], stage0_23[91], stage0_23[92]},
      {stage0_25[24], stage0_25[25], stage0_25[26], stage0_25[27], stage0_25[28], stage0_25[29]},
      {stage1_27[4],stage1_26[16],stage1_25[26],stage1_24[31],stage1_23[42]}
   );
   gpc606_5 gpc238 (
      {stage0_23[93], stage0_23[94], stage0_23[95], stage0_23[96], stage0_23[97], stage0_23[98]},
      {stage0_25[30], stage0_25[31], stage0_25[32], stage0_25[33], stage0_25[34], stage0_25[35]},
      {stage1_27[5],stage1_26[17],stage1_25[27],stage1_24[32],stage1_23[43]}
   );
   gpc606_5 gpc239 (
      {stage0_23[99], stage0_23[100], stage0_23[101], stage0_23[102], stage0_23[103], stage0_23[104]},
      {stage0_25[36], stage0_25[37], stage0_25[38], stage0_25[39], stage0_25[40], stage0_25[41]},
      {stage1_27[6],stage1_26[18],stage1_25[28],stage1_24[33],stage1_23[44]}
   );
   gpc606_5 gpc240 (
      {stage0_23[105], stage0_23[106], stage0_23[107], stage0_23[108], stage0_23[109], stage0_23[110]},
      {stage0_25[42], stage0_25[43], stage0_25[44], stage0_25[45], stage0_25[46], stage0_25[47]},
      {stage1_27[7],stage1_26[19],stage1_25[29],stage1_24[34],stage1_23[45]}
   );
   gpc606_5 gpc241 (
      {stage0_23[111], stage0_23[112], stage0_23[113], stage0_23[114], stage0_23[115], stage0_23[116]},
      {stage0_25[48], stage0_25[49], stage0_25[50], stage0_25[51], stage0_25[52], stage0_25[53]},
      {stage1_27[8],stage1_26[20],stage1_25[30],stage1_24[35],stage1_23[46]}
   );
   gpc615_5 gpc242 (
      {stage0_23[117], stage0_23[118], stage0_23[119], stage0_23[120], stage0_23[121]},
      {stage0_24[72]},
      {stage0_25[54], stage0_25[55], stage0_25[56], stage0_25[57], stage0_25[58], stage0_25[59]},
      {stage1_27[9],stage1_26[21],stage1_25[31],stage1_24[36],stage1_23[47]}
   );
   gpc606_5 gpc243 (
      {stage0_24[73], stage0_24[74], stage0_24[75], stage0_24[76], stage0_24[77], stage0_24[78]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[10],stage1_26[22],stage1_25[32],stage1_24[37]}
   );
   gpc606_5 gpc244 (
      {stage0_24[79], stage0_24[80], stage0_24[81], stage0_24[82], stage0_24[83], stage0_24[84]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[11],stage1_26[23],stage1_25[33],stage1_24[38]}
   );
   gpc606_5 gpc245 (
      {stage0_24[85], stage0_24[86], stage0_24[87], stage0_24[88], stage0_24[89], stage0_24[90]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[12],stage1_26[24],stage1_25[34],stage1_24[39]}
   );
   gpc606_5 gpc246 (
      {stage0_24[91], stage0_24[92], stage0_24[93], stage0_24[94], stage0_24[95], stage0_24[96]},
      {stage0_26[18], stage0_26[19], stage0_26[20], stage0_26[21], stage0_26[22], stage0_26[23]},
      {stage1_28[3],stage1_27[13],stage1_26[25],stage1_25[35],stage1_24[40]}
   );
   gpc606_5 gpc247 (
      {stage0_24[97], stage0_24[98], stage0_24[99], stage0_24[100], stage0_24[101], stage0_24[102]},
      {stage0_26[24], stage0_26[25], stage0_26[26], stage0_26[27], stage0_26[28], stage0_26[29]},
      {stage1_28[4],stage1_27[14],stage1_26[26],stage1_25[36],stage1_24[41]}
   );
   gpc606_5 gpc248 (
      {stage0_24[103], stage0_24[104], stage0_24[105], stage0_24[106], stage0_24[107], stage0_24[108]},
      {stage0_26[30], stage0_26[31], stage0_26[32], stage0_26[33], stage0_26[34], stage0_26[35]},
      {stage1_28[5],stage1_27[15],stage1_26[27],stage1_25[37],stage1_24[42]}
   );
   gpc606_5 gpc249 (
      {stage0_25[60], stage0_25[61], stage0_25[62], stage0_25[63], stage0_25[64], stage0_25[65]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[6],stage1_27[16],stage1_26[28],stage1_25[38]}
   );
   gpc606_5 gpc250 (
      {stage0_25[66], stage0_25[67], stage0_25[68], stage0_25[69], stage0_25[70], stage0_25[71]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[7],stage1_27[17],stage1_26[29],stage1_25[39]}
   );
   gpc606_5 gpc251 (
      {stage0_25[72], stage0_25[73], stage0_25[74], stage0_25[75], stage0_25[76], stage0_25[77]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[8],stage1_27[18],stage1_26[30],stage1_25[40]}
   );
   gpc606_5 gpc252 (
      {stage0_25[78], stage0_25[79], stage0_25[80], stage0_25[81], stage0_25[82], stage0_25[83]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[9],stage1_27[19],stage1_26[31],stage1_25[41]}
   );
   gpc606_5 gpc253 (
      {stage0_25[84], stage0_25[85], stage0_25[86], stage0_25[87], stage0_25[88], stage0_25[89]},
      {stage0_27[24], stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29]},
      {stage1_29[4],stage1_28[10],stage1_27[20],stage1_26[32],stage1_25[42]}
   );
   gpc606_5 gpc254 (
      {stage0_25[90], stage0_25[91], stage0_25[92], stage0_25[93], stage0_25[94], stage0_25[95]},
      {stage0_27[30], stage0_27[31], stage0_27[32], stage0_27[33], stage0_27[34], stage0_27[35]},
      {stage1_29[5],stage1_28[11],stage1_27[21],stage1_26[33],stage1_25[43]}
   );
   gpc606_5 gpc255 (
      {stage0_25[96], stage0_25[97], stage0_25[98], stage0_25[99], stage0_25[100], stage0_25[101]},
      {stage0_27[36], stage0_27[37], stage0_27[38], stage0_27[39], stage0_27[40], stage0_27[41]},
      {stage1_29[6],stage1_28[12],stage1_27[22],stage1_26[34],stage1_25[44]}
   );
   gpc606_5 gpc256 (
      {stage0_25[102], stage0_25[103], stage0_25[104], stage0_25[105], stage0_25[106], stage0_25[107]},
      {stage0_27[42], stage0_27[43], stage0_27[44], stage0_27[45], stage0_27[46], stage0_27[47]},
      {stage1_29[7],stage1_28[13],stage1_27[23],stage1_26[35],stage1_25[45]}
   );
   gpc606_5 gpc257 (
      {stage0_25[108], stage0_25[109], stage0_25[110], stage0_25[111], stage0_25[112], stage0_25[113]},
      {stage0_27[48], stage0_27[49], stage0_27[50], stage0_27[51], stage0_27[52], stage0_27[53]},
      {stage1_29[8],stage1_28[14],stage1_27[24],stage1_26[36],stage1_25[46]}
   );
   gpc1163_5 gpc258 (
      {stage0_26[36], stage0_26[37], stage0_26[38]},
      {stage0_27[54], stage0_27[55], stage0_27[56], stage0_27[57], stage0_27[58], stage0_27[59]},
      {stage0_28[0]},
      {stage0_29[0]},
      {stage1_30[0],stage1_29[9],stage1_28[15],stage1_27[25],stage1_26[37]}
   );
   gpc1163_5 gpc259 (
      {stage0_26[39], stage0_26[40], stage0_26[41]},
      {stage0_27[60], stage0_27[61], stage0_27[62], stage0_27[63], stage0_27[64], stage0_27[65]},
      {stage0_28[1]},
      {stage0_29[1]},
      {stage1_30[1],stage1_29[10],stage1_28[16],stage1_27[26],stage1_26[38]}
   );
   gpc1163_5 gpc260 (
      {stage0_26[42], stage0_26[43], stage0_26[44]},
      {stage0_27[66], stage0_27[67], stage0_27[68], stage0_27[69], stage0_27[70], stage0_27[71]},
      {stage0_28[2]},
      {stage0_29[2]},
      {stage1_30[2],stage1_29[11],stage1_28[17],stage1_27[27],stage1_26[39]}
   );
   gpc1163_5 gpc261 (
      {stage0_26[45], stage0_26[46], stage0_26[47]},
      {stage0_27[72], stage0_27[73], stage0_27[74], stage0_27[75], stage0_27[76], stage0_27[77]},
      {stage0_28[3]},
      {stage0_29[3]},
      {stage1_30[3],stage1_29[12],stage1_28[18],stage1_27[28],stage1_26[40]}
   );
   gpc1163_5 gpc262 (
      {stage0_26[48], stage0_26[49], stage0_26[50]},
      {stage0_27[78], stage0_27[79], stage0_27[80], stage0_27[81], stage0_27[82], stage0_27[83]},
      {stage0_28[4]},
      {stage0_29[4]},
      {stage1_30[4],stage1_29[13],stage1_28[19],stage1_27[29],stage1_26[41]}
   );
   gpc207_4 gpc263 (
      {stage0_26[51], stage0_26[52], stage0_26[53], stage0_26[54], stage0_26[55], stage0_26[56], stage0_26[57]},
      {stage0_28[5], stage0_28[6]},
      {stage1_29[14],stage1_28[20],stage1_27[30],stage1_26[42]}
   );
   gpc606_5 gpc264 (
      {stage0_26[58], stage0_26[59], stage0_26[60], stage0_26[61], stage0_26[62], stage0_26[63]},
      {stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11], stage0_28[12]},
      {stage1_30[5],stage1_29[15],stage1_28[21],stage1_27[31],stage1_26[43]}
   );
   gpc606_5 gpc265 (
      {stage0_26[64], stage0_26[65], stage0_26[66], stage0_26[67], stage0_26[68], stage0_26[69]},
      {stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17], stage0_28[18]},
      {stage1_30[6],stage1_29[16],stage1_28[22],stage1_27[32],stage1_26[44]}
   );
   gpc606_5 gpc266 (
      {stage0_26[70], stage0_26[71], stage0_26[72], stage0_26[73], stage0_26[74], stage0_26[75]},
      {stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23], stage0_28[24]},
      {stage1_30[7],stage1_29[17],stage1_28[23],stage1_27[33],stage1_26[45]}
   );
   gpc606_5 gpc267 (
      {stage0_26[76], stage0_26[77], stage0_26[78], stage0_26[79], stage0_26[80], stage0_26[81]},
      {stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28], stage0_28[29], stage0_28[30]},
      {stage1_30[8],stage1_29[18],stage1_28[24],stage1_27[34],stage1_26[46]}
   );
   gpc606_5 gpc268 (
      {stage0_26[82], stage0_26[83], stage0_26[84], stage0_26[85], stage0_26[86], stage0_26[87]},
      {stage0_28[31], stage0_28[32], stage0_28[33], stage0_28[34], stage0_28[35], stage0_28[36]},
      {stage1_30[9],stage1_29[19],stage1_28[25],stage1_27[35],stage1_26[47]}
   );
   gpc615_5 gpc269 (
      {stage0_26[88], stage0_26[89], stage0_26[90], stage0_26[91], stage0_26[92]},
      {stage0_27[84]},
      {stage0_28[37], stage0_28[38], stage0_28[39], stage0_28[40], stage0_28[41], stage0_28[42]},
      {stage1_30[10],stage1_29[20],stage1_28[26],stage1_27[36],stage1_26[48]}
   );
   gpc2135_5 gpc270 (
      {stage0_27[85], stage0_27[86], stage0_27[87], stage0_27[88], stage0_27[89]},
      {stage0_28[43], stage0_28[44], stage0_28[45]},
      {stage0_29[5]},
      {stage0_30[0], stage0_30[1]},
      {stage1_31[0],stage1_30[11],stage1_29[21],stage1_28[27],stage1_27[37]}
   );
   gpc606_5 gpc271 (
      {stage0_27[90], stage0_27[91], stage0_27[92], stage0_27[93], stage0_27[94], stage0_27[95]},
      {stage0_29[6], stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11]},
      {stage1_31[1],stage1_30[12],stage1_29[22],stage1_28[28],stage1_27[38]}
   );
   gpc606_5 gpc272 (
      {stage0_27[96], stage0_27[97], stage0_27[98], stage0_27[99], stage0_27[100], stage0_27[101]},
      {stage0_29[12], stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage1_31[2],stage1_30[13],stage1_29[23],stage1_28[29],stage1_27[39]}
   );
   gpc606_5 gpc273 (
      {stage0_27[102], stage0_27[103], stage0_27[104], stage0_27[105], stage0_27[106], stage0_27[107]},
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22], stage0_29[23]},
      {stage1_31[3],stage1_30[14],stage1_29[24],stage1_28[30],stage1_27[40]}
   );
   gpc606_5 gpc274 (
      {stage0_27[108], stage0_27[109], stage0_27[110], stage0_27[111], stage0_27[112], stage0_27[113]},
      {stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27], stage0_29[28], stage0_29[29]},
      {stage1_31[4],stage1_30[15],stage1_29[25],stage1_28[31],stage1_27[41]}
   );
   gpc606_5 gpc275 (
      {stage0_28[46], stage0_28[47], stage0_28[48], stage0_28[49], stage0_28[50], stage0_28[51]},
      {stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5], stage0_30[6], stage0_30[7]},
      {stage1_32[0],stage1_31[5],stage1_30[16],stage1_29[26],stage1_28[32]}
   );
   gpc606_5 gpc276 (
      {stage0_28[52], stage0_28[53], stage0_28[54], stage0_28[55], stage0_28[56], stage0_28[57]},
      {stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11], stage0_30[12], stage0_30[13]},
      {stage1_32[1],stage1_31[6],stage1_30[17],stage1_29[27],stage1_28[33]}
   );
   gpc606_5 gpc277 (
      {stage0_28[58], stage0_28[59], stage0_28[60], stage0_28[61], stage0_28[62], stage0_28[63]},
      {stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17], stage0_30[18], stage0_30[19]},
      {stage1_32[2],stage1_31[7],stage1_30[18],stage1_29[28],stage1_28[34]}
   );
   gpc606_5 gpc278 (
      {stage0_28[64], stage0_28[65], stage0_28[66], stage0_28[67], stage0_28[68], stage0_28[69]},
      {stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23], stage0_30[24], stage0_30[25]},
      {stage1_32[3],stage1_31[8],stage1_30[19],stage1_29[29],stage1_28[35]}
   );
   gpc606_5 gpc279 (
      {stage0_28[70], stage0_28[71], stage0_28[72], stage0_28[73], stage0_28[74], stage0_28[75]},
      {stage0_30[26], stage0_30[27], stage0_30[28], stage0_30[29], stage0_30[30], stage0_30[31]},
      {stage1_32[4],stage1_31[9],stage1_30[20],stage1_29[30],stage1_28[36]}
   );
   gpc606_5 gpc280 (
      {stage0_28[76], stage0_28[77], stage0_28[78], stage0_28[79], stage0_28[80], stage0_28[81]},
      {stage0_30[32], stage0_30[33], stage0_30[34], stage0_30[35], stage0_30[36], stage0_30[37]},
      {stage1_32[5],stage1_31[10],stage1_30[21],stage1_29[31],stage1_28[37]}
   );
   gpc606_5 gpc281 (
      {stage0_28[82], stage0_28[83], stage0_28[84], stage0_28[85], stage0_28[86], stage0_28[87]},
      {stage0_30[38], stage0_30[39], stage0_30[40], stage0_30[41], stage0_30[42], stage0_30[43]},
      {stage1_32[6],stage1_31[11],stage1_30[22],stage1_29[32],stage1_28[38]}
   );
   gpc606_5 gpc282 (
      {stage0_28[88], stage0_28[89], stage0_28[90], stage0_28[91], stage0_28[92], stage0_28[93]},
      {stage0_30[44], stage0_30[45], stage0_30[46], stage0_30[47], stage0_30[48], stage0_30[49]},
      {stage1_32[7],stage1_31[12],stage1_30[23],stage1_29[33],stage1_28[39]}
   );
   gpc606_5 gpc283 (
      {stage0_28[94], stage0_28[95], stage0_28[96], stage0_28[97], stage0_28[98], stage0_28[99]},
      {stage0_30[50], stage0_30[51], stage0_30[52], stage0_30[53], stage0_30[54], stage0_30[55]},
      {stage1_32[8],stage1_31[13],stage1_30[24],stage1_29[34],stage1_28[40]}
   );
   gpc606_5 gpc284 (
      {stage0_28[100], stage0_28[101], stage0_28[102], stage0_28[103], stage0_28[104], stage0_28[105]},
      {stage0_30[56], stage0_30[57], stage0_30[58], stage0_30[59], stage0_30[60], stage0_30[61]},
      {stage1_32[9],stage1_31[14],stage1_30[25],stage1_29[35],stage1_28[41]}
   );
   gpc615_5 gpc285 (
      {stage0_28[106], stage0_28[107], stage0_28[108], stage0_28[109], stage0_28[110]},
      {stage0_29[30]},
      {stage0_30[62], stage0_30[63], stage0_30[64], stage0_30[65], stage0_30[66], stage0_30[67]},
      {stage1_32[10],stage1_31[15],stage1_30[26],stage1_29[36],stage1_28[42]}
   );
   gpc615_5 gpc286 (
      {stage0_28[111], stage0_28[112], stage0_28[113], stage0_28[114], stage0_28[115]},
      {stage0_29[31]},
      {stage0_30[68], stage0_30[69], stage0_30[70], stage0_30[71], stage0_30[72], stage0_30[73]},
      {stage1_32[11],stage1_31[16],stage1_30[27],stage1_29[37],stage1_28[43]}
   );
   gpc615_5 gpc287 (
      {stage0_28[116], stage0_28[117], stage0_28[118], stage0_28[119], stage0_28[120]},
      {stage0_29[32]},
      {stage0_30[74], stage0_30[75], stage0_30[76], stage0_30[77], stage0_30[78], stage0_30[79]},
      {stage1_32[12],stage1_31[17],stage1_30[28],stage1_29[38],stage1_28[44]}
   );
   gpc615_5 gpc288 (
      {stage0_28[121], stage0_28[122], stage0_28[123], stage0_28[124], stage0_28[125]},
      {stage0_29[33]},
      {stage0_30[80], stage0_30[81], stage0_30[82], stage0_30[83], stage0_30[84], stage0_30[85]},
      {stage1_32[13],stage1_31[18],stage1_30[29],stage1_29[39],stage1_28[45]}
   );
   gpc135_4 gpc289 (
      {stage0_29[34], stage0_29[35], stage0_29[36], stage0_29[37], stage0_29[38]},
      {stage0_30[86], stage0_30[87], stage0_30[88]},
      {stage0_31[0]},
      {stage1_32[14],stage1_31[19],stage1_30[30],stage1_29[40]}
   );
   gpc606_5 gpc290 (
      {stage0_29[39], stage0_29[40], stage0_29[41], stage0_29[42], stage0_29[43], stage0_29[44]},
      {stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5], stage0_31[6]},
      {stage1_33[0],stage1_32[15],stage1_31[20],stage1_30[31],stage1_29[41]}
   );
   gpc606_5 gpc291 (
      {stage0_29[45], stage0_29[46], stage0_29[47], stage0_29[48], stage0_29[49], stage0_29[50]},
      {stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11], stage0_31[12]},
      {stage1_33[1],stage1_32[16],stage1_31[21],stage1_30[32],stage1_29[42]}
   );
   gpc606_5 gpc292 (
      {stage0_29[51], stage0_29[52], stage0_29[53], stage0_29[54], stage0_29[55], stage0_29[56]},
      {stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17], stage0_31[18]},
      {stage1_33[2],stage1_32[17],stage1_31[22],stage1_30[33],stage1_29[43]}
   );
   gpc606_5 gpc293 (
      {stage0_29[57], stage0_29[58], stage0_29[59], stage0_29[60], stage0_29[61], stage0_29[62]},
      {stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23], stage0_31[24]},
      {stage1_33[3],stage1_32[18],stage1_31[23],stage1_30[34],stage1_29[44]}
   );
   gpc606_5 gpc294 (
      {stage0_29[63], stage0_29[64], stage0_29[65], stage0_29[66], stage0_29[67], stage0_29[68]},
      {stage0_31[25], stage0_31[26], stage0_31[27], stage0_31[28], stage0_31[29], stage0_31[30]},
      {stage1_33[4],stage1_32[19],stage1_31[24],stage1_30[35],stage1_29[45]}
   );
   gpc606_5 gpc295 (
      {stage0_29[69], stage0_29[70], stage0_29[71], stage0_29[72], stage0_29[73], stage0_29[74]},
      {stage0_31[31], stage0_31[32], stage0_31[33], stage0_31[34], stage0_31[35], stage0_31[36]},
      {stage1_33[5],stage1_32[20],stage1_31[25],stage1_30[36],stage1_29[46]}
   );
   gpc606_5 gpc296 (
      {stage0_29[75], stage0_29[76], stage0_29[77], stage0_29[78], stage0_29[79], stage0_29[80]},
      {stage0_31[37], stage0_31[38], stage0_31[39], stage0_31[40], stage0_31[41], stage0_31[42]},
      {stage1_33[6],stage1_32[21],stage1_31[26],stage1_30[37],stage1_29[47]}
   );
   gpc606_5 gpc297 (
      {stage0_29[81], stage0_29[82], stage0_29[83], stage0_29[84], stage0_29[85], stage0_29[86]},
      {stage0_31[43], stage0_31[44], stage0_31[45], stage0_31[46], stage0_31[47], stage0_31[48]},
      {stage1_33[7],stage1_32[22],stage1_31[27],stage1_30[38],stage1_29[48]}
   );
   gpc606_5 gpc298 (
      {stage0_29[87], stage0_29[88], stage0_29[89], stage0_29[90], stage0_29[91], stage0_29[92]},
      {stage0_31[49], stage0_31[50], stage0_31[51], stage0_31[52], stage0_31[53], stage0_31[54]},
      {stage1_33[8],stage1_32[23],stage1_31[28],stage1_30[39],stage1_29[49]}
   );
   gpc606_5 gpc299 (
      {stage0_29[93], stage0_29[94], stage0_29[95], stage0_29[96], stage0_29[97], stage0_29[98]},
      {stage0_31[55], stage0_31[56], stage0_31[57], stage0_31[58], stage0_31[59], stage0_31[60]},
      {stage1_33[9],stage1_32[24],stage1_31[29],stage1_30[40],stage1_29[50]}
   );
   gpc615_5 gpc300 (
      {stage0_30[89], stage0_30[90], stage0_30[91], stage0_30[92], stage0_30[93]},
      {stage0_31[61]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3], stage0_32[4], stage0_32[5]},
      {stage1_34[0],stage1_33[10],stage1_32[25],stage1_31[30],stage1_30[41]}
   );
   gpc615_5 gpc301 (
      {stage0_30[94], stage0_30[95], stage0_30[96], stage0_30[97], stage0_30[98]},
      {stage0_31[62]},
      {stage0_32[6], stage0_32[7], stage0_32[8], stage0_32[9], stage0_32[10], stage0_32[11]},
      {stage1_34[1],stage1_33[11],stage1_32[26],stage1_31[31],stage1_30[42]}
   );
   gpc2116_5 gpc302 (
      {stage0_31[63], stage0_31[64], stage0_31[65], stage0_31[66], stage0_31[67], stage0_31[68]},
      {stage0_32[12]},
      {stage0_33[0]},
      {stage0_34[0], stage0_34[1]},
      {stage1_35[0],stage1_34[2],stage1_33[12],stage1_32[27],stage1_31[32]}
   );
   gpc615_5 gpc303 (
      {stage0_31[69], stage0_31[70], stage0_31[71], stage0_31[72], stage0_31[73]},
      {stage0_32[13]},
      {stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5], stage0_33[6]},
      {stage1_35[1],stage1_34[3],stage1_33[13],stage1_32[28],stage1_31[33]}
   );
   gpc615_5 gpc304 (
      {stage0_31[74], stage0_31[75], stage0_31[76], stage0_31[77], stage0_31[78]},
      {stage0_32[14]},
      {stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11], stage0_33[12]},
      {stage1_35[2],stage1_34[4],stage1_33[14],stage1_32[29],stage1_31[34]}
   );
   gpc615_5 gpc305 (
      {stage0_31[79], stage0_31[80], stage0_31[81], stage0_31[82], stage0_31[83]},
      {stage0_32[15]},
      {stage0_33[13], stage0_33[14], stage0_33[15], stage0_33[16], stage0_33[17], stage0_33[18]},
      {stage1_35[3],stage1_34[5],stage1_33[15],stage1_32[30],stage1_31[35]}
   );
   gpc615_5 gpc306 (
      {stage0_31[84], stage0_31[85], stage0_31[86], stage0_31[87], stage0_31[88]},
      {stage0_32[16]},
      {stage0_33[19], stage0_33[20], stage0_33[21], stage0_33[22], stage0_33[23], stage0_33[24]},
      {stage1_35[4],stage1_34[6],stage1_33[16],stage1_32[31],stage1_31[36]}
   );
   gpc615_5 gpc307 (
      {stage0_31[89], stage0_31[90], stage0_31[91], stage0_31[92], stage0_31[93]},
      {stage0_32[17]},
      {stage0_33[25], stage0_33[26], stage0_33[27], stage0_33[28], stage0_33[29], stage0_33[30]},
      {stage1_35[5],stage1_34[7],stage1_33[17],stage1_32[32],stage1_31[37]}
   );
   gpc615_5 gpc308 (
      {stage0_31[94], stage0_31[95], stage0_31[96], stage0_31[97], stage0_31[98]},
      {stage0_32[18]},
      {stage0_33[31], stage0_33[32], stage0_33[33], stage0_33[34], stage0_33[35], stage0_33[36]},
      {stage1_35[6],stage1_34[8],stage1_33[18],stage1_32[33],stage1_31[38]}
   );
   gpc615_5 gpc309 (
      {stage0_31[99], stage0_31[100], stage0_31[101], stage0_31[102], stage0_31[103]},
      {stage0_32[19]},
      {stage0_33[37], stage0_33[38], stage0_33[39], stage0_33[40], stage0_33[41], stage0_33[42]},
      {stage1_35[7],stage1_34[9],stage1_33[19],stage1_32[34],stage1_31[39]}
   );
   gpc615_5 gpc310 (
      {stage0_31[104], stage0_31[105], stage0_31[106], stage0_31[107], stage0_31[108]},
      {stage0_32[20]},
      {stage0_33[43], stage0_33[44], stage0_33[45], stage0_33[46], stage0_33[47], stage0_33[48]},
      {stage1_35[8],stage1_34[10],stage1_33[20],stage1_32[35],stage1_31[40]}
   );
   gpc606_5 gpc311 (
      {stage0_32[21], stage0_32[22], stage0_32[23], stage0_32[24], stage0_32[25], stage0_32[26]},
      {stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5], stage0_34[6], stage0_34[7]},
      {stage1_36[0],stage1_35[9],stage1_34[11],stage1_33[21],stage1_32[36]}
   );
   gpc606_5 gpc312 (
      {stage0_32[27], stage0_32[28], stage0_32[29], stage0_32[30], stage0_32[31], stage0_32[32]},
      {stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11], stage0_34[12], stage0_34[13]},
      {stage1_36[1],stage1_35[10],stage1_34[12],stage1_33[22],stage1_32[37]}
   );
   gpc606_5 gpc313 (
      {stage0_32[33], stage0_32[34], stage0_32[35], stage0_32[36], stage0_32[37], stage0_32[38]},
      {stage0_34[14], stage0_34[15], stage0_34[16], stage0_34[17], stage0_34[18], stage0_34[19]},
      {stage1_36[2],stage1_35[11],stage1_34[13],stage1_33[23],stage1_32[38]}
   );
   gpc606_5 gpc314 (
      {stage0_32[39], stage0_32[40], stage0_32[41], stage0_32[42], stage0_32[43], stage0_32[44]},
      {stage0_34[20], stage0_34[21], stage0_34[22], stage0_34[23], stage0_34[24], stage0_34[25]},
      {stage1_36[3],stage1_35[12],stage1_34[14],stage1_33[24],stage1_32[39]}
   );
   gpc606_5 gpc315 (
      {stage0_32[45], stage0_32[46], stage0_32[47], stage0_32[48], stage0_32[49], stage0_32[50]},
      {stage0_34[26], stage0_34[27], stage0_34[28], stage0_34[29], stage0_34[30], stage0_34[31]},
      {stage1_36[4],stage1_35[13],stage1_34[15],stage1_33[25],stage1_32[40]}
   );
   gpc606_5 gpc316 (
      {stage0_32[51], stage0_32[52], stage0_32[53], stage0_32[54], stage0_32[55], stage0_32[56]},
      {stage0_34[32], stage0_34[33], stage0_34[34], stage0_34[35], stage0_34[36], stage0_34[37]},
      {stage1_36[5],stage1_35[14],stage1_34[16],stage1_33[26],stage1_32[41]}
   );
   gpc606_5 gpc317 (
      {stage0_32[57], stage0_32[58], stage0_32[59], stage0_32[60], stage0_32[61], stage0_32[62]},
      {stage0_34[38], stage0_34[39], stage0_34[40], stage0_34[41], stage0_34[42], stage0_34[43]},
      {stage1_36[6],stage1_35[15],stage1_34[17],stage1_33[27],stage1_32[42]}
   );
   gpc606_5 gpc318 (
      {stage0_32[63], stage0_32[64], stage0_32[65], stage0_32[66], stage0_32[67], stage0_32[68]},
      {stage0_34[44], stage0_34[45], stage0_34[46], stage0_34[47], stage0_34[48], stage0_34[49]},
      {stage1_36[7],stage1_35[16],stage1_34[18],stage1_33[28],stage1_32[43]}
   );
   gpc606_5 gpc319 (
      {stage0_32[69], stage0_32[70], stage0_32[71], stage0_32[72], stage0_32[73], stage0_32[74]},
      {stage0_34[50], stage0_34[51], stage0_34[52], stage0_34[53], stage0_34[54], stage0_34[55]},
      {stage1_36[8],stage1_35[17],stage1_34[19],stage1_33[29],stage1_32[44]}
   );
   gpc606_5 gpc320 (
      {stage0_32[75], stage0_32[76], stage0_32[77], stage0_32[78], stage0_32[79], stage0_32[80]},
      {stage0_34[56], stage0_34[57], stage0_34[58], stage0_34[59], stage0_34[60], stage0_34[61]},
      {stage1_36[9],stage1_35[18],stage1_34[20],stage1_33[30],stage1_32[45]}
   );
   gpc606_5 gpc321 (
      {stage0_32[81], stage0_32[82], stage0_32[83], stage0_32[84], stage0_32[85], stage0_32[86]},
      {stage0_34[62], stage0_34[63], stage0_34[64], stage0_34[65], stage0_34[66], stage0_34[67]},
      {stage1_36[10],stage1_35[19],stage1_34[21],stage1_33[31],stage1_32[46]}
   );
   gpc606_5 gpc322 (
      {stage0_32[87], stage0_32[88], stage0_32[89], stage0_32[90], stage0_32[91], stage0_32[92]},
      {stage0_34[68], stage0_34[69], stage0_34[70], stage0_34[71], stage0_34[72], stage0_34[73]},
      {stage1_36[11],stage1_35[20],stage1_34[22],stage1_33[32],stage1_32[47]}
   );
   gpc606_5 gpc323 (
      {stage0_33[49], stage0_33[50], stage0_33[51], stage0_33[52], stage0_33[53], stage0_33[54]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[12],stage1_35[21],stage1_34[23],stage1_33[33]}
   );
   gpc606_5 gpc324 (
      {stage0_33[55], stage0_33[56], stage0_33[57], stage0_33[58], stage0_33[59], stage0_33[60]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[13],stage1_35[22],stage1_34[24],stage1_33[34]}
   );
   gpc606_5 gpc325 (
      {stage0_33[61], stage0_33[62], stage0_33[63], stage0_33[64], stage0_33[65], stage0_33[66]},
      {stage0_35[12], stage0_35[13], stage0_35[14], stage0_35[15], stage0_35[16], stage0_35[17]},
      {stage1_37[2],stage1_36[14],stage1_35[23],stage1_34[25],stage1_33[35]}
   );
   gpc606_5 gpc326 (
      {stage0_33[67], stage0_33[68], stage0_33[69], stage0_33[70], stage0_33[71], stage0_33[72]},
      {stage0_35[18], stage0_35[19], stage0_35[20], stage0_35[21], stage0_35[22], stage0_35[23]},
      {stage1_37[3],stage1_36[15],stage1_35[24],stage1_34[26],stage1_33[36]}
   );
   gpc606_5 gpc327 (
      {stage0_33[73], stage0_33[74], stage0_33[75], stage0_33[76], stage0_33[77], stage0_33[78]},
      {stage0_35[24], stage0_35[25], stage0_35[26], stage0_35[27], stage0_35[28], stage0_35[29]},
      {stage1_37[4],stage1_36[16],stage1_35[25],stage1_34[27],stage1_33[37]}
   );
   gpc615_5 gpc328 (
      {stage0_33[79], stage0_33[80], stage0_33[81], stage0_33[82], stage0_33[83]},
      {stage0_34[74]},
      {stage0_35[30], stage0_35[31], stage0_35[32], stage0_35[33], stage0_35[34], stage0_35[35]},
      {stage1_37[5],stage1_36[17],stage1_35[26],stage1_34[28],stage1_33[38]}
   );
   gpc615_5 gpc329 (
      {stage0_33[84], stage0_33[85], stage0_33[86], stage0_33[87], stage0_33[88]},
      {stage0_34[75]},
      {stage0_35[36], stage0_35[37], stage0_35[38], stage0_35[39], stage0_35[40], stage0_35[41]},
      {stage1_37[6],stage1_36[18],stage1_35[27],stage1_34[29],stage1_33[39]}
   );
   gpc615_5 gpc330 (
      {stage0_33[89], stage0_33[90], stage0_33[91], stage0_33[92], stage0_33[93]},
      {stage0_34[76]},
      {stage0_35[42], stage0_35[43], stage0_35[44], stage0_35[45], stage0_35[46], stage0_35[47]},
      {stage1_37[7],stage1_36[19],stage1_35[28],stage1_34[30],stage1_33[40]}
   );
   gpc615_5 gpc331 (
      {stage0_33[94], stage0_33[95], stage0_33[96], stage0_33[97], stage0_33[98]},
      {stage0_34[77]},
      {stage0_35[48], stage0_35[49], stage0_35[50], stage0_35[51], stage0_35[52], stage0_35[53]},
      {stage1_37[8],stage1_36[20],stage1_35[29],stage1_34[31],stage1_33[41]}
   );
   gpc615_5 gpc332 (
      {stage0_33[99], stage0_33[100], stage0_33[101], stage0_33[102], stage0_33[103]},
      {stage0_34[78]},
      {stage0_35[54], stage0_35[55], stage0_35[56], stage0_35[57], stage0_35[58], stage0_35[59]},
      {stage1_37[9],stage1_36[21],stage1_35[30],stage1_34[32],stage1_33[42]}
   );
   gpc615_5 gpc333 (
      {stage0_33[104], stage0_33[105], stage0_33[106], stage0_33[107], stage0_33[108]},
      {stage0_34[79]},
      {stage0_35[60], stage0_35[61], stage0_35[62], stage0_35[63], stage0_35[64], stage0_35[65]},
      {stage1_37[10],stage1_36[22],stage1_35[31],stage1_34[33],stage1_33[43]}
   );
   gpc606_5 gpc334 (
      {stage0_34[80], stage0_34[81], stage0_34[82], stage0_34[83], stage0_34[84], stage0_34[85]},
      {stage0_36[0], stage0_36[1], stage0_36[2], stage0_36[3], stage0_36[4], stage0_36[5]},
      {stage1_38[0],stage1_37[11],stage1_36[23],stage1_35[32],stage1_34[34]}
   );
   gpc606_5 gpc335 (
      {stage0_34[86], stage0_34[87], stage0_34[88], stage0_34[89], stage0_34[90], stage0_34[91]},
      {stage0_36[6], stage0_36[7], stage0_36[8], stage0_36[9], stage0_36[10], stage0_36[11]},
      {stage1_38[1],stage1_37[12],stage1_36[24],stage1_35[33],stage1_34[35]}
   );
   gpc615_5 gpc336 (
      {stage0_34[92], stage0_34[93], stage0_34[94], stage0_34[95], stage0_34[96]},
      {stage0_35[66]},
      {stage0_36[12], stage0_36[13], stage0_36[14], stage0_36[15], stage0_36[16], stage0_36[17]},
      {stage1_38[2],stage1_37[13],stage1_36[25],stage1_35[34],stage1_34[36]}
   );
   gpc615_5 gpc337 (
      {stage0_35[67], stage0_35[68], stage0_35[69], stage0_35[70], stage0_35[71]},
      {stage0_36[18]},
      {stage0_37[0], stage0_37[1], stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5]},
      {stage1_39[0],stage1_38[3],stage1_37[14],stage1_36[26],stage1_35[35]}
   );
   gpc615_5 gpc338 (
      {stage0_35[72], stage0_35[73], stage0_35[74], stage0_35[75], stage0_35[76]},
      {stage0_36[19]},
      {stage0_37[6], stage0_37[7], stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11]},
      {stage1_39[1],stage1_38[4],stage1_37[15],stage1_36[27],stage1_35[36]}
   );
   gpc615_5 gpc339 (
      {stage0_35[77], stage0_35[78], stage0_35[79], stage0_35[80], stage0_35[81]},
      {stage0_36[20]},
      {stage0_37[12], stage0_37[13], stage0_37[14], stage0_37[15], stage0_37[16], stage0_37[17]},
      {stage1_39[2],stage1_38[5],stage1_37[16],stage1_36[28],stage1_35[37]}
   );
   gpc615_5 gpc340 (
      {stage0_35[82], stage0_35[83], stage0_35[84], stage0_35[85], stage0_35[86]},
      {stage0_36[21]},
      {stage0_37[18], stage0_37[19], stage0_37[20], stage0_37[21], stage0_37[22], stage0_37[23]},
      {stage1_39[3],stage1_38[6],stage1_37[17],stage1_36[29],stage1_35[38]}
   );
   gpc615_5 gpc341 (
      {stage0_35[87], stage0_35[88], stage0_35[89], stage0_35[90], stage0_35[91]},
      {stage0_36[22]},
      {stage0_37[24], stage0_37[25], stage0_37[26], stage0_37[27], stage0_37[28], stage0_37[29]},
      {stage1_39[4],stage1_38[7],stage1_37[18],stage1_36[30],stage1_35[39]}
   );
   gpc615_5 gpc342 (
      {stage0_35[92], stage0_35[93], stage0_35[94], stage0_35[95], stage0_35[96]},
      {stage0_36[23]},
      {stage0_37[30], stage0_37[31], stage0_37[32], stage0_37[33], stage0_37[34], stage0_37[35]},
      {stage1_39[5],stage1_38[8],stage1_37[19],stage1_36[31],stage1_35[40]}
   );
   gpc615_5 gpc343 (
      {stage0_35[97], stage0_35[98], stage0_35[99], stage0_35[100], stage0_35[101]},
      {stage0_36[24]},
      {stage0_37[36], stage0_37[37], stage0_37[38], stage0_37[39], stage0_37[40], stage0_37[41]},
      {stage1_39[6],stage1_38[9],stage1_37[20],stage1_36[32],stage1_35[41]}
   );
   gpc615_5 gpc344 (
      {stage0_35[102], stage0_35[103], stage0_35[104], stage0_35[105], stage0_35[106]},
      {stage0_36[25]},
      {stage0_37[42], stage0_37[43], stage0_37[44], stage0_37[45], stage0_37[46], stage0_37[47]},
      {stage1_39[7],stage1_38[10],stage1_37[21],stage1_36[33],stage1_35[42]}
   );
   gpc615_5 gpc345 (
      {stage0_35[107], stage0_35[108], stage0_35[109], stage0_35[110], stage0_35[111]},
      {stage0_36[26]},
      {stage0_37[48], stage0_37[49], stage0_37[50], stage0_37[51], stage0_37[52], stage0_37[53]},
      {stage1_39[8],stage1_38[11],stage1_37[22],stage1_36[34],stage1_35[43]}
   );
   gpc615_5 gpc346 (
      {stage0_35[112], stage0_35[113], stage0_35[114], stage0_35[115], stage0_35[116]},
      {stage0_36[27]},
      {stage0_37[54], stage0_37[55], stage0_37[56], stage0_37[57], stage0_37[58], stage0_37[59]},
      {stage1_39[9],stage1_38[12],stage1_37[23],stage1_36[35],stage1_35[44]}
   );
   gpc615_5 gpc347 (
      {stage0_35[117], stage0_35[118], stage0_35[119], stage0_35[120], stage0_35[121]},
      {stage0_36[28]},
      {stage0_37[60], stage0_37[61], stage0_37[62], stage0_37[63], stage0_37[64], stage0_37[65]},
      {stage1_39[10],stage1_38[13],stage1_37[24],stage1_36[36],stage1_35[45]}
   );
   gpc615_5 gpc348 (
      {stage0_35[122], stage0_35[123], stage0_35[124], stage0_35[125], stage0_35[126]},
      {stage0_36[29]},
      {stage0_37[66], stage0_37[67], stage0_37[68], stage0_37[69], stage0_37[70], stage0_37[71]},
      {stage1_39[11],stage1_38[14],stage1_37[25],stage1_36[37],stage1_35[46]}
   );
   gpc606_5 gpc349 (
      {stage0_36[30], stage0_36[31], stage0_36[32], stage0_36[33], stage0_36[34], stage0_36[35]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[12],stage1_38[15],stage1_37[26],stage1_36[38]}
   );
   gpc606_5 gpc350 (
      {stage0_36[36], stage0_36[37], stage0_36[38], stage0_36[39], stage0_36[40], stage0_36[41]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[13],stage1_38[16],stage1_37[27],stage1_36[39]}
   );
   gpc606_5 gpc351 (
      {stage0_36[42], stage0_36[43], stage0_36[44], stage0_36[45], stage0_36[46], stage0_36[47]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[14],stage1_38[17],stage1_37[28],stage1_36[40]}
   );
   gpc606_5 gpc352 (
      {stage0_36[48], stage0_36[49], stage0_36[50], stage0_36[51], stage0_36[52], stage0_36[53]},
      {stage0_38[18], stage0_38[19], stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23]},
      {stage1_40[3],stage1_39[15],stage1_38[18],stage1_37[29],stage1_36[41]}
   );
   gpc606_5 gpc353 (
      {stage0_36[54], stage0_36[55], stage0_36[56], stage0_36[57], stage0_36[58], stage0_36[59]},
      {stage0_38[24], stage0_38[25], stage0_38[26], stage0_38[27], stage0_38[28], stage0_38[29]},
      {stage1_40[4],stage1_39[16],stage1_38[19],stage1_37[30],stage1_36[42]}
   );
   gpc606_5 gpc354 (
      {stage0_36[60], stage0_36[61], stage0_36[62], stage0_36[63], stage0_36[64], stage0_36[65]},
      {stage0_38[30], stage0_38[31], stage0_38[32], stage0_38[33], stage0_38[34], stage0_38[35]},
      {stage1_40[5],stage1_39[17],stage1_38[20],stage1_37[31],stage1_36[43]}
   );
   gpc606_5 gpc355 (
      {stage0_36[66], stage0_36[67], stage0_36[68], stage0_36[69], stage0_36[70], stage0_36[71]},
      {stage0_38[36], stage0_38[37], stage0_38[38], stage0_38[39], stage0_38[40], stage0_38[41]},
      {stage1_40[6],stage1_39[18],stage1_38[21],stage1_37[32],stage1_36[44]}
   );
   gpc606_5 gpc356 (
      {stage0_36[72], stage0_36[73], stage0_36[74], stage0_36[75], stage0_36[76], stage0_36[77]},
      {stage0_38[42], stage0_38[43], stage0_38[44], stage0_38[45], stage0_38[46], stage0_38[47]},
      {stage1_40[7],stage1_39[19],stage1_38[22],stage1_37[33],stage1_36[45]}
   );
   gpc606_5 gpc357 (
      {stage0_36[78], stage0_36[79], stage0_36[80], stage0_36[81], stage0_36[82], stage0_36[83]},
      {stage0_38[48], stage0_38[49], stage0_38[50], stage0_38[51], stage0_38[52], stage0_38[53]},
      {stage1_40[8],stage1_39[20],stage1_38[23],stage1_37[34],stage1_36[46]}
   );
   gpc606_5 gpc358 (
      {stage0_36[84], stage0_36[85], stage0_36[86], stage0_36[87], stage0_36[88], stage0_36[89]},
      {stage0_38[54], stage0_38[55], stage0_38[56], stage0_38[57], stage0_38[58], stage0_38[59]},
      {stage1_40[9],stage1_39[21],stage1_38[24],stage1_37[35],stage1_36[47]}
   );
   gpc606_5 gpc359 (
      {stage0_36[90], stage0_36[91], stage0_36[92], stage0_36[93], stage0_36[94], stage0_36[95]},
      {stage0_38[60], stage0_38[61], stage0_38[62], stage0_38[63], stage0_38[64], stage0_38[65]},
      {stage1_40[10],stage1_39[22],stage1_38[25],stage1_37[36],stage1_36[48]}
   );
   gpc606_5 gpc360 (
      {stage0_36[96], stage0_36[97], stage0_36[98], stage0_36[99], stage0_36[100], stage0_36[101]},
      {stage0_38[66], stage0_38[67], stage0_38[68], stage0_38[69], stage0_38[70], stage0_38[71]},
      {stage1_40[11],stage1_39[23],stage1_38[26],stage1_37[37],stage1_36[49]}
   );
   gpc606_5 gpc361 (
      {stage0_36[102], stage0_36[103], stage0_36[104], stage0_36[105], stage0_36[106], stage0_36[107]},
      {stage0_38[72], stage0_38[73], stage0_38[74], stage0_38[75], stage0_38[76], stage0_38[77]},
      {stage1_40[12],stage1_39[24],stage1_38[27],stage1_37[38],stage1_36[50]}
   );
   gpc606_5 gpc362 (
      {stage0_36[108], stage0_36[109], stage0_36[110], stage0_36[111], stage0_36[112], stage0_36[113]},
      {stage0_38[78], stage0_38[79], stage0_38[80], stage0_38[81], stage0_38[82], stage0_38[83]},
      {stage1_40[13],stage1_39[25],stage1_38[28],stage1_37[39],stage1_36[51]}
   );
   gpc606_5 gpc363 (
      {stage0_36[114], stage0_36[115], stage0_36[116], stage0_36[117], stage0_36[118], stage0_36[119]},
      {stage0_38[84], stage0_38[85], stage0_38[86], stage0_38[87], stage0_38[88], stage0_38[89]},
      {stage1_40[14],stage1_39[26],stage1_38[29],stage1_37[40],stage1_36[52]}
   );
   gpc615_5 gpc364 (
      {stage0_38[90], stage0_38[91], stage0_38[92], stage0_38[93], stage0_38[94]},
      {stage0_39[0]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[0],stage1_40[15],stage1_39[27],stage1_38[30]}
   );
   gpc615_5 gpc365 (
      {stage0_38[95], stage0_38[96], stage0_38[97], stage0_38[98], stage0_38[99]},
      {stage0_39[1]},
      {stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11]},
      {stage1_42[1],stage1_41[1],stage1_40[16],stage1_39[28],stage1_38[31]}
   );
   gpc615_5 gpc366 (
      {stage0_38[100], stage0_38[101], stage0_38[102], stage0_38[103], stage0_38[104]},
      {stage0_39[2]},
      {stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15], stage0_40[16], stage0_40[17]},
      {stage1_42[2],stage1_41[2],stage1_40[17],stage1_39[29],stage1_38[32]}
   );
   gpc615_5 gpc367 (
      {stage0_38[105], stage0_38[106], stage0_38[107], stage0_38[108], stage0_38[109]},
      {stage0_39[3]},
      {stage0_40[18], stage0_40[19], stage0_40[20], stage0_40[21], stage0_40[22], stage0_40[23]},
      {stage1_42[3],stage1_41[3],stage1_40[18],stage1_39[30],stage1_38[33]}
   );
   gpc615_5 gpc368 (
      {stage0_38[110], stage0_38[111], stage0_38[112], stage0_38[113], stage0_38[114]},
      {stage0_39[4]},
      {stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27], stage0_40[28], stage0_40[29]},
      {stage1_42[4],stage1_41[4],stage1_40[19],stage1_39[31],stage1_38[34]}
   );
   gpc615_5 gpc369 (
      {stage0_38[115], stage0_38[116], stage0_38[117], stage0_38[118], stage0_38[119]},
      {stage0_39[5]},
      {stage0_40[30], stage0_40[31], stage0_40[32], stage0_40[33], stage0_40[34], stage0_40[35]},
      {stage1_42[5],stage1_41[5],stage1_40[20],stage1_39[32],stage1_38[35]}
   );
   gpc606_5 gpc370 (
      {stage0_39[6], stage0_39[7], stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[6],stage1_41[6],stage1_40[21],stage1_39[33]}
   );
   gpc606_5 gpc371 (
      {stage0_39[12], stage0_39[13], stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17]},
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage1_43[1],stage1_42[7],stage1_41[7],stage1_40[22],stage1_39[34]}
   );
   gpc615_5 gpc372 (
      {stage0_39[18], stage0_39[19], stage0_39[20], stage0_39[21], stage0_39[22]},
      {stage0_40[36]},
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage1_43[2],stage1_42[8],stage1_41[8],stage1_40[23],stage1_39[35]}
   );
   gpc615_5 gpc373 (
      {stage0_39[23], stage0_39[24], stage0_39[25], stage0_39[26], stage0_39[27]},
      {stage0_40[37]},
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage1_43[3],stage1_42[9],stage1_41[9],stage1_40[24],stage1_39[36]}
   );
   gpc615_5 gpc374 (
      {stage0_39[28], stage0_39[29], stage0_39[30], stage0_39[31], stage0_39[32]},
      {stage0_40[38]},
      {stage0_41[24], stage0_41[25], stage0_41[26], stage0_41[27], stage0_41[28], stage0_41[29]},
      {stage1_43[4],stage1_42[10],stage1_41[10],stage1_40[25],stage1_39[37]}
   );
   gpc615_5 gpc375 (
      {stage0_39[33], stage0_39[34], stage0_39[35], stage0_39[36], stage0_39[37]},
      {stage0_40[39]},
      {stage0_41[30], stage0_41[31], stage0_41[32], stage0_41[33], stage0_41[34], stage0_41[35]},
      {stage1_43[5],stage1_42[11],stage1_41[11],stage1_40[26],stage1_39[38]}
   );
   gpc615_5 gpc376 (
      {stage0_39[38], stage0_39[39], stage0_39[40], stage0_39[41], stage0_39[42]},
      {stage0_40[40]},
      {stage0_41[36], stage0_41[37], stage0_41[38], stage0_41[39], stage0_41[40], stage0_41[41]},
      {stage1_43[6],stage1_42[12],stage1_41[12],stage1_40[27],stage1_39[39]}
   );
   gpc615_5 gpc377 (
      {stage0_39[43], stage0_39[44], stage0_39[45], stage0_39[46], stage0_39[47]},
      {stage0_40[41]},
      {stage0_41[42], stage0_41[43], stage0_41[44], stage0_41[45], stage0_41[46], stage0_41[47]},
      {stage1_43[7],stage1_42[13],stage1_41[13],stage1_40[28],stage1_39[40]}
   );
   gpc615_5 gpc378 (
      {stage0_39[48], stage0_39[49], stage0_39[50], stage0_39[51], stage0_39[52]},
      {stage0_40[42]},
      {stage0_41[48], stage0_41[49], stage0_41[50], stage0_41[51], stage0_41[52], stage0_41[53]},
      {stage1_43[8],stage1_42[14],stage1_41[14],stage1_40[29],stage1_39[41]}
   );
   gpc615_5 gpc379 (
      {stage0_39[53], stage0_39[54], stage0_39[55], stage0_39[56], stage0_39[57]},
      {stage0_40[43]},
      {stage0_41[54], stage0_41[55], stage0_41[56], stage0_41[57], stage0_41[58], stage0_41[59]},
      {stage1_43[9],stage1_42[15],stage1_41[15],stage1_40[30],stage1_39[42]}
   );
   gpc615_5 gpc380 (
      {stage0_39[58], stage0_39[59], stage0_39[60], stage0_39[61], stage0_39[62]},
      {stage0_40[44]},
      {stage0_41[60], stage0_41[61], stage0_41[62], stage0_41[63], stage0_41[64], stage0_41[65]},
      {stage1_43[10],stage1_42[16],stage1_41[16],stage1_40[31],stage1_39[43]}
   );
   gpc615_5 gpc381 (
      {stage0_39[63], stage0_39[64], stage0_39[65], stage0_39[66], stage0_39[67]},
      {stage0_40[45]},
      {stage0_41[66], stage0_41[67], stage0_41[68], stage0_41[69], stage0_41[70], stage0_41[71]},
      {stage1_43[11],stage1_42[17],stage1_41[17],stage1_40[32],stage1_39[44]}
   );
   gpc615_5 gpc382 (
      {stage0_39[68], stage0_39[69], stage0_39[70], stage0_39[71], stage0_39[72]},
      {stage0_40[46]},
      {stage0_41[72], stage0_41[73], stage0_41[74], stage0_41[75], stage0_41[76], stage0_41[77]},
      {stage1_43[12],stage1_42[18],stage1_41[18],stage1_40[33],stage1_39[45]}
   );
   gpc615_5 gpc383 (
      {stage0_39[73], stage0_39[74], stage0_39[75], stage0_39[76], stage0_39[77]},
      {stage0_40[47]},
      {stage0_41[78], stage0_41[79], stage0_41[80], stage0_41[81], stage0_41[82], stage0_41[83]},
      {stage1_43[13],stage1_42[19],stage1_41[19],stage1_40[34],stage1_39[46]}
   );
   gpc615_5 gpc384 (
      {stage0_39[78], stage0_39[79], stage0_39[80], stage0_39[81], stage0_39[82]},
      {stage0_40[48]},
      {stage0_41[84], stage0_41[85], stage0_41[86], stage0_41[87], stage0_41[88], stage0_41[89]},
      {stage1_43[14],stage1_42[20],stage1_41[20],stage1_40[35],stage1_39[47]}
   );
   gpc1163_5 gpc385 (
      {stage0_40[49], stage0_40[50], stage0_40[51]},
      {stage0_41[90], stage0_41[91], stage0_41[92], stage0_41[93], stage0_41[94], stage0_41[95]},
      {stage0_42[0]},
      {stage0_43[0]},
      {stage1_44[0],stage1_43[15],stage1_42[21],stage1_41[21],stage1_40[36]}
   );
   gpc606_5 gpc386 (
      {stage0_40[52], stage0_40[53], stage0_40[54], stage0_40[55], stage0_40[56], stage0_40[57]},
      {stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5], stage0_42[6]},
      {stage1_44[1],stage1_43[16],stage1_42[22],stage1_41[22],stage1_40[37]}
   );
   gpc606_5 gpc387 (
      {stage0_40[58], stage0_40[59], stage0_40[60], stage0_40[61], stage0_40[62], stage0_40[63]},
      {stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11], stage0_42[12]},
      {stage1_44[2],stage1_43[17],stage1_42[23],stage1_41[23],stage1_40[38]}
   );
   gpc606_5 gpc388 (
      {stage0_40[64], stage0_40[65], stage0_40[66], stage0_40[67], stage0_40[68], stage0_40[69]},
      {stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16], stage0_42[17], stage0_42[18]},
      {stage1_44[3],stage1_43[18],stage1_42[24],stage1_41[24],stage1_40[39]}
   );
   gpc606_5 gpc389 (
      {stage0_40[70], stage0_40[71], stage0_40[72], stage0_40[73], stage0_40[74], stage0_40[75]},
      {stage0_42[19], stage0_42[20], stage0_42[21], stage0_42[22], stage0_42[23], stage0_42[24]},
      {stage1_44[4],stage1_43[19],stage1_42[25],stage1_41[25],stage1_40[40]}
   );
   gpc606_5 gpc390 (
      {stage0_40[76], stage0_40[77], stage0_40[78], stage0_40[79], stage0_40[80], stage0_40[81]},
      {stage0_42[25], stage0_42[26], stage0_42[27], stage0_42[28], stage0_42[29], stage0_42[30]},
      {stage1_44[5],stage1_43[20],stage1_42[26],stage1_41[26],stage1_40[41]}
   );
   gpc606_5 gpc391 (
      {stage0_40[82], stage0_40[83], stage0_40[84], stage0_40[85], stage0_40[86], stage0_40[87]},
      {stage0_42[31], stage0_42[32], stage0_42[33], stage0_42[34], stage0_42[35], stage0_42[36]},
      {stage1_44[6],stage1_43[21],stage1_42[27],stage1_41[27],stage1_40[42]}
   );
   gpc606_5 gpc392 (
      {stage0_40[88], stage0_40[89], stage0_40[90], stage0_40[91], stage0_40[92], stage0_40[93]},
      {stage0_42[37], stage0_42[38], stage0_42[39], stage0_42[40], stage0_42[41], stage0_42[42]},
      {stage1_44[7],stage1_43[22],stage1_42[28],stage1_41[28],stage1_40[43]}
   );
   gpc606_5 gpc393 (
      {stage0_40[94], stage0_40[95], stage0_40[96], stage0_40[97], stage0_40[98], stage0_40[99]},
      {stage0_42[43], stage0_42[44], stage0_42[45], stage0_42[46], stage0_42[47], stage0_42[48]},
      {stage1_44[8],stage1_43[23],stage1_42[29],stage1_41[29],stage1_40[44]}
   );
   gpc606_5 gpc394 (
      {stage0_40[100], stage0_40[101], stage0_40[102], stage0_40[103], stage0_40[104], stage0_40[105]},
      {stage0_42[49], stage0_42[50], stage0_42[51], stage0_42[52], stage0_42[53], stage0_42[54]},
      {stage1_44[9],stage1_43[24],stage1_42[30],stage1_41[30],stage1_40[45]}
   );
   gpc606_5 gpc395 (
      {stage0_40[106], stage0_40[107], stage0_40[108], stage0_40[109], stage0_40[110], stage0_40[111]},
      {stage0_42[55], stage0_42[56], stage0_42[57], stage0_42[58], stage0_42[59], stage0_42[60]},
      {stage1_44[10],stage1_43[25],stage1_42[31],stage1_41[31],stage1_40[46]}
   );
   gpc615_5 gpc396 (
      {stage0_41[96], stage0_41[97], stage0_41[98], stage0_41[99], stage0_41[100]},
      {stage0_42[61]},
      {stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5], stage0_43[6]},
      {stage1_45[0],stage1_44[11],stage1_43[26],stage1_42[32],stage1_41[32]}
   );
   gpc615_5 gpc397 (
      {stage0_41[101], stage0_41[102], stage0_41[103], stage0_41[104], stage0_41[105]},
      {stage0_42[62]},
      {stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11], stage0_43[12]},
      {stage1_45[1],stage1_44[12],stage1_43[27],stage1_42[33],stage1_41[33]}
   );
   gpc615_5 gpc398 (
      {stage0_41[106], stage0_41[107], stage0_41[108], stage0_41[109], stage0_41[110]},
      {stage0_42[63]},
      {stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17], stage0_43[18]},
      {stage1_45[2],stage1_44[13],stage1_43[28],stage1_42[34],stage1_41[34]}
   );
   gpc615_5 gpc399 (
      {stage0_41[111], stage0_41[112], stage0_41[113], stage0_41[114], stage0_41[115]},
      {stage0_42[64]},
      {stage0_43[19], stage0_43[20], stage0_43[21], stage0_43[22], stage0_43[23], stage0_43[24]},
      {stage1_45[3],stage1_44[14],stage1_43[29],stage1_42[35],stage1_41[35]}
   );
   gpc615_5 gpc400 (
      {stage0_41[116], stage0_41[117], stage0_41[118], stage0_41[119], stage0_41[120]},
      {stage0_42[65]},
      {stage0_43[25], stage0_43[26], stage0_43[27], stage0_43[28], stage0_43[29], stage0_43[30]},
      {stage1_45[4],stage1_44[15],stage1_43[30],stage1_42[36],stage1_41[36]}
   );
   gpc615_5 gpc401 (
      {stage0_41[121], stage0_41[122], stage0_41[123], stage0_41[124], stage0_41[125]},
      {stage0_42[66]},
      {stage0_43[31], stage0_43[32], stage0_43[33], stage0_43[34], stage0_43[35], stage0_43[36]},
      {stage1_45[5],stage1_44[16],stage1_43[31],stage1_42[37],stage1_41[37]}
   );
   gpc615_5 gpc402 (
      {stage0_42[67], stage0_42[68], stage0_42[69], stage0_42[70], stage0_42[71]},
      {stage0_43[37]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[6],stage1_44[17],stage1_43[32],stage1_42[38]}
   );
   gpc615_5 gpc403 (
      {stage0_42[72], stage0_42[73], stage0_42[74], stage0_42[75], stage0_42[76]},
      {stage0_43[38]},
      {stage0_44[6], stage0_44[7], stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11]},
      {stage1_46[1],stage1_45[7],stage1_44[18],stage1_43[33],stage1_42[39]}
   );
   gpc615_5 gpc404 (
      {stage0_42[77], stage0_42[78], stage0_42[79], stage0_42[80], stage0_42[81]},
      {stage0_43[39]},
      {stage0_44[12], stage0_44[13], stage0_44[14], stage0_44[15], stage0_44[16], stage0_44[17]},
      {stage1_46[2],stage1_45[8],stage1_44[19],stage1_43[34],stage1_42[40]}
   );
   gpc615_5 gpc405 (
      {stage0_42[82], stage0_42[83], stage0_42[84], stage0_42[85], stage0_42[86]},
      {stage0_43[40]},
      {stage0_44[18], stage0_44[19], stage0_44[20], stage0_44[21], stage0_44[22], stage0_44[23]},
      {stage1_46[3],stage1_45[9],stage1_44[20],stage1_43[35],stage1_42[41]}
   );
   gpc615_5 gpc406 (
      {stage0_42[87], stage0_42[88], stage0_42[89], stage0_42[90], stage0_42[91]},
      {stage0_43[41]},
      {stage0_44[24], stage0_44[25], stage0_44[26], stage0_44[27], stage0_44[28], stage0_44[29]},
      {stage1_46[4],stage1_45[10],stage1_44[21],stage1_43[36],stage1_42[42]}
   );
   gpc615_5 gpc407 (
      {stage0_42[92], stage0_42[93], stage0_42[94], stage0_42[95], stage0_42[96]},
      {stage0_43[42]},
      {stage0_44[30], stage0_44[31], stage0_44[32], stage0_44[33], stage0_44[34], stage0_44[35]},
      {stage1_46[5],stage1_45[11],stage1_44[22],stage1_43[37],stage1_42[43]}
   );
   gpc615_5 gpc408 (
      {stage0_42[97], stage0_42[98], stage0_42[99], stage0_42[100], stage0_42[101]},
      {stage0_43[43]},
      {stage0_44[36], stage0_44[37], stage0_44[38], stage0_44[39], stage0_44[40], stage0_44[41]},
      {stage1_46[6],stage1_45[12],stage1_44[23],stage1_43[38],stage1_42[44]}
   );
   gpc615_5 gpc409 (
      {stage0_42[102], stage0_42[103], stage0_42[104], stage0_42[105], stage0_42[106]},
      {stage0_43[44]},
      {stage0_44[42], stage0_44[43], stage0_44[44], stage0_44[45], stage0_44[46], stage0_44[47]},
      {stage1_46[7],stage1_45[13],stage1_44[24],stage1_43[39],stage1_42[45]}
   );
   gpc615_5 gpc410 (
      {stage0_42[107], stage0_42[108], stage0_42[109], stage0_42[110], stage0_42[111]},
      {stage0_43[45]},
      {stage0_44[48], stage0_44[49], stage0_44[50], stage0_44[51], stage0_44[52], stage0_44[53]},
      {stage1_46[8],stage1_45[14],stage1_44[25],stage1_43[40],stage1_42[46]}
   );
   gpc615_5 gpc411 (
      {stage0_42[112], stage0_42[113], stage0_42[114], stage0_42[115], stage0_42[116]},
      {stage0_43[46]},
      {stage0_44[54], stage0_44[55], stage0_44[56], stage0_44[57], stage0_44[58], stage0_44[59]},
      {stage1_46[9],stage1_45[15],stage1_44[26],stage1_43[41],stage1_42[47]}
   );
   gpc615_5 gpc412 (
      {stage0_42[117], stage0_42[118], stage0_42[119], stage0_42[120], stage0_42[121]},
      {stage0_43[47]},
      {stage0_44[60], stage0_44[61], stage0_44[62], stage0_44[63], stage0_44[64], stage0_44[65]},
      {stage1_46[10],stage1_45[16],stage1_44[27],stage1_43[42],stage1_42[48]}
   );
   gpc615_5 gpc413 (
      {stage0_42[122], stage0_42[123], stage0_42[124], stage0_42[125], stage0_42[126]},
      {stage0_43[48]},
      {stage0_44[66], stage0_44[67], stage0_44[68], stage0_44[69], stage0_44[70], stage0_44[71]},
      {stage1_46[11],stage1_45[17],stage1_44[28],stage1_43[43],stage1_42[49]}
   );
   gpc615_5 gpc414 (
      {stage0_43[49], stage0_43[50], stage0_43[51], stage0_43[52], stage0_43[53]},
      {stage0_44[72]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[12],stage1_45[18],stage1_44[29],stage1_43[44]}
   );
   gpc615_5 gpc415 (
      {stage0_43[54], stage0_43[55], stage0_43[56], stage0_43[57], stage0_43[58]},
      {stage0_44[73]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[13],stage1_45[19],stage1_44[30],stage1_43[45]}
   );
   gpc615_5 gpc416 (
      {stage0_43[59], stage0_43[60], stage0_43[61], stage0_43[62], stage0_43[63]},
      {stage0_44[74]},
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage1_47[2],stage1_46[14],stage1_45[20],stage1_44[31],stage1_43[46]}
   );
   gpc615_5 gpc417 (
      {stage0_43[64], stage0_43[65], stage0_43[66], stage0_43[67], stage0_43[68]},
      {stage0_44[75]},
      {stage0_45[18], stage0_45[19], stage0_45[20], stage0_45[21], stage0_45[22], stage0_45[23]},
      {stage1_47[3],stage1_46[15],stage1_45[21],stage1_44[32],stage1_43[47]}
   );
   gpc615_5 gpc418 (
      {stage0_43[69], stage0_43[70], stage0_43[71], stage0_43[72], stage0_43[73]},
      {stage0_44[76]},
      {stage0_45[24], stage0_45[25], stage0_45[26], stage0_45[27], stage0_45[28], stage0_45[29]},
      {stage1_47[4],stage1_46[16],stage1_45[22],stage1_44[33],stage1_43[48]}
   );
   gpc615_5 gpc419 (
      {stage0_43[74], stage0_43[75], stage0_43[76], stage0_43[77], stage0_43[78]},
      {stage0_44[77]},
      {stage0_45[30], stage0_45[31], stage0_45[32], stage0_45[33], stage0_45[34], stage0_45[35]},
      {stage1_47[5],stage1_46[17],stage1_45[23],stage1_44[34],stage1_43[49]}
   );
   gpc615_5 gpc420 (
      {stage0_43[79], stage0_43[80], stage0_43[81], stage0_43[82], stage0_43[83]},
      {stage0_44[78]},
      {stage0_45[36], stage0_45[37], stage0_45[38], stage0_45[39], stage0_45[40], stage0_45[41]},
      {stage1_47[6],stage1_46[18],stage1_45[24],stage1_44[35],stage1_43[50]}
   );
   gpc615_5 gpc421 (
      {stage0_43[84], stage0_43[85], stage0_43[86], stage0_43[87], stage0_43[88]},
      {stage0_44[79]},
      {stage0_45[42], stage0_45[43], stage0_45[44], stage0_45[45], stage0_45[46], stage0_45[47]},
      {stage1_47[7],stage1_46[19],stage1_45[25],stage1_44[36],stage1_43[51]}
   );
   gpc615_5 gpc422 (
      {stage0_43[89], stage0_43[90], stage0_43[91], stage0_43[92], stage0_43[93]},
      {stage0_44[80]},
      {stage0_45[48], stage0_45[49], stage0_45[50], stage0_45[51], stage0_45[52], stage0_45[53]},
      {stage1_47[8],stage1_46[20],stage1_45[26],stage1_44[37],stage1_43[52]}
   );
   gpc615_5 gpc423 (
      {stage0_43[94], stage0_43[95], stage0_43[96], stage0_43[97], stage0_43[98]},
      {stage0_44[81]},
      {stage0_45[54], stage0_45[55], stage0_45[56], stage0_45[57], stage0_45[58], stage0_45[59]},
      {stage1_47[9],stage1_46[21],stage1_45[27],stage1_44[38],stage1_43[53]}
   );
   gpc615_5 gpc424 (
      {stage0_43[99], stage0_43[100], stage0_43[101], stage0_43[102], stage0_43[103]},
      {stage0_44[82]},
      {stage0_45[60], stage0_45[61], stage0_45[62], stage0_45[63], stage0_45[64], stage0_45[65]},
      {stage1_47[10],stage1_46[22],stage1_45[28],stage1_44[39],stage1_43[54]}
   );
   gpc606_5 gpc425 (
      {stage0_44[83], stage0_44[84], stage0_44[85], stage0_44[86], stage0_44[87], stage0_44[88]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[11],stage1_46[23],stage1_45[29],stage1_44[40]}
   );
   gpc606_5 gpc426 (
      {stage0_44[89], stage0_44[90], stage0_44[91], stage0_44[92], stage0_44[93], stage0_44[94]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[12],stage1_46[24],stage1_45[30],stage1_44[41]}
   );
   gpc606_5 gpc427 (
      {stage0_44[95], stage0_44[96], stage0_44[97], stage0_44[98], stage0_44[99], stage0_44[100]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[13],stage1_46[25],stage1_45[31],stage1_44[42]}
   );
   gpc606_5 gpc428 (
      {stage0_44[101], stage0_44[102], stage0_44[103], stage0_44[104], stage0_44[105], stage0_44[106]},
      {stage0_46[18], stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage1_48[3],stage1_47[14],stage1_46[26],stage1_45[32],stage1_44[43]}
   );
   gpc606_5 gpc429 (
      {stage0_44[107], stage0_44[108], stage0_44[109], stage0_44[110], stage0_44[111], stage0_44[112]},
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28], stage0_46[29]},
      {stage1_48[4],stage1_47[15],stage1_46[27],stage1_45[33],stage1_44[44]}
   );
   gpc606_5 gpc430 (
      {stage0_44[113], stage0_44[114], stage0_44[115], stage0_44[116], stage0_44[117], stage0_44[118]},
      {stage0_46[30], stage0_46[31], stage0_46[32], stage0_46[33], stage0_46[34], stage0_46[35]},
      {stage1_48[5],stage1_47[16],stage1_46[28],stage1_45[34],stage1_44[45]}
   );
   gpc606_5 gpc431 (
      {stage0_44[119], stage0_44[120], stage0_44[121], stage0_44[122], stage0_44[123], stage0_44[124]},
      {stage0_46[36], stage0_46[37], stage0_46[38], stage0_46[39], stage0_46[40], stage0_46[41]},
      {stage1_48[6],stage1_47[17],stage1_46[29],stage1_45[35],stage1_44[46]}
   );
   gpc606_5 gpc432 (
      {stage0_45[66], stage0_45[67], stage0_45[68], stage0_45[69], stage0_45[70], stage0_45[71]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[7],stage1_47[18],stage1_46[30],stage1_45[36]}
   );
   gpc606_5 gpc433 (
      {stage0_45[72], stage0_45[73], stage0_45[74], stage0_45[75], stage0_45[76], stage0_45[77]},
      {stage0_47[6], stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11]},
      {stage1_49[1],stage1_48[8],stage1_47[19],stage1_46[31],stage1_45[37]}
   );
   gpc606_5 gpc434 (
      {stage0_45[78], stage0_45[79], stage0_45[80], stage0_45[81], stage0_45[82], stage0_45[83]},
      {stage0_47[12], stage0_47[13], stage0_47[14], stage0_47[15], stage0_47[16], stage0_47[17]},
      {stage1_49[2],stage1_48[9],stage1_47[20],stage1_46[32],stage1_45[38]}
   );
   gpc606_5 gpc435 (
      {stage0_45[84], stage0_45[85], stage0_45[86], stage0_45[87], stage0_45[88], stage0_45[89]},
      {stage0_47[18], stage0_47[19], stage0_47[20], stage0_47[21], stage0_47[22], stage0_47[23]},
      {stage1_49[3],stage1_48[10],stage1_47[21],stage1_46[33],stage1_45[39]}
   );
   gpc606_5 gpc436 (
      {stage0_45[90], stage0_45[91], stage0_45[92], stage0_45[93], stage0_45[94], stage0_45[95]},
      {stage0_47[24], stage0_47[25], stage0_47[26], stage0_47[27], stage0_47[28], stage0_47[29]},
      {stage1_49[4],stage1_48[11],stage1_47[22],stage1_46[34],stage1_45[40]}
   );
   gpc606_5 gpc437 (
      {stage0_45[96], stage0_45[97], stage0_45[98], stage0_45[99], stage0_45[100], stage0_45[101]},
      {stage0_47[30], stage0_47[31], stage0_47[32], stage0_47[33], stage0_47[34], stage0_47[35]},
      {stage1_49[5],stage1_48[12],stage1_47[23],stage1_46[35],stage1_45[41]}
   );
   gpc606_5 gpc438 (
      {stage0_45[102], stage0_45[103], stage0_45[104], stage0_45[105], stage0_45[106], stage0_45[107]},
      {stage0_47[36], stage0_47[37], stage0_47[38], stage0_47[39], stage0_47[40], stage0_47[41]},
      {stage1_49[6],stage1_48[13],stage1_47[24],stage1_46[36],stage1_45[42]}
   );
   gpc606_5 gpc439 (
      {stage0_45[108], stage0_45[109], stage0_45[110], stage0_45[111], stage0_45[112], stage0_45[113]},
      {stage0_47[42], stage0_47[43], stage0_47[44], stage0_47[45], stage0_47[46], stage0_47[47]},
      {stage1_49[7],stage1_48[14],stage1_47[25],stage1_46[37],stage1_45[43]}
   );
   gpc606_5 gpc440 (
      {stage0_46[42], stage0_46[43], stage0_46[44], stage0_46[45], stage0_46[46], stage0_46[47]},
      {stage0_48[0], stage0_48[1], stage0_48[2], stage0_48[3], stage0_48[4], stage0_48[5]},
      {stage1_50[0],stage1_49[8],stage1_48[15],stage1_47[26],stage1_46[38]}
   );
   gpc606_5 gpc441 (
      {stage0_46[48], stage0_46[49], stage0_46[50], stage0_46[51], stage0_46[52], stage0_46[53]},
      {stage0_48[6], stage0_48[7], stage0_48[8], stage0_48[9], stage0_48[10], stage0_48[11]},
      {stage1_50[1],stage1_49[9],stage1_48[16],stage1_47[27],stage1_46[39]}
   );
   gpc606_5 gpc442 (
      {stage0_46[54], stage0_46[55], stage0_46[56], stage0_46[57], stage0_46[58], stage0_46[59]},
      {stage0_48[12], stage0_48[13], stage0_48[14], stage0_48[15], stage0_48[16], stage0_48[17]},
      {stage1_50[2],stage1_49[10],stage1_48[17],stage1_47[28],stage1_46[40]}
   );
   gpc606_5 gpc443 (
      {stage0_46[60], stage0_46[61], stage0_46[62], stage0_46[63], stage0_46[64], stage0_46[65]},
      {stage0_48[18], stage0_48[19], stage0_48[20], stage0_48[21], stage0_48[22], stage0_48[23]},
      {stage1_50[3],stage1_49[11],stage1_48[18],stage1_47[29],stage1_46[41]}
   );
   gpc615_5 gpc444 (
      {stage0_46[66], stage0_46[67], stage0_46[68], stage0_46[69], stage0_46[70]},
      {stage0_47[48]},
      {stage0_48[24], stage0_48[25], stage0_48[26], stage0_48[27], stage0_48[28], stage0_48[29]},
      {stage1_50[4],stage1_49[12],stage1_48[19],stage1_47[30],stage1_46[42]}
   );
   gpc615_5 gpc445 (
      {stage0_46[71], stage0_46[72], stage0_46[73], stage0_46[74], stage0_46[75]},
      {stage0_47[49]},
      {stage0_48[30], stage0_48[31], stage0_48[32], stage0_48[33], stage0_48[34], stage0_48[35]},
      {stage1_50[5],stage1_49[13],stage1_48[20],stage1_47[31],stage1_46[43]}
   );
   gpc615_5 gpc446 (
      {stage0_46[76], stage0_46[77], stage0_46[78], stage0_46[79], stage0_46[80]},
      {stage0_47[50]},
      {stage0_48[36], stage0_48[37], stage0_48[38], stage0_48[39], stage0_48[40], stage0_48[41]},
      {stage1_50[6],stage1_49[14],stage1_48[21],stage1_47[32],stage1_46[44]}
   );
   gpc615_5 gpc447 (
      {stage0_46[81], stage0_46[82], stage0_46[83], stage0_46[84], stage0_46[85]},
      {stage0_47[51]},
      {stage0_48[42], stage0_48[43], stage0_48[44], stage0_48[45], stage0_48[46], stage0_48[47]},
      {stage1_50[7],stage1_49[15],stage1_48[22],stage1_47[33],stage1_46[45]}
   );
   gpc1325_5 gpc448 (
      {stage0_46[86], stage0_46[87], stage0_46[88], stage0_46[89], stage0_46[90]},
      {stage0_47[52], stage0_47[53]},
      {stage0_48[48], stage0_48[49], stage0_48[50]},
      {stage0_49[0]},
      {stage1_50[8],stage1_49[16],stage1_48[23],stage1_47[34],stage1_46[46]}
   );
   gpc1325_5 gpc449 (
      {stage0_46[91], stage0_46[92], stage0_46[93], stage0_46[94], stage0_46[95]},
      {stage0_47[54], stage0_47[55]},
      {stage0_48[51], stage0_48[52], stage0_48[53]},
      {stage0_49[1]},
      {stage1_50[9],stage1_49[17],stage1_48[24],stage1_47[35],stage1_46[47]}
   );
   gpc2135_5 gpc450 (
      {stage0_47[56], stage0_47[57], stage0_47[58], stage0_47[59], stage0_47[60]},
      {stage0_48[54], stage0_48[55], stage0_48[56]},
      {stage0_49[2]},
      {stage0_50[0], stage0_50[1]},
      {stage1_51[0],stage1_50[10],stage1_49[18],stage1_48[25],stage1_47[36]}
   );
   gpc606_5 gpc451 (
      {stage0_47[61], stage0_47[62], stage0_47[63], stage0_47[64], stage0_47[65], stage0_47[66]},
      {stage0_49[3], stage0_49[4], stage0_49[5], stage0_49[6], stage0_49[7], stage0_49[8]},
      {stage1_51[1],stage1_50[11],stage1_49[19],stage1_48[26],stage1_47[37]}
   );
   gpc606_5 gpc452 (
      {stage0_47[67], stage0_47[68], stage0_47[69], stage0_47[70], stage0_47[71], stage0_47[72]},
      {stage0_49[9], stage0_49[10], stage0_49[11], stage0_49[12], stage0_49[13], stage0_49[14]},
      {stage1_51[2],stage1_50[12],stage1_49[20],stage1_48[27],stage1_47[38]}
   );
   gpc615_5 gpc453 (
      {stage0_47[73], stage0_47[74], stage0_47[75], stage0_47[76], stage0_47[77]},
      {stage0_48[57]},
      {stage0_49[15], stage0_49[16], stage0_49[17], stage0_49[18], stage0_49[19], stage0_49[20]},
      {stage1_51[3],stage1_50[13],stage1_49[21],stage1_48[28],stage1_47[39]}
   );
   gpc615_5 gpc454 (
      {stage0_47[78], stage0_47[79], stage0_47[80], stage0_47[81], stage0_47[82]},
      {stage0_48[58]},
      {stage0_49[21], stage0_49[22], stage0_49[23], stage0_49[24], stage0_49[25], stage0_49[26]},
      {stage1_51[4],stage1_50[14],stage1_49[22],stage1_48[29],stage1_47[40]}
   );
   gpc615_5 gpc455 (
      {stage0_47[83], stage0_47[84], stage0_47[85], stage0_47[86], stage0_47[87]},
      {stage0_48[59]},
      {stage0_49[27], stage0_49[28], stage0_49[29], stage0_49[30], stage0_49[31], stage0_49[32]},
      {stage1_51[5],stage1_50[15],stage1_49[23],stage1_48[30],stage1_47[41]}
   );
   gpc615_5 gpc456 (
      {stage0_47[88], stage0_47[89], stage0_47[90], stage0_47[91], stage0_47[92]},
      {stage0_48[60]},
      {stage0_49[33], stage0_49[34], stage0_49[35], stage0_49[36], stage0_49[37], stage0_49[38]},
      {stage1_51[6],stage1_50[16],stage1_49[24],stage1_48[31],stage1_47[42]}
   );
   gpc615_5 gpc457 (
      {stage0_47[93], stage0_47[94], stage0_47[95], stage0_47[96], stage0_47[97]},
      {stage0_48[61]},
      {stage0_49[39], stage0_49[40], stage0_49[41], stage0_49[42], stage0_49[43], stage0_49[44]},
      {stage1_51[7],stage1_50[17],stage1_49[25],stage1_48[32],stage1_47[43]}
   );
   gpc615_5 gpc458 (
      {stage0_47[98], stage0_47[99], stage0_47[100], stage0_47[101], stage0_47[102]},
      {stage0_48[62]},
      {stage0_49[45], stage0_49[46], stage0_49[47], stage0_49[48], stage0_49[49], stage0_49[50]},
      {stage1_51[8],stage1_50[18],stage1_49[26],stage1_48[33],stage1_47[44]}
   );
   gpc606_5 gpc459 (
      {stage0_48[63], stage0_48[64], stage0_48[65], stage0_48[66], stage0_48[67], stage0_48[68]},
      {stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5], stage0_50[6], stage0_50[7]},
      {stage1_52[0],stage1_51[9],stage1_50[19],stage1_49[27],stage1_48[34]}
   );
   gpc606_5 gpc460 (
      {stage0_48[69], stage0_48[70], stage0_48[71], stage0_48[72], stage0_48[73], stage0_48[74]},
      {stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11], stage0_50[12], stage0_50[13]},
      {stage1_52[1],stage1_51[10],stage1_50[20],stage1_49[28],stage1_48[35]}
   );
   gpc606_5 gpc461 (
      {stage0_48[75], stage0_48[76], stage0_48[77], stage0_48[78], stage0_48[79], stage0_48[80]},
      {stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17], stage0_50[18], stage0_50[19]},
      {stage1_52[2],stage1_51[11],stage1_50[21],stage1_49[29],stage1_48[36]}
   );
   gpc606_5 gpc462 (
      {stage0_48[81], stage0_48[82], stage0_48[83], stage0_48[84], stage0_48[85], stage0_48[86]},
      {stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23], stage0_50[24], stage0_50[25]},
      {stage1_52[3],stage1_51[12],stage1_50[22],stage1_49[30],stage1_48[37]}
   );
   gpc606_5 gpc463 (
      {stage0_48[87], stage0_48[88], stage0_48[89], stage0_48[90], stage0_48[91], stage0_48[92]},
      {stage0_50[26], stage0_50[27], stage0_50[28], stage0_50[29], stage0_50[30], stage0_50[31]},
      {stage1_52[4],stage1_51[13],stage1_50[23],stage1_49[31],stage1_48[38]}
   );
   gpc606_5 gpc464 (
      {stage0_48[93], stage0_48[94], stage0_48[95], stage0_48[96], stage0_48[97], stage0_48[98]},
      {stage0_50[32], stage0_50[33], stage0_50[34], stage0_50[35], stage0_50[36], stage0_50[37]},
      {stage1_52[5],stage1_51[14],stage1_50[24],stage1_49[32],stage1_48[39]}
   );
   gpc606_5 gpc465 (
      {stage0_48[99], stage0_48[100], stage0_48[101], stage0_48[102], stage0_48[103], stage0_48[104]},
      {stage0_50[38], stage0_50[39], stage0_50[40], stage0_50[41], stage0_50[42], stage0_50[43]},
      {stage1_52[6],stage1_51[15],stage1_50[25],stage1_49[33],stage1_48[40]}
   );
   gpc606_5 gpc466 (
      {stage0_48[105], stage0_48[106], stage0_48[107], stage0_48[108], stage0_48[109], stage0_48[110]},
      {stage0_50[44], stage0_50[45], stage0_50[46], stage0_50[47], stage0_50[48], stage0_50[49]},
      {stage1_52[7],stage1_51[16],stage1_50[26],stage1_49[34],stage1_48[41]}
   );
   gpc606_5 gpc467 (
      {stage0_48[111], stage0_48[112], stage0_48[113], stage0_48[114], stage0_48[115], stage0_48[116]},
      {stage0_50[50], stage0_50[51], stage0_50[52], stage0_50[53], stage0_50[54], stage0_50[55]},
      {stage1_52[8],stage1_51[17],stage1_50[27],stage1_49[35],stage1_48[42]}
   );
   gpc615_5 gpc468 (
      {stage0_48[117], stage0_48[118], stage0_48[119], stage0_48[120], stage0_48[121]},
      {stage0_49[51]},
      {stage0_50[56], stage0_50[57], stage0_50[58], stage0_50[59], stage0_50[60], stage0_50[61]},
      {stage1_52[9],stage1_51[18],stage1_50[28],stage1_49[36],stage1_48[43]}
   );
   gpc615_5 gpc469 (
      {stage0_48[122], stage0_48[123], stage0_48[124], stage0_48[125], stage0_48[126]},
      {stage0_49[52]},
      {stage0_50[62], stage0_50[63], stage0_50[64], stage0_50[65], stage0_50[66], stage0_50[67]},
      {stage1_52[10],stage1_51[19],stage1_50[29],stage1_49[37],stage1_48[44]}
   );
   gpc606_5 gpc470 (
      {stage0_49[53], stage0_49[54], stage0_49[55], stage0_49[56], stage0_49[57], stage0_49[58]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[11],stage1_51[20],stage1_50[30],stage1_49[38]}
   );
   gpc606_5 gpc471 (
      {stage0_49[59], stage0_49[60], stage0_49[61], stage0_49[62], stage0_49[63], stage0_49[64]},
      {stage0_51[6], stage0_51[7], stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11]},
      {stage1_53[1],stage1_52[12],stage1_51[21],stage1_50[31],stage1_49[39]}
   );
   gpc606_5 gpc472 (
      {stage0_49[65], stage0_49[66], stage0_49[67], stage0_49[68], stage0_49[69], stage0_49[70]},
      {stage0_51[12], stage0_51[13], stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17]},
      {stage1_53[2],stage1_52[13],stage1_51[22],stage1_50[32],stage1_49[40]}
   );
   gpc606_5 gpc473 (
      {stage0_49[71], stage0_49[72], stage0_49[73], stage0_49[74], stage0_49[75], stage0_49[76]},
      {stage0_51[18], stage0_51[19], stage0_51[20], stage0_51[21], stage0_51[22], stage0_51[23]},
      {stage1_53[3],stage1_52[14],stage1_51[23],stage1_50[33],stage1_49[41]}
   );
   gpc606_5 gpc474 (
      {stage0_49[77], stage0_49[78], stage0_49[79], stage0_49[80], stage0_49[81], stage0_49[82]},
      {stage0_51[24], stage0_51[25], stage0_51[26], stage0_51[27], stage0_51[28], stage0_51[29]},
      {stage1_53[4],stage1_52[15],stage1_51[24],stage1_50[34],stage1_49[42]}
   );
   gpc606_5 gpc475 (
      {stage0_49[83], stage0_49[84], stage0_49[85], stage0_49[86], stage0_49[87], stage0_49[88]},
      {stage0_51[30], stage0_51[31], stage0_51[32], stage0_51[33], stage0_51[34], stage0_51[35]},
      {stage1_53[5],stage1_52[16],stage1_51[25],stage1_50[35],stage1_49[43]}
   );
   gpc606_5 gpc476 (
      {stage0_49[89], stage0_49[90], stage0_49[91], stage0_49[92], stage0_49[93], stage0_49[94]},
      {stage0_51[36], stage0_51[37], stage0_51[38], stage0_51[39], stage0_51[40], stage0_51[41]},
      {stage1_53[6],stage1_52[17],stage1_51[26],stage1_50[36],stage1_49[44]}
   );
   gpc606_5 gpc477 (
      {stage0_49[95], stage0_49[96], stage0_49[97], stage0_49[98], stage0_49[99], stage0_49[100]},
      {stage0_51[42], stage0_51[43], stage0_51[44], stage0_51[45], stage0_51[46], stage0_51[47]},
      {stage1_53[7],stage1_52[18],stage1_51[27],stage1_50[37],stage1_49[45]}
   );
   gpc606_5 gpc478 (
      {stage0_49[101], stage0_49[102], stage0_49[103], stage0_49[104], stage0_49[105], stage0_49[106]},
      {stage0_51[48], stage0_51[49], stage0_51[50], stage0_51[51], stage0_51[52], stage0_51[53]},
      {stage1_53[8],stage1_52[19],stage1_51[28],stage1_50[38],stage1_49[46]}
   );
   gpc606_5 gpc479 (
      {stage0_49[107], stage0_49[108], stage0_49[109], stage0_49[110], stage0_49[111], stage0_49[112]},
      {stage0_51[54], stage0_51[55], stage0_51[56], stage0_51[57], stage0_51[58], stage0_51[59]},
      {stage1_53[9],stage1_52[20],stage1_51[29],stage1_50[39],stage1_49[47]}
   );
   gpc606_5 gpc480 (
      {stage0_49[113], stage0_49[114], stage0_49[115], stage0_49[116], stage0_49[117], stage0_49[118]},
      {stage0_51[60], stage0_51[61], stage0_51[62], stage0_51[63], stage0_51[64], stage0_51[65]},
      {stage1_53[10],stage1_52[21],stage1_51[30],stage1_50[40],stage1_49[48]}
   );
   gpc606_5 gpc481 (
      {stage0_49[119], stage0_49[120], stage0_49[121], stage0_49[122], stage0_49[123], stage0_49[124]},
      {stage0_51[66], stage0_51[67], stage0_51[68], stage0_51[69], stage0_51[70], stage0_51[71]},
      {stage1_53[11],stage1_52[22],stage1_51[31],stage1_50[41],stage1_49[49]}
   );
   gpc623_5 gpc482 (
      {stage0_49[125], stage0_49[126], stage0_49[127]},
      {stage0_50[68], stage0_50[69]},
      {stage0_51[72], stage0_51[73], stage0_51[74], stage0_51[75], stage0_51[76], stage0_51[77]},
      {stage1_53[12],stage1_52[23],stage1_51[32],stage1_50[42],stage1_49[50]}
   );
   gpc606_5 gpc483 (
      {stage0_50[70], stage0_50[71], stage0_50[72], stage0_50[73], stage0_50[74], stage0_50[75]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[13],stage1_52[24],stage1_51[33],stage1_50[43]}
   );
   gpc606_5 gpc484 (
      {stage0_50[76], stage0_50[77], stage0_50[78], stage0_50[79], stage0_50[80], stage0_50[81]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[14],stage1_52[25],stage1_51[34],stage1_50[44]}
   );
   gpc606_5 gpc485 (
      {stage0_50[82], stage0_50[83], stage0_50[84], stage0_50[85], stage0_50[86], stage0_50[87]},
      {stage0_52[12], stage0_52[13], stage0_52[14], stage0_52[15], stage0_52[16], stage0_52[17]},
      {stage1_54[2],stage1_53[15],stage1_52[26],stage1_51[35],stage1_50[45]}
   );
   gpc606_5 gpc486 (
      {stage0_50[88], stage0_50[89], stage0_50[90], stage0_50[91], stage0_50[92], stage0_50[93]},
      {stage0_52[18], stage0_52[19], stage0_52[20], stage0_52[21], stage0_52[22], stage0_52[23]},
      {stage1_54[3],stage1_53[16],stage1_52[27],stage1_51[36],stage1_50[46]}
   );
   gpc606_5 gpc487 (
      {stage0_50[94], stage0_50[95], stage0_50[96], stage0_50[97], stage0_50[98], stage0_50[99]},
      {stage0_52[24], stage0_52[25], stage0_52[26], stage0_52[27], stage0_52[28], stage0_52[29]},
      {stage1_54[4],stage1_53[17],stage1_52[28],stage1_51[37],stage1_50[47]}
   );
   gpc606_5 gpc488 (
      {stage0_50[100], stage0_50[101], stage0_50[102], stage0_50[103], stage0_50[104], stage0_50[105]},
      {stage0_52[30], stage0_52[31], stage0_52[32], stage0_52[33], stage0_52[34], stage0_52[35]},
      {stage1_54[5],stage1_53[18],stage1_52[29],stage1_51[38],stage1_50[48]}
   );
   gpc606_5 gpc489 (
      {stage0_51[78], stage0_51[79], stage0_51[80], stage0_51[81], stage0_51[82], stage0_51[83]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[6],stage1_53[19],stage1_52[30],stage1_51[39]}
   );
   gpc606_5 gpc490 (
      {stage0_51[84], stage0_51[85], stage0_51[86], stage0_51[87], stage0_51[88], stage0_51[89]},
      {stage0_53[6], stage0_53[7], stage0_53[8], stage0_53[9], stage0_53[10], stage0_53[11]},
      {stage1_55[1],stage1_54[7],stage1_53[20],stage1_52[31],stage1_51[40]}
   );
   gpc606_5 gpc491 (
      {stage0_51[90], stage0_51[91], stage0_51[92], stage0_51[93], stage0_51[94], stage0_51[95]},
      {stage0_53[12], stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage1_55[2],stage1_54[8],stage1_53[21],stage1_52[32],stage1_51[41]}
   );
   gpc606_5 gpc492 (
      {stage0_51[96], stage0_51[97], stage0_51[98], stage0_51[99], stage0_51[100], stage0_51[101]},
      {stage0_53[18], stage0_53[19], stage0_53[20], stage0_53[21], stage0_53[22], stage0_53[23]},
      {stage1_55[3],stage1_54[9],stage1_53[22],stage1_52[33],stage1_51[42]}
   );
   gpc606_5 gpc493 (
      {stage0_51[102], stage0_51[103], stage0_51[104], stage0_51[105], stage0_51[106], stage0_51[107]},
      {stage0_53[24], stage0_53[25], stage0_53[26], stage0_53[27], stage0_53[28], stage0_53[29]},
      {stage1_55[4],stage1_54[10],stage1_53[23],stage1_52[34],stage1_51[43]}
   );
   gpc606_5 gpc494 (
      {stage0_51[108], stage0_51[109], stage0_51[110], stage0_51[111], stage0_51[112], stage0_51[113]},
      {stage0_53[30], stage0_53[31], stage0_53[32], stage0_53[33], stage0_53[34], stage0_53[35]},
      {stage1_55[5],stage1_54[11],stage1_53[24],stage1_52[35],stage1_51[44]}
   );
   gpc606_5 gpc495 (
      {stage0_51[114], stage0_51[115], stage0_51[116], stage0_51[117], stage0_51[118], stage0_51[119]},
      {stage0_53[36], stage0_53[37], stage0_53[38], stage0_53[39], stage0_53[40], stage0_53[41]},
      {stage1_55[6],stage1_54[12],stage1_53[25],stage1_52[36],stage1_51[45]}
   );
   gpc606_5 gpc496 (
      {stage0_51[120], stage0_51[121], stage0_51[122], stage0_51[123], stage0_51[124], stage0_51[125]},
      {stage0_53[42], stage0_53[43], stage0_53[44], stage0_53[45], stage0_53[46], stage0_53[47]},
      {stage1_55[7],stage1_54[13],stage1_53[26],stage1_52[37],stage1_51[46]}
   );
   gpc606_5 gpc497 (
      {stage0_51[126], stage0_51[127], 1'b0, 1'b0, 1'b0, 1'b0},
      {stage0_53[48], stage0_53[49], stage0_53[50], stage0_53[51], stage0_53[52], stage0_53[53]},
      {stage1_55[8],stage1_54[14],stage1_53[27],stage1_52[38],stage1_51[47]}
   );
   gpc606_5 gpc498 (
      {stage0_52[36], stage0_52[37], stage0_52[38], stage0_52[39], stage0_52[40], stage0_52[41]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[9],stage1_54[15],stage1_53[28],stage1_52[39]}
   );
   gpc606_5 gpc499 (
      {stage0_52[42], stage0_52[43], stage0_52[44], stage0_52[45], stage0_52[46], stage0_52[47]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[10],stage1_54[16],stage1_53[29],stage1_52[40]}
   );
   gpc606_5 gpc500 (
      {stage0_52[48], stage0_52[49], stage0_52[50], stage0_52[51], stage0_52[52], stage0_52[53]},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[11],stage1_54[17],stage1_53[30],stage1_52[41]}
   );
   gpc606_5 gpc501 (
      {stage0_52[54], stage0_52[55], stage0_52[56], stage0_52[57], stage0_52[58], stage0_52[59]},
      {stage0_54[18], stage0_54[19], stage0_54[20], stage0_54[21], stage0_54[22], stage0_54[23]},
      {stage1_56[3],stage1_55[12],stage1_54[18],stage1_53[31],stage1_52[42]}
   );
   gpc606_5 gpc502 (
      {stage0_52[60], stage0_52[61], stage0_52[62], stage0_52[63], stage0_52[64], stage0_52[65]},
      {stage0_54[24], stage0_54[25], stage0_54[26], stage0_54[27], stage0_54[28], stage0_54[29]},
      {stage1_56[4],stage1_55[13],stage1_54[19],stage1_53[32],stage1_52[43]}
   );
   gpc606_5 gpc503 (
      {stage0_52[66], stage0_52[67], stage0_52[68], stage0_52[69], stage0_52[70], stage0_52[71]},
      {stage0_54[30], stage0_54[31], stage0_54[32], stage0_54[33], stage0_54[34], stage0_54[35]},
      {stage1_56[5],stage1_55[14],stage1_54[20],stage1_53[33],stage1_52[44]}
   );
   gpc606_5 gpc504 (
      {stage0_52[72], stage0_52[73], stage0_52[74], stage0_52[75], stage0_52[76], stage0_52[77]},
      {stage0_54[36], stage0_54[37], stage0_54[38], stage0_54[39], stage0_54[40], stage0_54[41]},
      {stage1_56[6],stage1_55[15],stage1_54[21],stage1_53[34],stage1_52[45]}
   );
   gpc606_5 gpc505 (
      {stage0_52[78], stage0_52[79], stage0_52[80], stage0_52[81], stage0_52[82], stage0_52[83]},
      {stage0_54[42], stage0_54[43], stage0_54[44], stage0_54[45], stage0_54[46], stage0_54[47]},
      {stage1_56[7],stage1_55[16],stage1_54[22],stage1_53[35],stage1_52[46]}
   );
   gpc606_5 gpc506 (
      {stage0_52[84], stage0_52[85], stage0_52[86], stage0_52[87], stage0_52[88], stage0_52[89]},
      {stage0_54[48], stage0_54[49], stage0_54[50], stage0_54[51], stage0_54[52], stage0_54[53]},
      {stage1_56[8],stage1_55[17],stage1_54[23],stage1_53[36],stage1_52[47]}
   );
   gpc606_5 gpc507 (
      {stage0_52[90], stage0_52[91], stage0_52[92], stage0_52[93], stage0_52[94], stage0_52[95]},
      {stage0_54[54], stage0_54[55], stage0_54[56], stage0_54[57], stage0_54[58], stage0_54[59]},
      {stage1_56[9],stage1_55[18],stage1_54[24],stage1_53[37],stage1_52[48]}
   );
   gpc606_5 gpc508 (
      {stage0_52[96], stage0_52[97], stage0_52[98], stage0_52[99], stage0_52[100], stage0_52[101]},
      {stage0_54[60], stage0_54[61], stage0_54[62], stage0_54[63], stage0_54[64], stage0_54[65]},
      {stage1_56[10],stage1_55[19],stage1_54[25],stage1_53[38],stage1_52[49]}
   );
   gpc606_5 gpc509 (
      {stage0_52[102], stage0_52[103], stage0_52[104], stage0_52[105], stage0_52[106], stage0_52[107]},
      {stage0_54[66], stage0_54[67], stage0_54[68], stage0_54[69], stage0_54[70], stage0_54[71]},
      {stage1_56[11],stage1_55[20],stage1_54[26],stage1_53[39],stage1_52[50]}
   );
   gpc606_5 gpc510 (
      {stage0_52[108], stage0_52[109], stage0_52[110], stage0_52[111], stage0_52[112], stage0_52[113]},
      {stage0_54[72], stage0_54[73], stage0_54[74], stage0_54[75], stage0_54[76], stage0_54[77]},
      {stage1_56[12],stage1_55[21],stage1_54[27],stage1_53[40],stage1_52[51]}
   );
   gpc606_5 gpc511 (
      {stage0_52[114], stage0_52[115], stage0_52[116], stage0_52[117], stage0_52[118], stage0_52[119]},
      {stage0_54[78], stage0_54[79], stage0_54[80], stage0_54[81], stage0_54[82], stage0_54[83]},
      {stage1_56[13],stage1_55[22],stage1_54[28],stage1_53[41],stage1_52[52]}
   );
   gpc1343_5 gpc512 (
      {stage0_53[54], stage0_53[55], stage0_53[56]},
      {stage0_54[84], stage0_54[85], stage0_54[86], stage0_54[87]},
      {stage0_55[0], stage0_55[1], stage0_55[2]},
      {stage0_56[0]},
      {stage1_57[0],stage1_56[14],stage1_55[23],stage1_54[29],stage1_53[42]}
   );
   gpc606_5 gpc513 (
      {stage0_53[57], stage0_53[58], stage0_53[59], stage0_53[60], stage0_53[61], stage0_53[62]},
      {stage0_55[3], stage0_55[4], stage0_55[5], stage0_55[6], stage0_55[7], stage0_55[8]},
      {stage1_57[1],stage1_56[15],stage1_55[24],stage1_54[30],stage1_53[43]}
   );
   gpc606_5 gpc514 (
      {stage0_53[63], stage0_53[64], stage0_53[65], stage0_53[66], stage0_53[67], stage0_53[68]},
      {stage0_55[9], stage0_55[10], stage0_55[11], stage0_55[12], stage0_55[13], stage0_55[14]},
      {stage1_57[2],stage1_56[16],stage1_55[25],stage1_54[31],stage1_53[44]}
   );
   gpc606_5 gpc515 (
      {stage0_53[69], stage0_53[70], stage0_53[71], stage0_53[72], stage0_53[73], stage0_53[74]},
      {stage0_55[15], stage0_55[16], stage0_55[17], stage0_55[18], stage0_55[19], stage0_55[20]},
      {stage1_57[3],stage1_56[17],stage1_55[26],stage1_54[32],stage1_53[45]}
   );
   gpc606_5 gpc516 (
      {stage0_53[75], stage0_53[76], stage0_53[77], stage0_53[78], stage0_53[79], stage0_53[80]},
      {stage0_55[21], stage0_55[22], stage0_55[23], stage0_55[24], stage0_55[25], stage0_55[26]},
      {stage1_57[4],stage1_56[18],stage1_55[27],stage1_54[33],stage1_53[46]}
   );
   gpc606_5 gpc517 (
      {stage0_53[81], stage0_53[82], stage0_53[83], stage0_53[84], stage0_53[85], stage0_53[86]},
      {stage0_55[27], stage0_55[28], stage0_55[29], stage0_55[30], stage0_55[31], stage0_55[32]},
      {stage1_57[5],stage1_56[19],stage1_55[28],stage1_54[34],stage1_53[47]}
   );
   gpc606_5 gpc518 (
      {stage0_53[87], stage0_53[88], stage0_53[89], stage0_53[90], stage0_53[91], stage0_53[92]},
      {stage0_55[33], stage0_55[34], stage0_55[35], stage0_55[36], stage0_55[37], stage0_55[38]},
      {stage1_57[6],stage1_56[20],stage1_55[29],stage1_54[35],stage1_53[48]}
   );
   gpc606_5 gpc519 (
      {stage0_53[93], stage0_53[94], stage0_53[95], stage0_53[96], stage0_53[97], stage0_53[98]},
      {stage0_55[39], stage0_55[40], stage0_55[41], stage0_55[42], stage0_55[43], stage0_55[44]},
      {stage1_57[7],stage1_56[21],stage1_55[30],stage1_54[36],stage1_53[49]}
   );
   gpc606_5 gpc520 (
      {stage0_53[99], stage0_53[100], stage0_53[101], stage0_53[102], stage0_53[103], stage0_53[104]},
      {stage0_55[45], stage0_55[46], stage0_55[47], stage0_55[48], stage0_55[49], stage0_55[50]},
      {stage1_57[8],stage1_56[22],stage1_55[31],stage1_54[37],stage1_53[50]}
   );
   gpc615_5 gpc521 (
      {stage0_53[105], stage0_53[106], stage0_53[107], stage0_53[108], stage0_53[109]},
      {stage0_54[88]},
      {stage0_55[51], stage0_55[52], stage0_55[53], stage0_55[54], stage0_55[55], stage0_55[56]},
      {stage1_57[9],stage1_56[23],stage1_55[32],stage1_54[38],stage1_53[51]}
   );
   gpc615_5 gpc522 (
      {stage0_53[110], stage0_53[111], stage0_53[112], stage0_53[113], stage0_53[114]},
      {stage0_54[89]},
      {stage0_55[57], stage0_55[58], stage0_55[59], stage0_55[60], stage0_55[61], stage0_55[62]},
      {stage1_57[10],stage1_56[24],stage1_55[33],stage1_54[39],stage1_53[52]}
   );
   gpc615_5 gpc523 (
      {stage0_53[115], stage0_53[116], stage0_53[117], stage0_53[118], stage0_53[119]},
      {stage0_54[90]},
      {stage0_55[63], stage0_55[64], stage0_55[65], stage0_55[66], stage0_55[67], stage0_55[68]},
      {stage1_57[11],stage1_56[25],stage1_55[34],stage1_54[40],stage1_53[53]}
   );
   gpc606_5 gpc524 (
      {stage0_54[91], stage0_54[92], stage0_54[93], stage0_54[94], stage0_54[95], stage0_54[96]},
      {stage0_56[1], stage0_56[2], stage0_56[3], stage0_56[4], stage0_56[5], stage0_56[6]},
      {stage1_58[0],stage1_57[12],stage1_56[26],stage1_55[35],stage1_54[41]}
   );
   gpc606_5 gpc525 (
      {stage0_54[97], stage0_54[98], stage0_54[99], stage0_54[100], stage0_54[101], stage0_54[102]},
      {stage0_56[7], stage0_56[8], stage0_56[9], stage0_56[10], stage0_56[11], stage0_56[12]},
      {stage1_58[1],stage1_57[13],stage1_56[27],stage1_55[36],stage1_54[42]}
   );
   gpc615_5 gpc526 (
      {stage0_54[103], stage0_54[104], stage0_54[105], stage0_54[106], stage0_54[107]},
      {stage0_55[69]},
      {stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17], stage0_56[18]},
      {stage1_58[2],stage1_57[14],stage1_56[28],stage1_55[37],stage1_54[43]}
   );
   gpc615_5 gpc527 (
      {stage0_54[108], stage0_54[109], stage0_54[110], stage0_54[111], stage0_54[112]},
      {stage0_55[70]},
      {stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22], stage0_56[23], stage0_56[24]},
      {stage1_58[3],stage1_57[15],stage1_56[29],stage1_55[38],stage1_54[44]}
   );
   gpc615_5 gpc528 (
      {stage0_54[113], stage0_54[114], stage0_54[115], stage0_54[116], stage0_54[117]},
      {stage0_55[71]},
      {stage0_56[25], stage0_56[26], stage0_56[27], stage0_56[28], stage0_56[29], stage0_56[30]},
      {stage1_58[4],stage1_57[16],stage1_56[30],stage1_55[39],stage1_54[45]}
   );
   gpc615_5 gpc529 (
      {stage0_54[118], stage0_54[119], stage0_54[120], stage0_54[121], stage0_54[122]},
      {stage0_55[72]},
      {stage0_56[31], stage0_56[32], stage0_56[33], stage0_56[34], stage0_56[35], stage0_56[36]},
      {stage1_58[5],stage1_57[17],stage1_56[31],stage1_55[40],stage1_54[46]}
   );
   gpc1163_5 gpc530 (
      {stage0_55[73], stage0_55[74], stage0_55[75]},
      {stage0_56[37], stage0_56[38], stage0_56[39], stage0_56[40], stage0_56[41], stage0_56[42]},
      {stage0_57[0]},
      {stage0_58[0]},
      {stage1_59[0],stage1_58[6],stage1_57[18],stage1_56[32],stage1_55[41]}
   );
   gpc1163_5 gpc531 (
      {stage0_55[76], stage0_55[77], stage0_55[78]},
      {stage0_56[43], stage0_56[44], stage0_56[45], stage0_56[46], stage0_56[47], stage0_56[48]},
      {stage0_57[1]},
      {stage0_58[1]},
      {stage1_59[1],stage1_58[7],stage1_57[19],stage1_56[33],stage1_55[42]}
   );
   gpc606_5 gpc532 (
      {stage0_55[79], stage0_55[80], stage0_55[81], stage0_55[82], stage0_55[83], stage0_55[84]},
      {stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5], stage0_57[6], stage0_57[7]},
      {stage1_59[2],stage1_58[8],stage1_57[20],stage1_56[34],stage1_55[43]}
   );
   gpc606_5 gpc533 (
      {stage0_55[85], stage0_55[86], stage0_55[87], stage0_55[88], stage0_55[89], stage0_55[90]},
      {stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11], stage0_57[12], stage0_57[13]},
      {stage1_59[3],stage1_58[9],stage1_57[21],stage1_56[35],stage1_55[44]}
   );
   gpc606_5 gpc534 (
      {stage0_55[91], stage0_55[92], stage0_55[93], stage0_55[94], stage0_55[95], stage0_55[96]},
      {stage0_57[14], stage0_57[15], stage0_57[16], stage0_57[17], stage0_57[18], stage0_57[19]},
      {stage1_59[4],stage1_58[10],stage1_57[22],stage1_56[36],stage1_55[45]}
   );
   gpc606_5 gpc535 (
      {stage0_55[97], stage0_55[98], stage0_55[99], stage0_55[100], stage0_55[101], stage0_55[102]},
      {stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23], stage0_57[24], stage0_57[25]},
      {stage1_59[5],stage1_58[11],stage1_57[23],stage1_56[37],stage1_55[46]}
   );
   gpc615_5 gpc536 (
      {stage0_55[103], stage0_55[104], stage0_55[105], stage0_55[106], stage0_55[107]},
      {stage0_56[49]},
      {stage0_57[26], stage0_57[27], stage0_57[28], stage0_57[29], stage0_57[30], stage0_57[31]},
      {stage1_59[6],stage1_58[12],stage1_57[24],stage1_56[38],stage1_55[47]}
   );
   gpc606_5 gpc537 (
      {stage0_56[50], stage0_56[51], stage0_56[52], stage0_56[53], stage0_56[54], stage0_56[55]},
      {stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5], stage0_58[6], stage0_58[7]},
      {stage1_60[0],stage1_59[7],stage1_58[13],stage1_57[25],stage1_56[39]}
   );
   gpc606_5 gpc538 (
      {stage0_56[56], stage0_56[57], stage0_56[58], stage0_56[59], stage0_56[60], stage0_56[61]},
      {stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11], stage0_58[12], stage0_58[13]},
      {stage1_60[1],stage1_59[8],stage1_58[14],stage1_57[26],stage1_56[40]}
   );
   gpc606_5 gpc539 (
      {stage0_56[62], stage0_56[63], stage0_56[64], stage0_56[65], stage0_56[66], stage0_56[67]},
      {stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17], stage0_58[18], stage0_58[19]},
      {stage1_60[2],stage1_59[9],stage1_58[15],stage1_57[27],stage1_56[41]}
   );
   gpc606_5 gpc540 (
      {stage0_56[68], stage0_56[69], stage0_56[70], stage0_56[71], stage0_56[72], stage0_56[73]},
      {stage0_58[20], stage0_58[21], stage0_58[22], stage0_58[23], stage0_58[24], stage0_58[25]},
      {stage1_60[3],stage1_59[10],stage1_58[16],stage1_57[28],stage1_56[42]}
   );
   gpc606_5 gpc541 (
      {stage0_56[74], stage0_56[75], stage0_56[76], stage0_56[77], stage0_56[78], stage0_56[79]},
      {stage0_58[26], stage0_58[27], stage0_58[28], stage0_58[29], stage0_58[30], stage0_58[31]},
      {stage1_60[4],stage1_59[11],stage1_58[17],stage1_57[29],stage1_56[43]}
   );
   gpc606_5 gpc542 (
      {stage0_56[80], stage0_56[81], stage0_56[82], stage0_56[83], stage0_56[84], stage0_56[85]},
      {stage0_58[32], stage0_58[33], stage0_58[34], stage0_58[35], stage0_58[36], stage0_58[37]},
      {stage1_60[5],stage1_59[12],stage1_58[18],stage1_57[30],stage1_56[44]}
   );
   gpc606_5 gpc543 (
      {stage0_56[86], stage0_56[87], stage0_56[88], stage0_56[89], stage0_56[90], stage0_56[91]},
      {stage0_58[38], stage0_58[39], stage0_58[40], stage0_58[41], stage0_58[42], stage0_58[43]},
      {stage1_60[6],stage1_59[13],stage1_58[19],stage1_57[31],stage1_56[45]}
   );
   gpc606_5 gpc544 (
      {stage0_56[92], stage0_56[93], stage0_56[94], stage0_56[95], stage0_56[96], stage0_56[97]},
      {stage0_58[44], stage0_58[45], stage0_58[46], stage0_58[47], stage0_58[48], stage0_58[49]},
      {stage1_60[7],stage1_59[14],stage1_58[20],stage1_57[32],stage1_56[46]}
   );
   gpc606_5 gpc545 (
      {stage0_56[98], stage0_56[99], stage0_56[100], stage0_56[101], stage0_56[102], stage0_56[103]},
      {stage0_58[50], stage0_58[51], stage0_58[52], stage0_58[53], stage0_58[54], stage0_58[55]},
      {stage1_60[8],stage1_59[15],stage1_58[21],stage1_57[33],stage1_56[47]}
   );
   gpc606_5 gpc546 (
      {stage0_56[104], stage0_56[105], stage0_56[106], stage0_56[107], stage0_56[108], stage0_56[109]},
      {stage0_58[56], stage0_58[57], stage0_58[58], stage0_58[59], stage0_58[60], stage0_58[61]},
      {stage1_60[9],stage1_59[16],stage1_58[22],stage1_57[34],stage1_56[48]}
   );
   gpc606_5 gpc547 (
      {stage0_56[110], stage0_56[111], stage0_56[112], stage0_56[113], stage0_56[114], stage0_56[115]},
      {stage0_58[62], stage0_58[63], stage0_58[64], stage0_58[65], stage0_58[66], stage0_58[67]},
      {stage1_60[10],stage1_59[17],stage1_58[23],stage1_57[35],stage1_56[49]}
   );
   gpc606_5 gpc548 (
      {stage0_56[116], stage0_56[117], stage0_56[118], stage0_56[119], stage0_56[120], stage0_56[121]},
      {stage0_58[68], stage0_58[69], stage0_58[70], stage0_58[71], stage0_58[72], stage0_58[73]},
      {stage1_60[11],stage1_59[18],stage1_58[24],stage1_57[36],stage1_56[50]}
   );
   gpc606_5 gpc549 (
      {stage0_57[32], stage0_57[33], stage0_57[34], stage0_57[35], stage0_57[36], stage0_57[37]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[12],stage1_59[19],stage1_58[25],stage1_57[37]}
   );
   gpc606_5 gpc550 (
      {stage0_57[38], stage0_57[39], stage0_57[40], stage0_57[41], stage0_57[42], stage0_57[43]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[13],stage1_59[20],stage1_58[26],stage1_57[38]}
   );
   gpc606_5 gpc551 (
      {stage0_57[44], stage0_57[45], stage0_57[46], stage0_57[47], stage0_57[48], stage0_57[49]},
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage1_61[2],stage1_60[14],stage1_59[21],stage1_58[27],stage1_57[39]}
   );
   gpc606_5 gpc552 (
      {stage0_57[50], stage0_57[51], stage0_57[52], stage0_57[53], stage0_57[54], stage0_57[55]},
      {stage0_59[18], stage0_59[19], stage0_59[20], stage0_59[21], stage0_59[22], stage0_59[23]},
      {stage1_61[3],stage1_60[15],stage1_59[22],stage1_58[28],stage1_57[40]}
   );
   gpc606_5 gpc553 (
      {stage0_57[56], stage0_57[57], stage0_57[58], stage0_57[59], stage0_57[60], stage0_57[61]},
      {stage0_59[24], stage0_59[25], stage0_59[26], stage0_59[27], stage0_59[28], stage0_59[29]},
      {stage1_61[4],stage1_60[16],stage1_59[23],stage1_58[29],stage1_57[41]}
   );
   gpc606_5 gpc554 (
      {stage0_57[62], stage0_57[63], stage0_57[64], stage0_57[65], stage0_57[66], stage0_57[67]},
      {stage0_59[30], stage0_59[31], stage0_59[32], stage0_59[33], stage0_59[34], stage0_59[35]},
      {stage1_61[5],stage1_60[17],stage1_59[24],stage1_58[30],stage1_57[42]}
   );
   gpc606_5 gpc555 (
      {stage0_57[68], stage0_57[69], stage0_57[70], stage0_57[71], stage0_57[72], stage0_57[73]},
      {stage0_59[36], stage0_59[37], stage0_59[38], stage0_59[39], stage0_59[40], stage0_59[41]},
      {stage1_61[6],stage1_60[18],stage1_59[25],stage1_58[31],stage1_57[43]}
   );
   gpc606_5 gpc556 (
      {stage0_57[74], stage0_57[75], stage0_57[76], stage0_57[77], stage0_57[78], stage0_57[79]},
      {stage0_59[42], stage0_59[43], stage0_59[44], stage0_59[45], stage0_59[46], stage0_59[47]},
      {stage1_61[7],stage1_60[19],stage1_59[26],stage1_58[32],stage1_57[44]}
   );
   gpc606_5 gpc557 (
      {stage0_57[80], stage0_57[81], stage0_57[82], stage0_57[83], stage0_57[84], stage0_57[85]},
      {stage0_59[48], stage0_59[49], stage0_59[50], stage0_59[51], stage0_59[52], stage0_59[53]},
      {stage1_61[8],stage1_60[20],stage1_59[27],stage1_58[33],stage1_57[45]}
   );
   gpc606_5 gpc558 (
      {stage0_57[86], stage0_57[87], stage0_57[88], stage0_57[89], stage0_57[90], stage0_57[91]},
      {stage0_59[54], stage0_59[55], stage0_59[56], stage0_59[57], stage0_59[58], stage0_59[59]},
      {stage1_61[9],stage1_60[21],stage1_59[28],stage1_58[34],stage1_57[46]}
   );
   gpc606_5 gpc559 (
      {stage0_57[92], stage0_57[93], stage0_57[94], stage0_57[95], stage0_57[96], stage0_57[97]},
      {stage0_59[60], stage0_59[61], stage0_59[62], stage0_59[63], stage0_59[64], stage0_59[65]},
      {stage1_61[10],stage1_60[22],stage1_59[29],stage1_58[35],stage1_57[47]}
   );
   gpc606_5 gpc560 (
      {stage0_57[98], stage0_57[99], stage0_57[100], stage0_57[101], stage0_57[102], stage0_57[103]},
      {stage0_59[66], stage0_59[67], stage0_59[68], stage0_59[69], stage0_59[70], stage0_59[71]},
      {stage1_61[11],stage1_60[23],stage1_59[30],stage1_58[36],stage1_57[48]}
   );
   gpc606_5 gpc561 (
      {stage0_57[104], stage0_57[105], stage0_57[106], stage0_57[107], stage0_57[108], stage0_57[109]},
      {stage0_59[72], stage0_59[73], stage0_59[74], stage0_59[75], stage0_59[76], stage0_59[77]},
      {stage1_61[12],stage1_60[24],stage1_59[31],stage1_58[37],stage1_57[49]}
   );
   gpc606_5 gpc562 (
      {stage0_57[110], stage0_57[111], stage0_57[112], stage0_57[113], stage0_57[114], stage0_57[115]},
      {stage0_59[78], stage0_59[79], stage0_59[80], stage0_59[81], stage0_59[82], stage0_59[83]},
      {stage1_61[13],stage1_60[25],stage1_59[32],stage1_58[38],stage1_57[50]}
   );
   gpc606_5 gpc563 (
      {stage0_57[116], stage0_57[117], stage0_57[118], stage0_57[119], stage0_57[120], stage0_57[121]},
      {stage0_59[84], stage0_59[85], stage0_59[86], stage0_59[87], stage0_59[88], stage0_59[89]},
      {stage1_61[14],stage1_60[26],stage1_59[33],stage1_58[39],stage1_57[51]}
   );
   gpc615_5 gpc564 (
      {stage0_58[74], stage0_58[75], stage0_58[76], stage0_58[77], stage0_58[78]},
      {stage0_59[90]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3], stage0_60[4], stage0_60[5]},
      {stage1_62[0],stage1_61[15],stage1_60[27],stage1_59[34],stage1_58[40]}
   );
   gpc615_5 gpc565 (
      {stage0_58[79], stage0_58[80], stage0_58[81], stage0_58[82], stage0_58[83]},
      {stage0_59[91]},
      {stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9], stage0_60[10], stage0_60[11]},
      {stage1_62[1],stage1_61[16],stage1_60[28],stage1_59[35],stage1_58[41]}
   );
   gpc615_5 gpc566 (
      {stage0_58[84], stage0_58[85], stage0_58[86], stage0_58[87], stage0_58[88]},
      {stage0_59[92]},
      {stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15], stage0_60[16], stage0_60[17]},
      {stage1_62[2],stage1_61[17],stage1_60[29],stage1_59[36],stage1_58[42]}
   );
   gpc615_5 gpc567 (
      {stage0_58[89], stage0_58[90], stage0_58[91], stage0_58[92], stage0_58[93]},
      {stage0_59[93]},
      {stage0_60[18], stage0_60[19], stage0_60[20], stage0_60[21], stage0_60[22], stage0_60[23]},
      {stage1_62[3],stage1_61[18],stage1_60[30],stage1_59[37],stage1_58[43]}
   );
   gpc615_5 gpc568 (
      {stage0_58[94], stage0_58[95], stage0_58[96], stage0_58[97], stage0_58[98]},
      {stage0_59[94]},
      {stage0_60[24], stage0_60[25], stage0_60[26], stage0_60[27], stage0_60[28], stage0_60[29]},
      {stage1_62[4],stage1_61[19],stage1_60[31],stage1_59[38],stage1_58[44]}
   );
   gpc615_5 gpc569 (
      {stage0_58[99], stage0_58[100], stage0_58[101], stage0_58[102], stage0_58[103]},
      {stage0_59[95]},
      {stage0_60[30], stage0_60[31], stage0_60[32], stage0_60[33], stage0_60[34], stage0_60[35]},
      {stage1_62[5],stage1_61[20],stage1_60[32],stage1_59[39],stage1_58[45]}
   );
   gpc615_5 gpc570 (
      {stage0_58[104], stage0_58[105], stage0_58[106], stage0_58[107], stage0_58[108]},
      {stage0_59[96]},
      {stage0_60[36], stage0_60[37], stage0_60[38], stage0_60[39], stage0_60[40], stage0_60[41]},
      {stage1_62[6],stage1_61[21],stage1_60[33],stage1_59[40],stage1_58[46]}
   );
   gpc615_5 gpc571 (
      {stage0_58[109], stage0_58[110], stage0_58[111], stage0_58[112], stage0_58[113]},
      {stage0_59[97]},
      {stage0_60[42], stage0_60[43], stage0_60[44], stage0_60[45], stage0_60[46], stage0_60[47]},
      {stage1_62[7],stage1_61[22],stage1_60[34],stage1_59[41],stage1_58[47]}
   );
   gpc623_5 gpc572 (
      {stage0_58[114], stage0_58[115], stage0_58[116]},
      {stage0_59[98], stage0_59[99]},
      {stage0_60[48], stage0_60[49], stage0_60[50], stage0_60[51], stage0_60[52], stage0_60[53]},
      {stage1_62[8],stage1_61[23],stage1_60[35],stage1_59[42],stage1_58[48]}
   );
   gpc606_5 gpc573 (
      {stage0_59[100], stage0_59[101], stage0_59[102], stage0_59[103], stage0_59[104], stage0_59[105]},
      {stage0_61[0], stage0_61[1], stage0_61[2], stage0_61[3], stage0_61[4], stage0_61[5]},
      {stage1_63[0],stage1_62[9],stage1_61[24],stage1_60[36],stage1_59[43]}
   );
   gpc606_5 gpc574 (
      {stage0_59[106], stage0_59[107], stage0_59[108], stage0_59[109], stage0_59[110], stage0_59[111]},
      {stage0_61[6], stage0_61[7], stage0_61[8], stage0_61[9], stage0_61[10], stage0_61[11]},
      {stage1_63[1],stage1_62[10],stage1_61[25],stage1_60[37],stage1_59[44]}
   );
   gpc606_5 gpc575 (
      {stage0_59[112], stage0_59[113], stage0_59[114], stage0_59[115], stage0_59[116], stage0_59[117]},
      {stage0_61[12], stage0_61[13], stage0_61[14], stage0_61[15], stage0_61[16], stage0_61[17]},
      {stage1_63[2],stage1_62[11],stage1_61[26],stage1_60[38],stage1_59[45]}
   );
   gpc606_5 gpc576 (
      {stage0_60[54], stage0_60[55], stage0_60[56], stage0_60[57], stage0_60[58], stage0_60[59]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3], stage0_62[4], stage0_62[5]},
      {stage1_64[0],stage1_63[3],stage1_62[12],stage1_61[27],stage1_60[39]}
   );
   gpc606_5 gpc577 (
      {stage0_60[60], stage0_60[61], stage0_60[62], stage0_60[63], stage0_60[64], stage0_60[65]},
      {stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9], stage0_62[10], stage0_62[11]},
      {stage1_64[1],stage1_63[4],stage1_62[13],stage1_61[28],stage1_60[40]}
   );
   gpc606_5 gpc578 (
      {stage0_60[66], stage0_60[67], stage0_60[68], stage0_60[69], stage0_60[70], stage0_60[71]},
      {stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15], stage0_62[16], stage0_62[17]},
      {stage1_64[2],stage1_63[5],stage1_62[14],stage1_61[29],stage1_60[41]}
   );
   gpc606_5 gpc579 (
      {stage0_60[72], stage0_60[73], stage0_60[74], stage0_60[75], stage0_60[76], stage0_60[77]},
      {stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21], stage0_62[22], stage0_62[23]},
      {stage1_64[3],stage1_63[6],stage1_62[15],stage1_61[30],stage1_60[42]}
   );
   gpc606_5 gpc580 (
      {stage0_60[78], stage0_60[79], stage0_60[80], stage0_60[81], stage0_60[82], stage0_60[83]},
      {stage0_62[24], stage0_62[25], stage0_62[26], stage0_62[27], stage0_62[28], stage0_62[29]},
      {stage1_64[4],stage1_63[7],stage1_62[16],stage1_61[31],stage1_60[43]}
   );
   gpc606_5 gpc581 (
      {stage0_60[84], stage0_60[85], stage0_60[86], stage0_60[87], stage0_60[88], stage0_60[89]},
      {stage0_62[30], stage0_62[31], stage0_62[32], stage0_62[33], stage0_62[34], stage0_62[35]},
      {stage1_64[5],stage1_63[8],stage1_62[17],stage1_61[32],stage1_60[44]}
   );
   gpc606_5 gpc582 (
      {stage0_60[90], stage0_60[91], stage0_60[92], stage0_60[93], stage0_60[94], stage0_60[95]},
      {stage0_62[36], stage0_62[37], stage0_62[38], stage0_62[39], stage0_62[40], stage0_62[41]},
      {stage1_64[6],stage1_63[9],stage1_62[18],stage1_61[33],stage1_60[45]}
   );
   gpc606_5 gpc583 (
      {stage0_60[96], stage0_60[97], stage0_60[98], stage0_60[99], stage0_60[100], stage0_60[101]},
      {stage0_62[42], stage0_62[43], stage0_62[44], stage0_62[45], stage0_62[46], stage0_62[47]},
      {stage1_64[7],stage1_63[10],stage1_62[19],stage1_61[34],stage1_60[46]}
   );
   gpc606_5 gpc584 (
      {stage0_60[102], stage0_60[103], stage0_60[104], stage0_60[105], stage0_60[106], stage0_60[107]},
      {stage0_62[48], stage0_62[49], stage0_62[50], stage0_62[51], stage0_62[52], stage0_62[53]},
      {stage1_64[8],stage1_63[11],stage1_62[20],stage1_61[35],stage1_60[47]}
   );
   gpc606_5 gpc585 (
      {stage0_60[108], stage0_60[109], stage0_60[110], stage0_60[111], stage0_60[112], stage0_60[113]},
      {stage0_62[54], stage0_62[55], stage0_62[56], stage0_62[57], stage0_62[58], stage0_62[59]},
      {stage1_64[9],stage1_63[12],stage1_62[21],stage1_61[36],stage1_60[48]}
   );
   gpc606_5 gpc586 (
      {stage0_60[114], stage0_60[115], stage0_60[116], stage0_60[117], stage0_60[118], stage0_60[119]},
      {stage0_62[60], stage0_62[61], stage0_62[62], stage0_62[63], stage0_62[64], stage0_62[65]},
      {stage1_64[10],stage1_63[13],stage1_62[22],stage1_61[37],stage1_60[49]}
   );
   gpc606_5 gpc587 (
      {stage0_60[120], stage0_60[121], stage0_60[122], stage0_60[123], stage0_60[124], stage0_60[125]},
      {stage0_62[66], stage0_62[67], stage0_62[68], stage0_62[69], stage0_62[70], stage0_62[71]},
      {stage1_64[11],stage1_63[14],stage1_62[23],stage1_61[38],stage1_60[50]}
   );
   gpc606_5 gpc588 (
      {stage0_61[18], stage0_61[19], stage0_61[20], stage0_61[21], stage0_61[22], stage0_61[23]},
      {stage0_63[0], stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5]},
      {stage1_65[0],stage1_64[12],stage1_63[15],stage1_62[24],stage1_61[39]}
   );
   gpc606_5 gpc589 (
      {stage0_61[24], stage0_61[25], stage0_61[26], stage0_61[27], stage0_61[28], stage0_61[29]},
      {stage0_63[6], stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11]},
      {stage1_65[1],stage1_64[13],stage1_63[16],stage1_62[25],stage1_61[40]}
   );
   gpc606_5 gpc590 (
      {stage0_61[30], stage0_61[31], stage0_61[32], stage0_61[33], stage0_61[34], stage0_61[35]},
      {stage0_63[12], stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17]},
      {stage1_65[2],stage1_64[14],stage1_63[17],stage1_62[26],stage1_61[41]}
   );
   gpc606_5 gpc591 (
      {stage0_61[36], stage0_61[37], stage0_61[38], stage0_61[39], stage0_61[40], stage0_61[41]},
      {stage0_63[18], stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23]},
      {stage1_65[3],stage1_64[15],stage1_63[18],stage1_62[27],stage1_61[42]}
   );
   gpc606_5 gpc592 (
      {stage0_61[42], stage0_61[43], stage0_61[44], stage0_61[45], stage0_61[46], stage0_61[47]},
      {stage0_63[24], stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29]},
      {stage1_65[4],stage1_64[16],stage1_63[19],stage1_62[28],stage1_61[43]}
   );
   gpc606_5 gpc593 (
      {stage0_61[48], stage0_61[49], stage0_61[50], stage0_61[51], stage0_61[52], stage0_61[53]},
      {stage0_63[30], stage0_63[31], stage0_63[32], stage0_63[33], stage0_63[34], stage0_63[35]},
      {stage1_65[5],stage1_64[17],stage1_63[20],stage1_62[29],stage1_61[44]}
   );
   gpc606_5 gpc594 (
      {stage0_61[54], stage0_61[55], stage0_61[56], stage0_61[57], stage0_61[58], stage0_61[59]},
      {stage0_63[36], stage0_63[37], stage0_63[38], stage0_63[39], stage0_63[40], stage0_63[41]},
      {stage1_65[6],stage1_64[18],stage1_63[21],stage1_62[30],stage1_61[45]}
   );
   gpc606_5 gpc595 (
      {stage0_61[60], stage0_61[61], stage0_61[62], stage0_61[63], stage0_61[64], stage0_61[65]},
      {stage0_63[42], stage0_63[43], stage0_63[44], stage0_63[45], stage0_63[46], stage0_63[47]},
      {stage1_65[7],stage1_64[19],stage1_63[22],stage1_62[31],stage1_61[46]}
   );
   gpc606_5 gpc596 (
      {stage0_61[66], stage0_61[67], stage0_61[68], stage0_61[69], stage0_61[70], stage0_61[71]},
      {stage0_63[48], stage0_63[49], stage0_63[50], stage0_63[51], stage0_63[52], stage0_63[53]},
      {stage1_65[8],stage1_64[20],stage1_63[23],stage1_62[32],stage1_61[47]}
   );
   gpc606_5 gpc597 (
      {stage0_61[72], stage0_61[73], stage0_61[74], stage0_61[75], stage0_61[76], stage0_61[77]},
      {stage0_63[54], stage0_63[55], stage0_63[56], stage0_63[57], stage0_63[58], stage0_63[59]},
      {stage1_65[9],stage1_64[21],stage1_63[24],stage1_62[33],stage1_61[48]}
   );
   gpc606_5 gpc598 (
      {stage0_61[78], stage0_61[79], stage0_61[80], stage0_61[81], stage0_61[82], stage0_61[83]},
      {stage0_63[60], stage0_63[61], stage0_63[62], stage0_63[63], stage0_63[64], stage0_63[65]},
      {stage1_65[10],stage1_64[22],stage1_63[25],stage1_62[34],stage1_61[49]}
   );
   gpc606_5 gpc599 (
      {stage0_61[84], stage0_61[85], stage0_61[86], stage0_61[87], stage0_61[88], stage0_61[89]},
      {stage0_63[66], stage0_63[67], stage0_63[68], stage0_63[69], stage0_63[70], stage0_63[71]},
      {stage1_65[11],stage1_64[23],stage1_63[26],stage1_62[35],stage1_61[50]}
   );
   gpc606_5 gpc600 (
      {stage0_61[90], stage0_61[91], stage0_61[92], stage0_61[93], stage0_61[94], stage0_61[95]},
      {stage0_63[72], stage0_63[73], stage0_63[74], stage0_63[75], stage0_63[76], stage0_63[77]},
      {stage1_65[12],stage1_64[24],stage1_63[27],stage1_62[36],stage1_61[51]}
   );
   gpc606_5 gpc601 (
      {stage0_61[96], stage0_61[97], stage0_61[98], stage0_61[99], stage0_61[100], stage0_61[101]},
      {stage0_63[78], stage0_63[79], stage0_63[80], stage0_63[81], stage0_63[82], stage0_63[83]},
      {stage1_65[13],stage1_64[25],stage1_63[28],stage1_62[37],stage1_61[52]}
   );
   gpc606_5 gpc602 (
      {stage0_61[102], stage0_61[103], stage0_61[104], stage0_61[105], stage0_61[106], stage0_61[107]},
      {stage0_63[84], stage0_63[85], stage0_63[86], stage0_63[87], stage0_63[88], stage0_63[89]},
      {stage1_65[14],stage1_64[26],stage1_63[29],stage1_62[38],stage1_61[53]}
   );
   gpc606_5 gpc603 (
      {stage0_61[108], stage0_61[109], stage0_61[110], stage0_61[111], stage0_61[112], stage0_61[113]},
      {stage0_63[90], stage0_63[91], stage0_63[92], stage0_63[93], stage0_63[94], stage0_63[95]},
      {stage1_65[15],stage1_64[27],stage1_63[30],stage1_62[39],stage1_61[54]}
   );
   gpc606_5 gpc604 (
      {stage0_61[114], stage0_61[115], stage0_61[116], stage0_61[117], stage0_61[118], stage0_61[119]},
      {stage0_63[96], stage0_63[97], stage0_63[98], stage0_63[99], stage0_63[100], stage0_63[101]},
      {stage1_65[16],stage1_64[28],stage1_63[31],stage1_62[40],stage1_61[55]}
   );
   gpc606_5 gpc605 (
      {stage0_61[120], stage0_61[121], stage0_61[122], stage0_61[123], stage0_61[124], stage0_61[125]},
      {stage0_63[102], stage0_63[103], stage0_63[104], stage0_63[105], stage0_63[106], stage0_63[107]},
      {stage1_65[17],stage1_64[29],stage1_63[32],stage1_62[41],stage1_61[56]}
   );
   gpc1_1 gpc606 (
      {stage0_2[121]},
      {stage1_2[40]}
   );
   gpc1_1 gpc607 (
      {stage0_2[122]},
      {stage1_2[41]}
   );
   gpc1_1 gpc608 (
      {stage0_2[123]},
      {stage1_2[42]}
   );
   gpc1_1 gpc609 (
      {stage0_2[124]},
      {stage1_2[43]}
   );
   gpc1_1 gpc610 (
      {stage0_2[125]},
      {stage1_2[44]}
   );
   gpc1_1 gpc611 (
      {stage0_2[126]},
      {stage1_2[45]}
   );
   gpc1_1 gpc612 (
      {stage0_2[127]},
      {stage1_2[46]}
   );
   gpc1_1 gpc613 (
      {stage0_3[117]},
      {stage1_3[56]}
   );
   gpc1_1 gpc614 (
      {stage0_3[118]},
      {stage1_3[57]}
   );
   gpc1_1 gpc615 (
      {stage0_3[119]},
      {stage1_3[58]}
   );
   gpc1_1 gpc616 (
      {stage0_3[120]},
      {stage1_3[59]}
   );
   gpc1_1 gpc617 (
      {stage0_3[121]},
      {stage1_3[60]}
   );
   gpc1_1 gpc618 (
      {stage0_3[122]},
      {stage1_3[61]}
   );
   gpc1_1 gpc619 (
      {stage0_3[123]},
      {stage1_3[62]}
   );
   gpc1_1 gpc620 (
      {stage0_3[124]},
      {stage1_3[63]}
   );
   gpc1_1 gpc621 (
      {stage0_3[125]},
      {stage1_3[64]}
   );
   gpc1_1 gpc622 (
      {stage0_3[126]},
      {stage1_3[65]}
   );
   gpc1_1 gpc623 (
      {stage0_3[127]},
      {stage1_3[66]}
   );
   gpc1_1 gpc624 (
      {stage0_5[118]},
      {stage1_5[42]}
   );
   gpc1_1 gpc625 (
      {stage0_5[119]},
      {stage1_5[43]}
   );
   gpc1_1 gpc626 (
      {stage0_5[120]},
      {stage1_5[44]}
   );
   gpc1_1 gpc627 (
      {stage0_5[121]},
      {stage1_5[45]}
   );
   gpc1_1 gpc628 (
      {stage0_5[122]},
      {stage1_5[46]}
   );
   gpc1_1 gpc629 (
      {stage0_5[123]},
      {stage1_5[47]}
   );
   gpc1_1 gpc630 (
      {stage0_5[124]},
      {stage1_5[48]}
   );
   gpc1_1 gpc631 (
      {stage0_5[125]},
      {stage1_5[49]}
   );
   gpc1_1 gpc632 (
      {stage0_5[126]},
      {stage1_5[50]}
   );
   gpc1_1 gpc633 (
      {stage0_5[127]},
      {stage1_5[51]}
   );
   gpc1_1 gpc634 (
      {stage0_6[79]},
      {stage1_6[40]}
   );
   gpc1_1 gpc635 (
      {stage0_6[80]},
      {stage1_6[41]}
   );
   gpc1_1 gpc636 (
      {stage0_6[81]},
      {stage1_6[42]}
   );
   gpc1_1 gpc637 (
      {stage0_6[82]},
      {stage1_6[43]}
   );
   gpc1_1 gpc638 (
      {stage0_6[83]},
      {stage1_6[44]}
   );
   gpc1_1 gpc639 (
      {stage0_6[84]},
      {stage1_6[45]}
   );
   gpc1_1 gpc640 (
      {stage0_6[85]},
      {stage1_6[46]}
   );
   gpc1_1 gpc641 (
      {stage0_6[86]},
      {stage1_6[47]}
   );
   gpc1_1 gpc642 (
      {stage0_6[87]},
      {stage1_6[48]}
   );
   gpc1_1 gpc643 (
      {stage0_6[88]},
      {stage1_6[49]}
   );
   gpc1_1 gpc644 (
      {stage0_6[89]},
      {stage1_6[50]}
   );
   gpc1_1 gpc645 (
      {stage0_6[90]},
      {stage1_6[51]}
   );
   gpc1_1 gpc646 (
      {stage0_6[91]},
      {stage1_6[52]}
   );
   gpc1_1 gpc647 (
      {stage0_6[92]},
      {stage1_6[53]}
   );
   gpc1_1 gpc648 (
      {stage0_6[93]},
      {stage1_6[54]}
   );
   gpc1_1 gpc649 (
      {stage0_6[94]},
      {stage1_6[55]}
   );
   gpc1_1 gpc650 (
      {stage0_6[95]},
      {stage1_6[56]}
   );
   gpc1_1 gpc651 (
      {stage0_6[96]},
      {stage1_6[57]}
   );
   gpc1_1 gpc652 (
      {stage0_6[97]},
      {stage1_6[58]}
   );
   gpc1_1 gpc653 (
      {stage0_6[98]},
      {stage1_6[59]}
   );
   gpc1_1 gpc654 (
      {stage0_6[99]},
      {stage1_6[60]}
   );
   gpc1_1 gpc655 (
      {stage0_6[100]},
      {stage1_6[61]}
   );
   gpc1_1 gpc656 (
      {stage0_6[101]},
      {stage1_6[62]}
   );
   gpc1_1 gpc657 (
      {stage0_6[102]},
      {stage1_6[63]}
   );
   gpc1_1 gpc658 (
      {stage0_6[103]},
      {stage1_6[64]}
   );
   gpc1_1 gpc659 (
      {stage0_6[104]},
      {stage1_6[65]}
   );
   gpc1_1 gpc660 (
      {stage0_6[105]},
      {stage1_6[66]}
   );
   gpc1_1 gpc661 (
      {stage0_6[106]},
      {stage1_6[67]}
   );
   gpc1_1 gpc662 (
      {stage0_6[107]},
      {stage1_6[68]}
   );
   gpc1_1 gpc663 (
      {stage0_6[108]},
      {stage1_6[69]}
   );
   gpc1_1 gpc664 (
      {stage0_6[109]},
      {stage1_6[70]}
   );
   gpc1_1 gpc665 (
      {stage0_6[110]},
      {stage1_6[71]}
   );
   gpc1_1 gpc666 (
      {stage0_6[111]},
      {stage1_6[72]}
   );
   gpc1_1 gpc667 (
      {stage0_6[112]},
      {stage1_6[73]}
   );
   gpc1_1 gpc668 (
      {stage0_6[113]},
      {stage1_6[74]}
   );
   gpc1_1 gpc669 (
      {stage0_6[114]},
      {stage1_6[75]}
   );
   gpc1_1 gpc670 (
      {stage0_6[115]},
      {stage1_6[76]}
   );
   gpc1_1 gpc671 (
      {stage0_6[116]},
      {stage1_6[77]}
   );
   gpc1_1 gpc672 (
      {stage0_6[117]},
      {stage1_6[78]}
   );
   gpc1_1 gpc673 (
      {stage0_6[118]},
      {stage1_6[79]}
   );
   gpc1_1 gpc674 (
      {stage0_6[119]},
      {stage1_6[80]}
   );
   gpc1_1 gpc675 (
      {stage0_6[120]},
      {stage1_6[81]}
   );
   gpc1_1 gpc676 (
      {stage0_6[121]},
      {stage1_6[82]}
   );
   gpc1_1 gpc677 (
      {stage0_6[122]},
      {stage1_6[83]}
   );
   gpc1_1 gpc678 (
      {stage0_6[123]},
      {stage1_6[84]}
   );
   gpc1_1 gpc679 (
      {stage0_6[124]},
      {stage1_6[85]}
   );
   gpc1_1 gpc680 (
      {stage0_6[125]},
      {stage1_6[86]}
   );
   gpc1_1 gpc681 (
      {stage0_6[126]},
      {stage1_6[87]}
   );
   gpc1_1 gpc682 (
      {stage0_6[127]},
      {stage1_6[88]}
   );
   gpc1_1 gpc683 (
      {stage0_7[103]},
      {stage1_7[46]}
   );
   gpc1_1 gpc684 (
      {stage0_7[104]},
      {stage1_7[47]}
   );
   gpc1_1 gpc685 (
      {stage0_7[105]},
      {stage1_7[48]}
   );
   gpc1_1 gpc686 (
      {stage0_7[106]},
      {stage1_7[49]}
   );
   gpc1_1 gpc687 (
      {stage0_7[107]},
      {stage1_7[50]}
   );
   gpc1_1 gpc688 (
      {stage0_7[108]},
      {stage1_7[51]}
   );
   gpc1_1 gpc689 (
      {stage0_7[109]},
      {stage1_7[52]}
   );
   gpc1_1 gpc690 (
      {stage0_7[110]},
      {stage1_7[53]}
   );
   gpc1_1 gpc691 (
      {stage0_7[111]},
      {stage1_7[54]}
   );
   gpc1_1 gpc692 (
      {stage0_7[112]},
      {stage1_7[55]}
   );
   gpc1_1 gpc693 (
      {stage0_7[113]},
      {stage1_7[56]}
   );
   gpc1_1 gpc694 (
      {stage0_7[114]},
      {stage1_7[57]}
   );
   gpc1_1 gpc695 (
      {stage0_7[115]},
      {stage1_7[58]}
   );
   gpc1_1 gpc696 (
      {stage0_7[116]},
      {stage1_7[59]}
   );
   gpc1_1 gpc697 (
      {stage0_7[117]},
      {stage1_7[60]}
   );
   gpc1_1 gpc698 (
      {stage0_7[118]},
      {stage1_7[61]}
   );
   gpc1_1 gpc699 (
      {stage0_7[119]},
      {stage1_7[62]}
   );
   gpc1_1 gpc700 (
      {stage0_7[120]},
      {stage1_7[63]}
   );
   gpc1_1 gpc701 (
      {stage0_7[121]},
      {stage1_7[64]}
   );
   gpc1_1 gpc702 (
      {stage0_7[122]},
      {stage1_7[65]}
   );
   gpc1_1 gpc703 (
      {stage0_7[123]},
      {stage1_7[66]}
   );
   gpc1_1 gpc704 (
      {stage0_7[124]},
      {stage1_7[67]}
   );
   gpc1_1 gpc705 (
      {stage0_7[125]},
      {stage1_7[68]}
   );
   gpc1_1 gpc706 (
      {stage0_7[126]},
      {stage1_7[69]}
   );
   gpc1_1 gpc707 (
      {stage0_7[127]},
      {stage1_7[70]}
   );
   gpc1_1 gpc708 (
      {stage0_8[109]},
      {stage1_8[47]}
   );
   gpc1_1 gpc709 (
      {stage0_8[110]},
      {stage1_8[48]}
   );
   gpc1_1 gpc710 (
      {stage0_8[111]},
      {stage1_8[49]}
   );
   gpc1_1 gpc711 (
      {stage0_8[112]},
      {stage1_8[50]}
   );
   gpc1_1 gpc712 (
      {stage0_8[113]},
      {stage1_8[51]}
   );
   gpc1_1 gpc713 (
      {stage0_8[114]},
      {stage1_8[52]}
   );
   gpc1_1 gpc714 (
      {stage0_8[115]},
      {stage1_8[53]}
   );
   gpc1_1 gpc715 (
      {stage0_8[116]},
      {stage1_8[54]}
   );
   gpc1_1 gpc716 (
      {stage0_8[117]},
      {stage1_8[55]}
   );
   gpc1_1 gpc717 (
      {stage0_8[118]},
      {stage1_8[56]}
   );
   gpc1_1 gpc718 (
      {stage0_8[119]},
      {stage1_8[57]}
   );
   gpc1_1 gpc719 (
      {stage0_8[120]},
      {stage1_8[58]}
   );
   gpc1_1 gpc720 (
      {stage0_8[121]},
      {stage1_8[59]}
   );
   gpc1_1 gpc721 (
      {stage0_8[122]},
      {stage1_8[60]}
   );
   gpc1_1 gpc722 (
      {stage0_8[123]},
      {stage1_8[61]}
   );
   gpc1_1 gpc723 (
      {stage0_8[124]},
      {stage1_8[62]}
   );
   gpc1_1 gpc724 (
      {stage0_8[125]},
      {stage1_8[63]}
   );
   gpc1_1 gpc725 (
      {stage0_8[126]},
      {stage1_8[64]}
   );
   gpc1_1 gpc726 (
      {stage0_8[127]},
      {stage1_8[65]}
   );
   gpc1_1 gpc727 (
      {stage0_9[108]},
      {stage1_9[41]}
   );
   gpc1_1 gpc728 (
      {stage0_9[109]},
      {stage1_9[42]}
   );
   gpc1_1 gpc729 (
      {stage0_9[110]},
      {stage1_9[43]}
   );
   gpc1_1 gpc730 (
      {stage0_9[111]},
      {stage1_9[44]}
   );
   gpc1_1 gpc731 (
      {stage0_9[112]},
      {stage1_9[45]}
   );
   gpc1_1 gpc732 (
      {stage0_9[113]},
      {stage1_9[46]}
   );
   gpc1_1 gpc733 (
      {stage0_9[114]},
      {stage1_9[47]}
   );
   gpc1_1 gpc734 (
      {stage0_9[115]},
      {stage1_9[48]}
   );
   gpc1_1 gpc735 (
      {stage0_9[116]},
      {stage1_9[49]}
   );
   gpc1_1 gpc736 (
      {stage0_9[117]},
      {stage1_9[50]}
   );
   gpc1_1 gpc737 (
      {stage0_9[118]},
      {stage1_9[51]}
   );
   gpc1_1 gpc738 (
      {stage0_9[119]},
      {stage1_9[52]}
   );
   gpc1_1 gpc739 (
      {stage0_9[120]},
      {stage1_9[53]}
   );
   gpc1_1 gpc740 (
      {stage0_9[121]},
      {stage1_9[54]}
   );
   gpc1_1 gpc741 (
      {stage0_9[122]},
      {stage1_9[55]}
   );
   gpc1_1 gpc742 (
      {stage0_9[123]},
      {stage1_9[56]}
   );
   gpc1_1 gpc743 (
      {stage0_9[124]},
      {stage1_9[57]}
   );
   gpc1_1 gpc744 (
      {stage0_9[125]},
      {stage1_9[58]}
   );
   gpc1_1 gpc745 (
      {stage0_9[126]},
      {stage1_9[59]}
   );
   gpc1_1 gpc746 (
      {stage0_9[127]},
      {stage1_9[60]}
   );
   gpc1_1 gpc747 (
      {stage0_11[118]},
      {stage1_11[54]}
   );
   gpc1_1 gpc748 (
      {stage0_11[119]},
      {stage1_11[55]}
   );
   gpc1_1 gpc749 (
      {stage0_11[120]},
      {stage1_11[56]}
   );
   gpc1_1 gpc750 (
      {stage0_11[121]},
      {stage1_11[57]}
   );
   gpc1_1 gpc751 (
      {stage0_11[122]},
      {stage1_11[58]}
   );
   gpc1_1 gpc752 (
      {stage0_11[123]},
      {stage1_11[59]}
   );
   gpc1_1 gpc753 (
      {stage0_11[124]},
      {stage1_11[60]}
   );
   gpc1_1 gpc754 (
      {stage0_11[125]},
      {stage1_11[61]}
   );
   gpc1_1 gpc755 (
      {stage0_11[126]},
      {stage1_11[62]}
   );
   gpc1_1 gpc756 (
      {stage0_11[127]},
      {stage1_11[63]}
   );
   gpc1_1 gpc757 (
      {stage0_13[124]},
      {stage1_13[50]}
   );
   gpc1_1 gpc758 (
      {stage0_13[125]},
      {stage1_13[51]}
   );
   gpc1_1 gpc759 (
      {stage0_13[126]},
      {stage1_13[52]}
   );
   gpc1_1 gpc760 (
      {stage0_13[127]},
      {stage1_13[53]}
   );
   gpc1_1 gpc761 (
      {stage0_14[109]},
      {stage1_14[47]}
   );
   gpc1_1 gpc762 (
      {stage0_14[110]},
      {stage1_14[48]}
   );
   gpc1_1 gpc763 (
      {stage0_14[111]},
      {stage1_14[49]}
   );
   gpc1_1 gpc764 (
      {stage0_14[112]},
      {stage1_14[50]}
   );
   gpc1_1 gpc765 (
      {stage0_14[113]},
      {stage1_14[51]}
   );
   gpc1_1 gpc766 (
      {stage0_14[114]},
      {stage1_14[52]}
   );
   gpc1_1 gpc767 (
      {stage0_14[115]},
      {stage1_14[53]}
   );
   gpc1_1 gpc768 (
      {stage0_14[116]},
      {stage1_14[54]}
   );
   gpc1_1 gpc769 (
      {stage0_14[117]},
      {stage1_14[55]}
   );
   gpc1_1 gpc770 (
      {stage0_14[118]},
      {stage1_14[56]}
   );
   gpc1_1 gpc771 (
      {stage0_14[119]},
      {stage1_14[57]}
   );
   gpc1_1 gpc772 (
      {stage0_14[120]},
      {stage1_14[58]}
   );
   gpc1_1 gpc773 (
      {stage0_14[121]},
      {stage1_14[59]}
   );
   gpc1_1 gpc774 (
      {stage0_14[122]},
      {stage1_14[60]}
   );
   gpc1_1 gpc775 (
      {stage0_14[123]},
      {stage1_14[61]}
   );
   gpc1_1 gpc776 (
      {stage0_14[124]},
      {stage1_14[62]}
   );
   gpc1_1 gpc777 (
      {stage0_14[125]},
      {stage1_14[63]}
   );
   gpc1_1 gpc778 (
      {stage0_14[126]},
      {stage1_14[64]}
   );
   gpc1_1 gpc779 (
      {stage0_14[127]},
      {stage1_14[65]}
   );
   gpc1_1 gpc780 (
      {stage0_15[106]},
      {stage1_15[46]}
   );
   gpc1_1 gpc781 (
      {stage0_15[107]},
      {stage1_15[47]}
   );
   gpc1_1 gpc782 (
      {stage0_15[108]},
      {stage1_15[48]}
   );
   gpc1_1 gpc783 (
      {stage0_15[109]},
      {stage1_15[49]}
   );
   gpc1_1 gpc784 (
      {stage0_15[110]},
      {stage1_15[50]}
   );
   gpc1_1 gpc785 (
      {stage0_15[111]},
      {stage1_15[51]}
   );
   gpc1_1 gpc786 (
      {stage0_15[112]},
      {stage1_15[52]}
   );
   gpc1_1 gpc787 (
      {stage0_15[113]},
      {stage1_15[53]}
   );
   gpc1_1 gpc788 (
      {stage0_15[114]},
      {stage1_15[54]}
   );
   gpc1_1 gpc789 (
      {stage0_15[115]},
      {stage1_15[55]}
   );
   gpc1_1 gpc790 (
      {stage0_15[116]},
      {stage1_15[56]}
   );
   gpc1_1 gpc791 (
      {stage0_15[117]},
      {stage1_15[57]}
   );
   gpc1_1 gpc792 (
      {stage0_15[118]},
      {stage1_15[58]}
   );
   gpc1_1 gpc793 (
      {stage0_15[119]},
      {stage1_15[59]}
   );
   gpc1_1 gpc794 (
      {stage0_15[120]},
      {stage1_15[60]}
   );
   gpc1_1 gpc795 (
      {stage0_15[121]},
      {stage1_15[61]}
   );
   gpc1_1 gpc796 (
      {stage0_15[122]},
      {stage1_15[62]}
   );
   gpc1_1 gpc797 (
      {stage0_15[123]},
      {stage1_15[63]}
   );
   gpc1_1 gpc798 (
      {stage0_15[124]},
      {stage1_15[64]}
   );
   gpc1_1 gpc799 (
      {stage0_15[125]},
      {stage1_15[65]}
   );
   gpc1_1 gpc800 (
      {stage0_15[126]},
      {stage1_15[66]}
   );
   gpc1_1 gpc801 (
      {stage0_15[127]},
      {stage1_15[67]}
   );
   gpc1_1 gpc802 (
      {stage0_16[85]},
      {stage1_16[46]}
   );
   gpc1_1 gpc803 (
      {stage0_16[86]},
      {stage1_16[47]}
   );
   gpc1_1 gpc804 (
      {stage0_16[87]},
      {stage1_16[48]}
   );
   gpc1_1 gpc805 (
      {stage0_16[88]},
      {stage1_16[49]}
   );
   gpc1_1 gpc806 (
      {stage0_16[89]},
      {stage1_16[50]}
   );
   gpc1_1 gpc807 (
      {stage0_16[90]},
      {stage1_16[51]}
   );
   gpc1_1 gpc808 (
      {stage0_16[91]},
      {stage1_16[52]}
   );
   gpc1_1 gpc809 (
      {stage0_16[92]},
      {stage1_16[53]}
   );
   gpc1_1 gpc810 (
      {stage0_16[93]},
      {stage1_16[54]}
   );
   gpc1_1 gpc811 (
      {stage0_16[94]},
      {stage1_16[55]}
   );
   gpc1_1 gpc812 (
      {stage0_16[95]},
      {stage1_16[56]}
   );
   gpc1_1 gpc813 (
      {stage0_16[96]},
      {stage1_16[57]}
   );
   gpc1_1 gpc814 (
      {stage0_16[97]},
      {stage1_16[58]}
   );
   gpc1_1 gpc815 (
      {stage0_16[98]},
      {stage1_16[59]}
   );
   gpc1_1 gpc816 (
      {stage0_16[99]},
      {stage1_16[60]}
   );
   gpc1_1 gpc817 (
      {stage0_16[100]},
      {stage1_16[61]}
   );
   gpc1_1 gpc818 (
      {stage0_16[101]},
      {stage1_16[62]}
   );
   gpc1_1 gpc819 (
      {stage0_16[102]},
      {stage1_16[63]}
   );
   gpc1_1 gpc820 (
      {stage0_16[103]},
      {stage1_16[64]}
   );
   gpc1_1 gpc821 (
      {stage0_16[104]},
      {stage1_16[65]}
   );
   gpc1_1 gpc822 (
      {stage0_16[105]},
      {stage1_16[66]}
   );
   gpc1_1 gpc823 (
      {stage0_16[106]},
      {stage1_16[67]}
   );
   gpc1_1 gpc824 (
      {stage0_16[107]},
      {stage1_16[68]}
   );
   gpc1_1 gpc825 (
      {stage0_16[108]},
      {stage1_16[69]}
   );
   gpc1_1 gpc826 (
      {stage0_16[109]},
      {stage1_16[70]}
   );
   gpc1_1 gpc827 (
      {stage0_16[110]},
      {stage1_16[71]}
   );
   gpc1_1 gpc828 (
      {stage0_16[111]},
      {stage1_16[72]}
   );
   gpc1_1 gpc829 (
      {stage0_16[112]},
      {stage1_16[73]}
   );
   gpc1_1 gpc830 (
      {stage0_16[113]},
      {stage1_16[74]}
   );
   gpc1_1 gpc831 (
      {stage0_16[114]},
      {stage1_16[75]}
   );
   gpc1_1 gpc832 (
      {stage0_16[115]},
      {stage1_16[76]}
   );
   gpc1_1 gpc833 (
      {stage0_16[116]},
      {stage1_16[77]}
   );
   gpc1_1 gpc834 (
      {stage0_16[117]},
      {stage1_16[78]}
   );
   gpc1_1 gpc835 (
      {stage0_16[118]},
      {stage1_16[79]}
   );
   gpc1_1 gpc836 (
      {stage0_16[119]},
      {stage1_16[80]}
   );
   gpc1_1 gpc837 (
      {stage0_16[120]},
      {stage1_16[81]}
   );
   gpc1_1 gpc838 (
      {stage0_16[121]},
      {stage1_16[82]}
   );
   gpc1_1 gpc839 (
      {stage0_16[122]},
      {stage1_16[83]}
   );
   gpc1_1 gpc840 (
      {stage0_16[123]},
      {stage1_16[84]}
   );
   gpc1_1 gpc841 (
      {stage0_16[124]},
      {stage1_16[85]}
   );
   gpc1_1 gpc842 (
      {stage0_16[125]},
      {stage1_16[86]}
   );
   gpc1_1 gpc843 (
      {stage0_16[126]},
      {stage1_16[87]}
   );
   gpc1_1 gpc844 (
      {stage0_16[127]},
      {stage1_16[88]}
   );
   gpc1_1 gpc845 (
      {stage0_17[103]},
      {stage1_17[42]}
   );
   gpc1_1 gpc846 (
      {stage0_17[104]},
      {stage1_17[43]}
   );
   gpc1_1 gpc847 (
      {stage0_17[105]},
      {stage1_17[44]}
   );
   gpc1_1 gpc848 (
      {stage0_17[106]},
      {stage1_17[45]}
   );
   gpc1_1 gpc849 (
      {stage0_17[107]},
      {stage1_17[46]}
   );
   gpc1_1 gpc850 (
      {stage0_17[108]},
      {stage1_17[47]}
   );
   gpc1_1 gpc851 (
      {stage0_17[109]},
      {stage1_17[48]}
   );
   gpc1_1 gpc852 (
      {stage0_17[110]},
      {stage1_17[49]}
   );
   gpc1_1 gpc853 (
      {stage0_17[111]},
      {stage1_17[50]}
   );
   gpc1_1 gpc854 (
      {stage0_17[112]},
      {stage1_17[51]}
   );
   gpc1_1 gpc855 (
      {stage0_17[113]},
      {stage1_17[52]}
   );
   gpc1_1 gpc856 (
      {stage0_17[114]},
      {stage1_17[53]}
   );
   gpc1_1 gpc857 (
      {stage0_17[115]},
      {stage1_17[54]}
   );
   gpc1_1 gpc858 (
      {stage0_17[116]},
      {stage1_17[55]}
   );
   gpc1_1 gpc859 (
      {stage0_17[117]},
      {stage1_17[56]}
   );
   gpc1_1 gpc860 (
      {stage0_17[118]},
      {stage1_17[57]}
   );
   gpc1_1 gpc861 (
      {stage0_17[119]},
      {stage1_17[58]}
   );
   gpc1_1 gpc862 (
      {stage0_17[120]},
      {stage1_17[59]}
   );
   gpc1_1 gpc863 (
      {stage0_17[121]},
      {stage1_17[60]}
   );
   gpc1_1 gpc864 (
      {stage0_17[122]},
      {stage1_17[61]}
   );
   gpc1_1 gpc865 (
      {stage0_17[123]},
      {stage1_17[62]}
   );
   gpc1_1 gpc866 (
      {stage0_17[124]},
      {stage1_17[63]}
   );
   gpc1_1 gpc867 (
      {stage0_17[125]},
      {stage1_17[64]}
   );
   gpc1_1 gpc868 (
      {stage0_17[126]},
      {stage1_17[65]}
   );
   gpc1_1 gpc869 (
      {stage0_17[127]},
      {stage1_17[66]}
   );
   gpc1_1 gpc870 (
      {stage0_19[123]},
      {stage1_19[50]}
   );
   gpc1_1 gpc871 (
      {stage0_19[124]},
      {stage1_19[51]}
   );
   gpc1_1 gpc872 (
      {stage0_19[125]},
      {stage1_19[52]}
   );
   gpc1_1 gpc873 (
      {stage0_19[126]},
      {stage1_19[53]}
   );
   gpc1_1 gpc874 (
      {stage0_19[127]},
      {stage1_19[54]}
   );
   gpc1_1 gpc875 (
      {stage0_20[104]},
      {stage1_20[48]}
   );
   gpc1_1 gpc876 (
      {stage0_20[105]},
      {stage1_20[49]}
   );
   gpc1_1 gpc877 (
      {stage0_20[106]},
      {stage1_20[50]}
   );
   gpc1_1 gpc878 (
      {stage0_20[107]},
      {stage1_20[51]}
   );
   gpc1_1 gpc879 (
      {stage0_20[108]},
      {stage1_20[52]}
   );
   gpc1_1 gpc880 (
      {stage0_20[109]},
      {stage1_20[53]}
   );
   gpc1_1 gpc881 (
      {stage0_20[110]},
      {stage1_20[54]}
   );
   gpc1_1 gpc882 (
      {stage0_20[111]},
      {stage1_20[55]}
   );
   gpc1_1 gpc883 (
      {stage0_20[112]},
      {stage1_20[56]}
   );
   gpc1_1 gpc884 (
      {stage0_20[113]},
      {stage1_20[57]}
   );
   gpc1_1 gpc885 (
      {stage0_20[114]},
      {stage1_20[58]}
   );
   gpc1_1 gpc886 (
      {stage0_20[115]},
      {stage1_20[59]}
   );
   gpc1_1 gpc887 (
      {stage0_20[116]},
      {stage1_20[60]}
   );
   gpc1_1 gpc888 (
      {stage0_20[117]},
      {stage1_20[61]}
   );
   gpc1_1 gpc889 (
      {stage0_20[118]},
      {stage1_20[62]}
   );
   gpc1_1 gpc890 (
      {stage0_20[119]},
      {stage1_20[63]}
   );
   gpc1_1 gpc891 (
      {stage0_20[120]},
      {stage1_20[64]}
   );
   gpc1_1 gpc892 (
      {stage0_20[121]},
      {stage1_20[65]}
   );
   gpc1_1 gpc893 (
      {stage0_20[122]},
      {stage1_20[66]}
   );
   gpc1_1 gpc894 (
      {stage0_20[123]},
      {stage1_20[67]}
   );
   gpc1_1 gpc895 (
      {stage0_20[124]},
      {stage1_20[68]}
   );
   gpc1_1 gpc896 (
      {stage0_20[125]},
      {stage1_20[69]}
   );
   gpc1_1 gpc897 (
      {stage0_20[126]},
      {stage1_20[70]}
   );
   gpc1_1 gpc898 (
      {stage0_20[127]},
      {stage1_20[71]}
   );
   gpc1_1 gpc899 (
      {stage0_21[121]},
      {stage1_21[48]}
   );
   gpc1_1 gpc900 (
      {stage0_21[122]},
      {stage1_21[49]}
   );
   gpc1_1 gpc901 (
      {stage0_21[123]},
      {stage1_21[50]}
   );
   gpc1_1 gpc902 (
      {stage0_21[124]},
      {stage1_21[51]}
   );
   gpc1_1 gpc903 (
      {stage0_21[125]},
      {stage1_21[52]}
   );
   gpc1_1 gpc904 (
      {stage0_21[126]},
      {stage1_21[53]}
   );
   gpc1_1 gpc905 (
      {stage0_21[127]},
      {stage1_21[54]}
   );
   gpc1_1 gpc906 (
      {stage0_22[106]},
      {stage1_22[49]}
   );
   gpc1_1 gpc907 (
      {stage0_22[107]},
      {stage1_22[50]}
   );
   gpc1_1 gpc908 (
      {stage0_22[108]},
      {stage1_22[51]}
   );
   gpc1_1 gpc909 (
      {stage0_22[109]},
      {stage1_22[52]}
   );
   gpc1_1 gpc910 (
      {stage0_22[110]},
      {stage1_22[53]}
   );
   gpc1_1 gpc911 (
      {stage0_22[111]},
      {stage1_22[54]}
   );
   gpc1_1 gpc912 (
      {stage0_22[112]},
      {stage1_22[55]}
   );
   gpc1_1 gpc913 (
      {stage0_22[113]},
      {stage1_22[56]}
   );
   gpc1_1 gpc914 (
      {stage0_22[114]},
      {stage1_22[57]}
   );
   gpc1_1 gpc915 (
      {stage0_22[115]},
      {stage1_22[58]}
   );
   gpc1_1 gpc916 (
      {stage0_22[116]},
      {stage1_22[59]}
   );
   gpc1_1 gpc917 (
      {stage0_22[117]},
      {stage1_22[60]}
   );
   gpc1_1 gpc918 (
      {stage0_22[118]},
      {stage1_22[61]}
   );
   gpc1_1 gpc919 (
      {stage0_22[119]},
      {stage1_22[62]}
   );
   gpc1_1 gpc920 (
      {stage0_22[120]},
      {stage1_22[63]}
   );
   gpc1_1 gpc921 (
      {stage0_22[121]},
      {stage1_22[64]}
   );
   gpc1_1 gpc922 (
      {stage0_22[122]},
      {stage1_22[65]}
   );
   gpc1_1 gpc923 (
      {stage0_22[123]},
      {stage1_22[66]}
   );
   gpc1_1 gpc924 (
      {stage0_22[124]},
      {stage1_22[67]}
   );
   gpc1_1 gpc925 (
      {stage0_22[125]},
      {stage1_22[68]}
   );
   gpc1_1 gpc926 (
      {stage0_22[126]},
      {stage1_22[69]}
   );
   gpc1_1 gpc927 (
      {stage0_22[127]},
      {stage1_22[70]}
   );
   gpc1_1 gpc928 (
      {stage0_23[122]},
      {stage1_23[48]}
   );
   gpc1_1 gpc929 (
      {stage0_23[123]},
      {stage1_23[49]}
   );
   gpc1_1 gpc930 (
      {stage0_23[124]},
      {stage1_23[50]}
   );
   gpc1_1 gpc931 (
      {stage0_23[125]},
      {stage1_23[51]}
   );
   gpc1_1 gpc932 (
      {stage0_23[126]},
      {stage1_23[52]}
   );
   gpc1_1 gpc933 (
      {stage0_23[127]},
      {stage1_23[53]}
   );
   gpc1_1 gpc934 (
      {stage0_24[109]},
      {stage1_24[43]}
   );
   gpc1_1 gpc935 (
      {stage0_24[110]},
      {stage1_24[44]}
   );
   gpc1_1 gpc936 (
      {stage0_24[111]},
      {stage1_24[45]}
   );
   gpc1_1 gpc937 (
      {stage0_24[112]},
      {stage1_24[46]}
   );
   gpc1_1 gpc938 (
      {stage0_24[113]},
      {stage1_24[47]}
   );
   gpc1_1 gpc939 (
      {stage0_24[114]},
      {stage1_24[48]}
   );
   gpc1_1 gpc940 (
      {stage0_24[115]},
      {stage1_24[49]}
   );
   gpc1_1 gpc941 (
      {stage0_24[116]},
      {stage1_24[50]}
   );
   gpc1_1 gpc942 (
      {stage0_24[117]},
      {stage1_24[51]}
   );
   gpc1_1 gpc943 (
      {stage0_24[118]},
      {stage1_24[52]}
   );
   gpc1_1 gpc944 (
      {stage0_24[119]},
      {stage1_24[53]}
   );
   gpc1_1 gpc945 (
      {stage0_24[120]},
      {stage1_24[54]}
   );
   gpc1_1 gpc946 (
      {stage0_24[121]},
      {stage1_24[55]}
   );
   gpc1_1 gpc947 (
      {stage0_24[122]},
      {stage1_24[56]}
   );
   gpc1_1 gpc948 (
      {stage0_24[123]},
      {stage1_24[57]}
   );
   gpc1_1 gpc949 (
      {stage0_24[124]},
      {stage1_24[58]}
   );
   gpc1_1 gpc950 (
      {stage0_24[125]},
      {stage1_24[59]}
   );
   gpc1_1 gpc951 (
      {stage0_24[126]},
      {stage1_24[60]}
   );
   gpc1_1 gpc952 (
      {stage0_24[127]},
      {stage1_24[61]}
   );
   gpc1_1 gpc953 (
      {stage0_25[114]},
      {stage1_25[47]}
   );
   gpc1_1 gpc954 (
      {stage0_25[115]},
      {stage1_25[48]}
   );
   gpc1_1 gpc955 (
      {stage0_25[116]},
      {stage1_25[49]}
   );
   gpc1_1 gpc956 (
      {stage0_25[117]},
      {stage1_25[50]}
   );
   gpc1_1 gpc957 (
      {stage0_25[118]},
      {stage1_25[51]}
   );
   gpc1_1 gpc958 (
      {stage0_25[119]},
      {stage1_25[52]}
   );
   gpc1_1 gpc959 (
      {stage0_25[120]},
      {stage1_25[53]}
   );
   gpc1_1 gpc960 (
      {stage0_25[121]},
      {stage1_25[54]}
   );
   gpc1_1 gpc961 (
      {stage0_25[122]},
      {stage1_25[55]}
   );
   gpc1_1 gpc962 (
      {stage0_25[123]},
      {stage1_25[56]}
   );
   gpc1_1 gpc963 (
      {stage0_25[124]},
      {stage1_25[57]}
   );
   gpc1_1 gpc964 (
      {stage0_25[125]},
      {stage1_25[58]}
   );
   gpc1_1 gpc965 (
      {stage0_25[126]},
      {stage1_25[59]}
   );
   gpc1_1 gpc966 (
      {stage0_25[127]},
      {stage1_25[60]}
   );
   gpc1_1 gpc967 (
      {stage0_26[93]},
      {stage1_26[49]}
   );
   gpc1_1 gpc968 (
      {stage0_26[94]},
      {stage1_26[50]}
   );
   gpc1_1 gpc969 (
      {stage0_26[95]},
      {stage1_26[51]}
   );
   gpc1_1 gpc970 (
      {stage0_26[96]},
      {stage1_26[52]}
   );
   gpc1_1 gpc971 (
      {stage0_26[97]},
      {stage1_26[53]}
   );
   gpc1_1 gpc972 (
      {stage0_26[98]},
      {stage1_26[54]}
   );
   gpc1_1 gpc973 (
      {stage0_26[99]},
      {stage1_26[55]}
   );
   gpc1_1 gpc974 (
      {stage0_26[100]},
      {stage1_26[56]}
   );
   gpc1_1 gpc975 (
      {stage0_26[101]},
      {stage1_26[57]}
   );
   gpc1_1 gpc976 (
      {stage0_26[102]},
      {stage1_26[58]}
   );
   gpc1_1 gpc977 (
      {stage0_26[103]},
      {stage1_26[59]}
   );
   gpc1_1 gpc978 (
      {stage0_26[104]},
      {stage1_26[60]}
   );
   gpc1_1 gpc979 (
      {stage0_26[105]},
      {stage1_26[61]}
   );
   gpc1_1 gpc980 (
      {stage0_26[106]},
      {stage1_26[62]}
   );
   gpc1_1 gpc981 (
      {stage0_26[107]},
      {stage1_26[63]}
   );
   gpc1_1 gpc982 (
      {stage0_26[108]},
      {stage1_26[64]}
   );
   gpc1_1 gpc983 (
      {stage0_26[109]},
      {stage1_26[65]}
   );
   gpc1_1 gpc984 (
      {stage0_26[110]},
      {stage1_26[66]}
   );
   gpc1_1 gpc985 (
      {stage0_26[111]},
      {stage1_26[67]}
   );
   gpc1_1 gpc986 (
      {stage0_26[112]},
      {stage1_26[68]}
   );
   gpc1_1 gpc987 (
      {stage0_26[113]},
      {stage1_26[69]}
   );
   gpc1_1 gpc988 (
      {stage0_26[114]},
      {stage1_26[70]}
   );
   gpc1_1 gpc989 (
      {stage0_26[115]},
      {stage1_26[71]}
   );
   gpc1_1 gpc990 (
      {stage0_26[116]},
      {stage1_26[72]}
   );
   gpc1_1 gpc991 (
      {stage0_26[117]},
      {stage1_26[73]}
   );
   gpc1_1 gpc992 (
      {stage0_26[118]},
      {stage1_26[74]}
   );
   gpc1_1 gpc993 (
      {stage0_26[119]},
      {stage1_26[75]}
   );
   gpc1_1 gpc994 (
      {stage0_26[120]},
      {stage1_26[76]}
   );
   gpc1_1 gpc995 (
      {stage0_26[121]},
      {stage1_26[77]}
   );
   gpc1_1 gpc996 (
      {stage0_26[122]},
      {stage1_26[78]}
   );
   gpc1_1 gpc997 (
      {stage0_26[123]},
      {stage1_26[79]}
   );
   gpc1_1 gpc998 (
      {stage0_26[124]},
      {stage1_26[80]}
   );
   gpc1_1 gpc999 (
      {stage0_26[125]},
      {stage1_26[81]}
   );
   gpc1_1 gpc1000 (
      {stage0_26[126]},
      {stage1_26[82]}
   );
   gpc1_1 gpc1001 (
      {stage0_26[127]},
      {stage1_26[83]}
   );
   gpc1_1 gpc1002 (
      {stage0_27[114]},
      {stage1_27[42]}
   );
   gpc1_1 gpc1003 (
      {stage0_27[115]},
      {stage1_27[43]}
   );
   gpc1_1 gpc1004 (
      {stage0_27[116]},
      {stage1_27[44]}
   );
   gpc1_1 gpc1005 (
      {stage0_27[117]},
      {stage1_27[45]}
   );
   gpc1_1 gpc1006 (
      {stage0_27[118]},
      {stage1_27[46]}
   );
   gpc1_1 gpc1007 (
      {stage0_27[119]},
      {stage1_27[47]}
   );
   gpc1_1 gpc1008 (
      {stage0_27[120]},
      {stage1_27[48]}
   );
   gpc1_1 gpc1009 (
      {stage0_27[121]},
      {stage1_27[49]}
   );
   gpc1_1 gpc1010 (
      {stage0_27[122]},
      {stage1_27[50]}
   );
   gpc1_1 gpc1011 (
      {stage0_27[123]},
      {stage1_27[51]}
   );
   gpc1_1 gpc1012 (
      {stage0_27[124]},
      {stage1_27[52]}
   );
   gpc1_1 gpc1013 (
      {stage0_27[125]},
      {stage1_27[53]}
   );
   gpc1_1 gpc1014 (
      {stage0_27[126]},
      {stage1_27[54]}
   );
   gpc1_1 gpc1015 (
      {stage0_27[127]},
      {stage1_27[55]}
   );
   gpc1_1 gpc1016 (
      {stage0_28[126]},
      {stage1_28[46]}
   );
   gpc1_1 gpc1017 (
      {stage0_28[127]},
      {stage1_28[47]}
   );
   gpc1_1 gpc1018 (
      {stage0_29[99]},
      {stage1_29[51]}
   );
   gpc1_1 gpc1019 (
      {stage0_29[100]},
      {stage1_29[52]}
   );
   gpc1_1 gpc1020 (
      {stage0_29[101]},
      {stage1_29[53]}
   );
   gpc1_1 gpc1021 (
      {stage0_29[102]},
      {stage1_29[54]}
   );
   gpc1_1 gpc1022 (
      {stage0_29[103]},
      {stage1_29[55]}
   );
   gpc1_1 gpc1023 (
      {stage0_29[104]},
      {stage1_29[56]}
   );
   gpc1_1 gpc1024 (
      {stage0_29[105]},
      {stage1_29[57]}
   );
   gpc1_1 gpc1025 (
      {stage0_29[106]},
      {stage1_29[58]}
   );
   gpc1_1 gpc1026 (
      {stage0_29[107]},
      {stage1_29[59]}
   );
   gpc1_1 gpc1027 (
      {stage0_29[108]},
      {stage1_29[60]}
   );
   gpc1_1 gpc1028 (
      {stage0_29[109]},
      {stage1_29[61]}
   );
   gpc1_1 gpc1029 (
      {stage0_29[110]},
      {stage1_29[62]}
   );
   gpc1_1 gpc1030 (
      {stage0_29[111]},
      {stage1_29[63]}
   );
   gpc1_1 gpc1031 (
      {stage0_29[112]},
      {stage1_29[64]}
   );
   gpc1_1 gpc1032 (
      {stage0_29[113]},
      {stage1_29[65]}
   );
   gpc1_1 gpc1033 (
      {stage0_29[114]},
      {stage1_29[66]}
   );
   gpc1_1 gpc1034 (
      {stage0_29[115]},
      {stage1_29[67]}
   );
   gpc1_1 gpc1035 (
      {stage0_29[116]},
      {stage1_29[68]}
   );
   gpc1_1 gpc1036 (
      {stage0_29[117]},
      {stage1_29[69]}
   );
   gpc1_1 gpc1037 (
      {stage0_29[118]},
      {stage1_29[70]}
   );
   gpc1_1 gpc1038 (
      {stage0_29[119]},
      {stage1_29[71]}
   );
   gpc1_1 gpc1039 (
      {stage0_29[120]},
      {stage1_29[72]}
   );
   gpc1_1 gpc1040 (
      {stage0_29[121]},
      {stage1_29[73]}
   );
   gpc1_1 gpc1041 (
      {stage0_29[122]},
      {stage1_29[74]}
   );
   gpc1_1 gpc1042 (
      {stage0_29[123]},
      {stage1_29[75]}
   );
   gpc1_1 gpc1043 (
      {stage0_29[124]},
      {stage1_29[76]}
   );
   gpc1_1 gpc1044 (
      {stage0_29[125]},
      {stage1_29[77]}
   );
   gpc1_1 gpc1045 (
      {stage0_29[126]},
      {stage1_29[78]}
   );
   gpc1_1 gpc1046 (
      {stage0_29[127]},
      {stage1_29[79]}
   );
   gpc1_1 gpc1047 (
      {stage0_30[99]},
      {stage1_30[43]}
   );
   gpc1_1 gpc1048 (
      {stage0_30[100]},
      {stage1_30[44]}
   );
   gpc1_1 gpc1049 (
      {stage0_30[101]},
      {stage1_30[45]}
   );
   gpc1_1 gpc1050 (
      {stage0_30[102]},
      {stage1_30[46]}
   );
   gpc1_1 gpc1051 (
      {stage0_30[103]},
      {stage1_30[47]}
   );
   gpc1_1 gpc1052 (
      {stage0_30[104]},
      {stage1_30[48]}
   );
   gpc1_1 gpc1053 (
      {stage0_30[105]},
      {stage1_30[49]}
   );
   gpc1_1 gpc1054 (
      {stage0_30[106]},
      {stage1_30[50]}
   );
   gpc1_1 gpc1055 (
      {stage0_30[107]},
      {stage1_30[51]}
   );
   gpc1_1 gpc1056 (
      {stage0_30[108]},
      {stage1_30[52]}
   );
   gpc1_1 gpc1057 (
      {stage0_30[109]},
      {stage1_30[53]}
   );
   gpc1_1 gpc1058 (
      {stage0_30[110]},
      {stage1_30[54]}
   );
   gpc1_1 gpc1059 (
      {stage0_30[111]},
      {stage1_30[55]}
   );
   gpc1_1 gpc1060 (
      {stage0_30[112]},
      {stage1_30[56]}
   );
   gpc1_1 gpc1061 (
      {stage0_30[113]},
      {stage1_30[57]}
   );
   gpc1_1 gpc1062 (
      {stage0_30[114]},
      {stage1_30[58]}
   );
   gpc1_1 gpc1063 (
      {stage0_30[115]},
      {stage1_30[59]}
   );
   gpc1_1 gpc1064 (
      {stage0_30[116]},
      {stage1_30[60]}
   );
   gpc1_1 gpc1065 (
      {stage0_30[117]},
      {stage1_30[61]}
   );
   gpc1_1 gpc1066 (
      {stage0_30[118]},
      {stage1_30[62]}
   );
   gpc1_1 gpc1067 (
      {stage0_30[119]},
      {stage1_30[63]}
   );
   gpc1_1 gpc1068 (
      {stage0_30[120]},
      {stage1_30[64]}
   );
   gpc1_1 gpc1069 (
      {stage0_30[121]},
      {stage1_30[65]}
   );
   gpc1_1 gpc1070 (
      {stage0_30[122]},
      {stage1_30[66]}
   );
   gpc1_1 gpc1071 (
      {stage0_30[123]},
      {stage1_30[67]}
   );
   gpc1_1 gpc1072 (
      {stage0_30[124]},
      {stage1_30[68]}
   );
   gpc1_1 gpc1073 (
      {stage0_30[125]},
      {stage1_30[69]}
   );
   gpc1_1 gpc1074 (
      {stage0_30[126]},
      {stage1_30[70]}
   );
   gpc1_1 gpc1075 (
      {stage0_30[127]},
      {stage1_30[71]}
   );
   gpc1_1 gpc1076 (
      {stage0_31[109]},
      {stage1_31[41]}
   );
   gpc1_1 gpc1077 (
      {stage0_31[110]},
      {stage1_31[42]}
   );
   gpc1_1 gpc1078 (
      {stage0_31[111]},
      {stage1_31[43]}
   );
   gpc1_1 gpc1079 (
      {stage0_31[112]},
      {stage1_31[44]}
   );
   gpc1_1 gpc1080 (
      {stage0_31[113]},
      {stage1_31[45]}
   );
   gpc1_1 gpc1081 (
      {stage0_31[114]},
      {stage1_31[46]}
   );
   gpc1_1 gpc1082 (
      {stage0_31[115]},
      {stage1_31[47]}
   );
   gpc1_1 gpc1083 (
      {stage0_31[116]},
      {stage1_31[48]}
   );
   gpc1_1 gpc1084 (
      {stage0_31[117]},
      {stage1_31[49]}
   );
   gpc1_1 gpc1085 (
      {stage0_31[118]},
      {stage1_31[50]}
   );
   gpc1_1 gpc1086 (
      {stage0_31[119]},
      {stage1_31[51]}
   );
   gpc1_1 gpc1087 (
      {stage0_31[120]},
      {stage1_31[52]}
   );
   gpc1_1 gpc1088 (
      {stage0_31[121]},
      {stage1_31[53]}
   );
   gpc1_1 gpc1089 (
      {stage0_31[122]},
      {stage1_31[54]}
   );
   gpc1_1 gpc1090 (
      {stage0_31[123]},
      {stage1_31[55]}
   );
   gpc1_1 gpc1091 (
      {stage0_31[124]},
      {stage1_31[56]}
   );
   gpc1_1 gpc1092 (
      {stage0_31[125]},
      {stage1_31[57]}
   );
   gpc1_1 gpc1093 (
      {stage0_31[126]},
      {stage1_31[58]}
   );
   gpc1_1 gpc1094 (
      {stage0_31[127]},
      {stage1_31[59]}
   );
   gpc1_1 gpc1095 (
      {stage0_32[93]},
      {stage1_32[48]}
   );
   gpc1_1 gpc1096 (
      {stage0_32[94]},
      {stage1_32[49]}
   );
   gpc1_1 gpc1097 (
      {stage0_32[95]},
      {stage1_32[50]}
   );
   gpc1_1 gpc1098 (
      {stage0_32[96]},
      {stage1_32[51]}
   );
   gpc1_1 gpc1099 (
      {stage0_32[97]},
      {stage1_32[52]}
   );
   gpc1_1 gpc1100 (
      {stage0_32[98]},
      {stage1_32[53]}
   );
   gpc1_1 gpc1101 (
      {stage0_32[99]},
      {stage1_32[54]}
   );
   gpc1_1 gpc1102 (
      {stage0_32[100]},
      {stage1_32[55]}
   );
   gpc1_1 gpc1103 (
      {stage0_32[101]},
      {stage1_32[56]}
   );
   gpc1_1 gpc1104 (
      {stage0_32[102]},
      {stage1_32[57]}
   );
   gpc1_1 gpc1105 (
      {stage0_32[103]},
      {stage1_32[58]}
   );
   gpc1_1 gpc1106 (
      {stage0_32[104]},
      {stage1_32[59]}
   );
   gpc1_1 gpc1107 (
      {stage0_32[105]},
      {stage1_32[60]}
   );
   gpc1_1 gpc1108 (
      {stage0_32[106]},
      {stage1_32[61]}
   );
   gpc1_1 gpc1109 (
      {stage0_32[107]},
      {stage1_32[62]}
   );
   gpc1_1 gpc1110 (
      {stage0_32[108]},
      {stage1_32[63]}
   );
   gpc1_1 gpc1111 (
      {stage0_32[109]},
      {stage1_32[64]}
   );
   gpc1_1 gpc1112 (
      {stage0_32[110]},
      {stage1_32[65]}
   );
   gpc1_1 gpc1113 (
      {stage0_32[111]},
      {stage1_32[66]}
   );
   gpc1_1 gpc1114 (
      {stage0_32[112]},
      {stage1_32[67]}
   );
   gpc1_1 gpc1115 (
      {stage0_32[113]},
      {stage1_32[68]}
   );
   gpc1_1 gpc1116 (
      {stage0_32[114]},
      {stage1_32[69]}
   );
   gpc1_1 gpc1117 (
      {stage0_32[115]},
      {stage1_32[70]}
   );
   gpc1_1 gpc1118 (
      {stage0_32[116]},
      {stage1_32[71]}
   );
   gpc1_1 gpc1119 (
      {stage0_32[117]},
      {stage1_32[72]}
   );
   gpc1_1 gpc1120 (
      {stage0_32[118]},
      {stage1_32[73]}
   );
   gpc1_1 gpc1121 (
      {stage0_32[119]},
      {stage1_32[74]}
   );
   gpc1_1 gpc1122 (
      {stage0_32[120]},
      {stage1_32[75]}
   );
   gpc1_1 gpc1123 (
      {stage0_32[121]},
      {stage1_32[76]}
   );
   gpc1_1 gpc1124 (
      {stage0_32[122]},
      {stage1_32[77]}
   );
   gpc1_1 gpc1125 (
      {stage0_32[123]},
      {stage1_32[78]}
   );
   gpc1_1 gpc1126 (
      {stage0_32[124]},
      {stage1_32[79]}
   );
   gpc1_1 gpc1127 (
      {stage0_32[125]},
      {stage1_32[80]}
   );
   gpc1_1 gpc1128 (
      {stage0_32[126]},
      {stage1_32[81]}
   );
   gpc1_1 gpc1129 (
      {stage0_32[127]},
      {stage1_32[82]}
   );
   gpc1_1 gpc1130 (
      {stage0_33[109]},
      {stage1_33[44]}
   );
   gpc1_1 gpc1131 (
      {stage0_33[110]},
      {stage1_33[45]}
   );
   gpc1_1 gpc1132 (
      {stage0_33[111]},
      {stage1_33[46]}
   );
   gpc1_1 gpc1133 (
      {stage0_33[112]},
      {stage1_33[47]}
   );
   gpc1_1 gpc1134 (
      {stage0_33[113]},
      {stage1_33[48]}
   );
   gpc1_1 gpc1135 (
      {stage0_33[114]},
      {stage1_33[49]}
   );
   gpc1_1 gpc1136 (
      {stage0_33[115]},
      {stage1_33[50]}
   );
   gpc1_1 gpc1137 (
      {stage0_33[116]},
      {stage1_33[51]}
   );
   gpc1_1 gpc1138 (
      {stage0_33[117]},
      {stage1_33[52]}
   );
   gpc1_1 gpc1139 (
      {stage0_33[118]},
      {stage1_33[53]}
   );
   gpc1_1 gpc1140 (
      {stage0_33[119]},
      {stage1_33[54]}
   );
   gpc1_1 gpc1141 (
      {stage0_33[120]},
      {stage1_33[55]}
   );
   gpc1_1 gpc1142 (
      {stage0_33[121]},
      {stage1_33[56]}
   );
   gpc1_1 gpc1143 (
      {stage0_33[122]},
      {stage1_33[57]}
   );
   gpc1_1 gpc1144 (
      {stage0_33[123]},
      {stage1_33[58]}
   );
   gpc1_1 gpc1145 (
      {stage0_33[124]},
      {stage1_33[59]}
   );
   gpc1_1 gpc1146 (
      {stage0_33[125]},
      {stage1_33[60]}
   );
   gpc1_1 gpc1147 (
      {stage0_33[126]},
      {stage1_33[61]}
   );
   gpc1_1 gpc1148 (
      {stage0_33[127]},
      {stage1_33[62]}
   );
   gpc1_1 gpc1149 (
      {stage0_34[97]},
      {stage1_34[37]}
   );
   gpc1_1 gpc1150 (
      {stage0_34[98]},
      {stage1_34[38]}
   );
   gpc1_1 gpc1151 (
      {stage0_34[99]},
      {stage1_34[39]}
   );
   gpc1_1 gpc1152 (
      {stage0_34[100]},
      {stage1_34[40]}
   );
   gpc1_1 gpc1153 (
      {stage0_34[101]},
      {stage1_34[41]}
   );
   gpc1_1 gpc1154 (
      {stage0_34[102]},
      {stage1_34[42]}
   );
   gpc1_1 gpc1155 (
      {stage0_34[103]},
      {stage1_34[43]}
   );
   gpc1_1 gpc1156 (
      {stage0_34[104]},
      {stage1_34[44]}
   );
   gpc1_1 gpc1157 (
      {stage0_34[105]},
      {stage1_34[45]}
   );
   gpc1_1 gpc1158 (
      {stage0_34[106]},
      {stage1_34[46]}
   );
   gpc1_1 gpc1159 (
      {stage0_34[107]},
      {stage1_34[47]}
   );
   gpc1_1 gpc1160 (
      {stage0_34[108]},
      {stage1_34[48]}
   );
   gpc1_1 gpc1161 (
      {stage0_34[109]},
      {stage1_34[49]}
   );
   gpc1_1 gpc1162 (
      {stage0_34[110]},
      {stage1_34[50]}
   );
   gpc1_1 gpc1163 (
      {stage0_34[111]},
      {stage1_34[51]}
   );
   gpc1_1 gpc1164 (
      {stage0_34[112]},
      {stage1_34[52]}
   );
   gpc1_1 gpc1165 (
      {stage0_34[113]},
      {stage1_34[53]}
   );
   gpc1_1 gpc1166 (
      {stage0_34[114]},
      {stage1_34[54]}
   );
   gpc1_1 gpc1167 (
      {stage0_34[115]},
      {stage1_34[55]}
   );
   gpc1_1 gpc1168 (
      {stage0_34[116]},
      {stage1_34[56]}
   );
   gpc1_1 gpc1169 (
      {stage0_34[117]},
      {stage1_34[57]}
   );
   gpc1_1 gpc1170 (
      {stage0_34[118]},
      {stage1_34[58]}
   );
   gpc1_1 gpc1171 (
      {stage0_34[119]},
      {stage1_34[59]}
   );
   gpc1_1 gpc1172 (
      {stage0_34[120]},
      {stage1_34[60]}
   );
   gpc1_1 gpc1173 (
      {stage0_34[121]},
      {stage1_34[61]}
   );
   gpc1_1 gpc1174 (
      {stage0_34[122]},
      {stage1_34[62]}
   );
   gpc1_1 gpc1175 (
      {stage0_34[123]},
      {stage1_34[63]}
   );
   gpc1_1 gpc1176 (
      {stage0_34[124]},
      {stage1_34[64]}
   );
   gpc1_1 gpc1177 (
      {stage0_34[125]},
      {stage1_34[65]}
   );
   gpc1_1 gpc1178 (
      {stage0_34[126]},
      {stage1_34[66]}
   );
   gpc1_1 gpc1179 (
      {stage0_34[127]},
      {stage1_34[67]}
   );
   gpc1_1 gpc1180 (
      {stage0_35[127]},
      {stage1_35[47]}
   );
   gpc1_1 gpc1181 (
      {stage0_36[120]},
      {stage1_36[53]}
   );
   gpc1_1 gpc1182 (
      {stage0_36[121]},
      {stage1_36[54]}
   );
   gpc1_1 gpc1183 (
      {stage0_36[122]},
      {stage1_36[55]}
   );
   gpc1_1 gpc1184 (
      {stage0_36[123]},
      {stage1_36[56]}
   );
   gpc1_1 gpc1185 (
      {stage0_36[124]},
      {stage1_36[57]}
   );
   gpc1_1 gpc1186 (
      {stage0_36[125]},
      {stage1_36[58]}
   );
   gpc1_1 gpc1187 (
      {stage0_36[126]},
      {stage1_36[59]}
   );
   gpc1_1 gpc1188 (
      {stage0_36[127]},
      {stage1_36[60]}
   );
   gpc1_1 gpc1189 (
      {stage0_37[72]},
      {stage1_37[41]}
   );
   gpc1_1 gpc1190 (
      {stage0_37[73]},
      {stage1_37[42]}
   );
   gpc1_1 gpc1191 (
      {stage0_37[74]},
      {stage1_37[43]}
   );
   gpc1_1 gpc1192 (
      {stage0_37[75]},
      {stage1_37[44]}
   );
   gpc1_1 gpc1193 (
      {stage0_37[76]},
      {stage1_37[45]}
   );
   gpc1_1 gpc1194 (
      {stage0_37[77]},
      {stage1_37[46]}
   );
   gpc1_1 gpc1195 (
      {stage0_37[78]},
      {stage1_37[47]}
   );
   gpc1_1 gpc1196 (
      {stage0_37[79]},
      {stage1_37[48]}
   );
   gpc1_1 gpc1197 (
      {stage0_37[80]},
      {stage1_37[49]}
   );
   gpc1_1 gpc1198 (
      {stage0_37[81]},
      {stage1_37[50]}
   );
   gpc1_1 gpc1199 (
      {stage0_37[82]},
      {stage1_37[51]}
   );
   gpc1_1 gpc1200 (
      {stage0_37[83]},
      {stage1_37[52]}
   );
   gpc1_1 gpc1201 (
      {stage0_37[84]},
      {stage1_37[53]}
   );
   gpc1_1 gpc1202 (
      {stage0_37[85]},
      {stage1_37[54]}
   );
   gpc1_1 gpc1203 (
      {stage0_37[86]},
      {stage1_37[55]}
   );
   gpc1_1 gpc1204 (
      {stage0_37[87]},
      {stage1_37[56]}
   );
   gpc1_1 gpc1205 (
      {stage0_37[88]},
      {stage1_37[57]}
   );
   gpc1_1 gpc1206 (
      {stage0_37[89]},
      {stage1_37[58]}
   );
   gpc1_1 gpc1207 (
      {stage0_37[90]},
      {stage1_37[59]}
   );
   gpc1_1 gpc1208 (
      {stage0_37[91]},
      {stage1_37[60]}
   );
   gpc1_1 gpc1209 (
      {stage0_37[92]},
      {stage1_37[61]}
   );
   gpc1_1 gpc1210 (
      {stage0_37[93]},
      {stage1_37[62]}
   );
   gpc1_1 gpc1211 (
      {stage0_37[94]},
      {stage1_37[63]}
   );
   gpc1_1 gpc1212 (
      {stage0_37[95]},
      {stage1_37[64]}
   );
   gpc1_1 gpc1213 (
      {stage0_37[96]},
      {stage1_37[65]}
   );
   gpc1_1 gpc1214 (
      {stage0_37[97]},
      {stage1_37[66]}
   );
   gpc1_1 gpc1215 (
      {stage0_37[98]},
      {stage1_37[67]}
   );
   gpc1_1 gpc1216 (
      {stage0_37[99]},
      {stage1_37[68]}
   );
   gpc1_1 gpc1217 (
      {stage0_37[100]},
      {stage1_37[69]}
   );
   gpc1_1 gpc1218 (
      {stage0_37[101]},
      {stage1_37[70]}
   );
   gpc1_1 gpc1219 (
      {stage0_37[102]},
      {stage1_37[71]}
   );
   gpc1_1 gpc1220 (
      {stage0_37[103]},
      {stage1_37[72]}
   );
   gpc1_1 gpc1221 (
      {stage0_37[104]},
      {stage1_37[73]}
   );
   gpc1_1 gpc1222 (
      {stage0_37[105]},
      {stage1_37[74]}
   );
   gpc1_1 gpc1223 (
      {stage0_37[106]},
      {stage1_37[75]}
   );
   gpc1_1 gpc1224 (
      {stage0_37[107]},
      {stage1_37[76]}
   );
   gpc1_1 gpc1225 (
      {stage0_37[108]},
      {stage1_37[77]}
   );
   gpc1_1 gpc1226 (
      {stage0_37[109]},
      {stage1_37[78]}
   );
   gpc1_1 gpc1227 (
      {stage0_37[110]},
      {stage1_37[79]}
   );
   gpc1_1 gpc1228 (
      {stage0_37[111]},
      {stage1_37[80]}
   );
   gpc1_1 gpc1229 (
      {stage0_37[112]},
      {stage1_37[81]}
   );
   gpc1_1 gpc1230 (
      {stage0_37[113]},
      {stage1_37[82]}
   );
   gpc1_1 gpc1231 (
      {stage0_37[114]},
      {stage1_37[83]}
   );
   gpc1_1 gpc1232 (
      {stage0_37[115]},
      {stage1_37[84]}
   );
   gpc1_1 gpc1233 (
      {stage0_37[116]},
      {stage1_37[85]}
   );
   gpc1_1 gpc1234 (
      {stage0_37[117]},
      {stage1_37[86]}
   );
   gpc1_1 gpc1235 (
      {stage0_37[118]},
      {stage1_37[87]}
   );
   gpc1_1 gpc1236 (
      {stage0_37[119]},
      {stage1_37[88]}
   );
   gpc1_1 gpc1237 (
      {stage0_37[120]},
      {stage1_37[89]}
   );
   gpc1_1 gpc1238 (
      {stage0_37[121]},
      {stage1_37[90]}
   );
   gpc1_1 gpc1239 (
      {stage0_37[122]},
      {stage1_37[91]}
   );
   gpc1_1 gpc1240 (
      {stage0_37[123]},
      {stage1_37[92]}
   );
   gpc1_1 gpc1241 (
      {stage0_37[124]},
      {stage1_37[93]}
   );
   gpc1_1 gpc1242 (
      {stage0_37[125]},
      {stage1_37[94]}
   );
   gpc1_1 gpc1243 (
      {stage0_37[126]},
      {stage1_37[95]}
   );
   gpc1_1 gpc1244 (
      {stage0_37[127]},
      {stage1_37[96]}
   );
   gpc1_1 gpc1245 (
      {stage0_38[120]},
      {stage1_38[36]}
   );
   gpc1_1 gpc1246 (
      {stage0_38[121]},
      {stage1_38[37]}
   );
   gpc1_1 gpc1247 (
      {stage0_38[122]},
      {stage1_38[38]}
   );
   gpc1_1 gpc1248 (
      {stage0_38[123]},
      {stage1_38[39]}
   );
   gpc1_1 gpc1249 (
      {stage0_38[124]},
      {stage1_38[40]}
   );
   gpc1_1 gpc1250 (
      {stage0_38[125]},
      {stage1_38[41]}
   );
   gpc1_1 gpc1251 (
      {stage0_38[126]},
      {stage1_38[42]}
   );
   gpc1_1 gpc1252 (
      {stage0_38[127]},
      {stage1_38[43]}
   );
   gpc1_1 gpc1253 (
      {stage0_39[83]},
      {stage1_39[48]}
   );
   gpc1_1 gpc1254 (
      {stage0_39[84]},
      {stage1_39[49]}
   );
   gpc1_1 gpc1255 (
      {stage0_39[85]},
      {stage1_39[50]}
   );
   gpc1_1 gpc1256 (
      {stage0_39[86]},
      {stage1_39[51]}
   );
   gpc1_1 gpc1257 (
      {stage0_39[87]},
      {stage1_39[52]}
   );
   gpc1_1 gpc1258 (
      {stage0_39[88]},
      {stage1_39[53]}
   );
   gpc1_1 gpc1259 (
      {stage0_39[89]},
      {stage1_39[54]}
   );
   gpc1_1 gpc1260 (
      {stage0_39[90]},
      {stage1_39[55]}
   );
   gpc1_1 gpc1261 (
      {stage0_39[91]},
      {stage1_39[56]}
   );
   gpc1_1 gpc1262 (
      {stage0_39[92]},
      {stage1_39[57]}
   );
   gpc1_1 gpc1263 (
      {stage0_39[93]},
      {stage1_39[58]}
   );
   gpc1_1 gpc1264 (
      {stage0_39[94]},
      {stage1_39[59]}
   );
   gpc1_1 gpc1265 (
      {stage0_39[95]},
      {stage1_39[60]}
   );
   gpc1_1 gpc1266 (
      {stage0_39[96]},
      {stage1_39[61]}
   );
   gpc1_1 gpc1267 (
      {stage0_39[97]},
      {stage1_39[62]}
   );
   gpc1_1 gpc1268 (
      {stage0_39[98]},
      {stage1_39[63]}
   );
   gpc1_1 gpc1269 (
      {stage0_39[99]},
      {stage1_39[64]}
   );
   gpc1_1 gpc1270 (
      {stage0_39[100]},
      {stage1_39[65]}
   );
   gpc1_1 gpc1271 (
      {stage0_39[101]},
      {stage1_39[66]}
   );
   gpc1_1 gpc1272 (
      {stage0_39[102]},
      {stage1_39[67]}
   );
   gpc1_1 gpc1273 (
      {stage0_39[103]},
      {stage1_39[68]}
   );
   gpc1_1 gpc1274 (
      {stage0_39[104]},
      {stage1_39[69]}
   );
   gpc1_1 gpc1275 (
      {stage0_39[105]},
      {stage1_39[70]}
   );
   gpc1_1 gpc1276 (
      {stage0_39[106]},
      {stage1_39[71]}
   );
   gpc1_1 gpc1277 (
      {stage0_39[107]},
      {stage1_39[72]}
   );
   gpc1_1 gpc1278 (
      {stage0_39[108]},
      {stage1_39[73]}
   );
   gpc1_1 gpc1279 (
      {stage0_39[109]},
      {stage1_39[74]}
   );
   gpc1_1 gpc1280 (
      {stage0_39[110]},
      {stage1_39[75]}
   );
   gpc1_1 gpc1281 (
      {stage0_39[111]},
      {stage1_39[76]}
   );
   gpc1_1 gpc1282 (
      {stage0_39[112]},
      {stage1_39[77]}
   );
   gpc1_1 gpc1283 (
      {stage0_39[113]},
      {stage1_39[78]}
   );
   gpc1_1 gpc1284 (
      {stage0_39[114]},
      {stage1_39[79]}
   );
   gpc1_1 gpc1285 (
      {stage0_39[115]},
      {stage1_39[80]}
   );
   gpc1_1 gpc1286 (
      {stage0_39[116]},
      {stage1_39[81]}
   );
   gpc1_1 gpc1287 (
      {stage0_39[117]},
      {stage1_39[82]}
   );
   gpc1_1 gpc1288 (
      {stage0_39[118]},
      {stage1_39[83]}
   );
   gpc1_1 gpc1289 (
      {stage0_39[119]},
      {stage1_39[84]}
   );
   gpc1_1 gpc1290 (
      {stage0_39[120]},
      {stage1_39[85]}
   );
   gpc1_1 gpc1291 (
      {stage0_39[121]},
      {stage1_39[86]}
   );
   gpc1_1 gpc1292 (
      {stage0_39[122]},
      {stage1_39[87]}
   );
   gpc1_1 gpc1293 (
      {stage0_39[123]},
      {stage1_39[88]}
   );
   gpc1_1 gpc1294 (
      {stage0_39[124]},
      {stage1_39[89]}
   );
   gpc1_1 gpc1295 (
      {stage0_39[125]},
      {stage1_39[90]}
   );
   gpc1_1 gpc1296 (
      {stage0_39[126]},
      {stage1_39[91]}
   );
   gpc1_1 gpc1297 (
      {stage0_39[127]},
      {stage1_39[92]}
   );
   gpc1_1 gpc1298 (
      {stage0_40[112]},
      {stage1_40[47]}
   );
   gpc1_1 gpc1299 (
      {stage0_40[113]},
      {stage1_40[48]}
   );
   gpc1_1 gpc1300 (
      {stage0_40[114]},
      {stage1_40[49]}
   );
   gpc1_1 gpc1301 (
      {stage0_40[115]},
      {stage1_40[50]}
   );
   gpc1_1 gpc1302 (
      {stage0_40[116]},
      {stage1_40[51]}
   );
   gpc1_1 gpc1303 (
      {stage0_40[117]},
      {stage1_40[52]}
   );
   gpc1_1 gpc1304 (
      {stage0_40[118]},
      {stage1_40[53]}
   );
   gpc1_1 gpc1305 (
      {stage0_40[119]},
      {stage1_40[54]}
   );
   gpc1_1 gpc1306 (
      {stage0_40[120]},
      {stage1_40[55]}
   );
   gpc1_1 gpc1307 (
      {stage0_40[121]},
      {stage1_40[56]}
   );
   gpc1_1 gpc1308 (
      {stage0_40[122]},
      {stage1_40[57]}
   );
   gpc1_1 gpc1309 (
      {stage0_40[123]},
      {stage1_40[58]}
   );
   gpc1_1 gpc1310 (
      {stage0_40[124]},
      {stage1_40[59]}
   );
   gpc1_1 gpc1311 (
      {stage0_40[125]},
      {stage1_40[60]}
   );
   gpc1_1 gpc1312 (
      {stage0_40[126]},
      {stage1_40[61]}
   );
   gpc1_1 gpc1313 (
      {stage0_40[127]},
      {stage1_40[62]}
   );
   gpc1_1 gpc1314 (
      {stage0_41[126]},
      {stage1_41[38]}
   );
   gpc1_1 gpc1315 (
      {stage0_41[127]},
      {stage1_41[39]}
   );
   gpc1_1 gpc1316 (
      {stage0_42[127]},
      {stage1_42[50]}
   );
   gpc1_1 gpc1317 (
      {stage0_43[104]},
      {stage1_43[55]}
   );
   gpc1_1 gpc1318 (
      {stage0_43[105]},
      {stage1_43[56]}
   );
   gpc1_1 gpc1319 (
      {stage0_43[106]},
      {stage1_43[57]}
   );
   gpc1_1 gpc1320 (
      {stage0_43[107]},
      {stage1_43[58]}
   );
   gpc1_1 gpc1321 (
      {stage0_43[108]},
      {stage1_43[59]}
   );
   gpc1_1 gpc1322 (
      {stage0_43[109]},
      {stage1_43[60]}
   );
   gpc1_1 gpc1323 (
      {stage0_43[110]},
      {stage1_43[61]}
   );
   gpc1_1 gpc1324 (
      {stage0_43[111]},
      {stage1_43[62]}
   );
   gpc1_1 gpc1325 (
      {stage0_43[112]},
      {stage1_43[63]}
   );
   gpc1_1 gpc1326 (
      {stage0_43[113]},
      {stage1_43[64]}
   );
   gpc1_1 gpc1327 (
      {stage0_43[114]},
      {stage1_43[65]}
   );
   gpc1_1 gpc1328 (
      {stage0_43[115]},
      {stage1_43[66]}
   );
   gpc1_1 gpc1329 (
      {stage0_43[116]},
      {stage1_43[67]}
   );
   gpc1_1 gpc1330 (
      {stage0_43[117]},
      {stage1_43[68]}
   );
   gpc1_1 gpc1331 (
      {stage0_43[118]},
      {stage1_43[69]}
   );
   gpc1_1 gpc1332 (
      {stage0_43[119]},
      {stage1_43[70]}
   );
   gpc1_1 gpc1333 (
      {stage0_43[120]},
      {stage1_43[71]}
   );
   gpc1_1 gpc1334 (
      {stage0_43[121]},
      {stage1_43[72]}
   );
   gpc1_1 gpc1335 (
      {stage0_43[122]},
      {stage1_43[73]}
   );
   gpc1_1 gpc1336 (
      {stage0_43[123]},
      {stage1_43[74]}
   );
   gpc1_1 gpc1337 (
      {stage0_43[124]},
      {stage1_43[75]}
   );
   gpc1_1 gpc1338 (
      {stage0_43[125]},
      {stage1_43[76]}
   );
   gpc1_1 gpc1339 (
      {stage0_43[126]},
      {stage1_43[77]}
   );
   gpc1_1 gpc1340 (
      {stage0_43[127]},
      {stage1_43[78]}
   );
   gpc1_1 gpc1341 (
      {stage0_44[125]},
      {stage1_44[47]}
   );
   gpc1_1 gpc1342 (
      {stage0_44[126]},
      {stage1_44[48]}
   );
   gpc1_1 gpc1343 (
      {stage0_44[127]},
      {stage1_44[49]}
   );
   gpc1_1 gpc1344 (
      {stage0_45[114]},
      {stage1_45[44]}
   );
   gpc1_1 gpc1345 (
      {stage0_45[115]},
      {stage1_45[45]}
   );
   gpc1_1 gpc1346 (
      {stage0_45[116]},
      {stage1_45[46]}
   );
   gpc1_1 gpc1347 (
      {stage0_45[117]},
      {stage1_45[47]}
   );
   gpc1_1 gpc1348 (
      {stage0_45[118]},
      {stage1_45[48]}
   );
   gpc1_1 gpc1349 (
      {stage0_45[119]},
      {stage1_45[49]}
   );
   gpc1_1 gpc1350 (
      {stage0_45[120]},
      {stage1_45[50]}
   );
   gpc1_1 gpc1351 (
      {stage0_45[121]},
      {stage1_45[51]}
   );
   gpc1_1 gpc1352 (
      {stage0_45[122]},
      {stage1_45[52]}
   );
   gpc1_1 gpc1353 (
      {stage0_45[123]},
      {stage1_45[53]}
   );
   gpc1_1 gpc1354 (
      {stage0_45[124]},
      {stage1_45[54]}
   );
   gpc1_1 gpc1355 (
      {stage0_45[125]},
      {stage1_45[55]}
   );
   gpc1_1 gpc1356 (
      {stage0_45[126]},
      {stage1_45[56]}
   );
   gpc1_1 gpc1357 (
      {stage0_45[127]},
      {stage1_45[57]}
   );
   gpc1_1 gpc1358 (
      {stage0_46[96]},
      {stage1_46[48]}
   );
   gpc1_1 gpc1359 (
      {stage0_46[97]},
      {stage1_46[49]}
   );
   gpc1_1 gpc1360 (
      {stage0_46[98]},
      {stage1_46[50]}
   );
   gpc1_1 gpc1361 (
      {stage0_46[99]},
      {stage1_46[51]}
   );
   gpc1_1 gpc1362 (
      {stage0_46[100]},
      {stage1_46[52]}
   );
   gpc1_1 gpc1363 (
      {stage0_46[101]},
      {stage1_46[53]}
   );
   gpc1_1 gpc1364 (
      {stage0_46[102]},
      {stage1_46[54]}
   );
   gpc1_1 gpc1365 (
      {stage0_46[103]},
      {stage1_46[55]}
   );
   gpc1_1 gpc1366 (
      {stage0_46[104]},
      {stage1_46[56]}
   );
   gpc1_1 gpc1367 (
      {stage0_46[105]},
      {stage1_46[57]}
   );
   gpc1_1 gpc1368 (
      {stage0_46[106]},
      {stage1_46[58]}
   );
   gpc1_1 gpc1369 (
      {stage0_46[107]},
      {stage1_46[59]}
   );
   gpc1_1 gpc1370 (
      {stage0_46[108]},
      {stage1_46[60]}
   );
   gpc1_1 gpc1371 (
      {stage0_46[109]},
      {stage1_46[61]}
   );
   gpc1_1 gpc1372 (
      {stage0_46[110]},
      {stage1_46[62]}
   );
   gpc1_1 gpc1373 (
      {stage0_46[111]},
      {stage1_46[63]}
   );
   gpc1_1 gpc1374 (
      {stage0_46[112]},
      {stage1_46[64]}
   );
   gpc1_1 gpc1375 (
      {stage0_46[113]},
      {stage1_46[65]}
   );
   gpc1_1 gpc1376 (
      {stage0_46[114]},
      {stage1_46[66]}
   );
   gpc1_1 gpc1377 (
      {stage0_46[115]},
      {stage1_46[67]}
   );
   gpc1_1 gpc1378 (
      {stage0_46[116]},
      {stage1_46[68]}
   );
   gpc1_1 gpc1379 (
      {stage0_46[117]},
      {stage1_46[69]}
   );
   gpc1_1 gpc1380 (
      {stage0_46[118]},
      {stage1_46[70]}
   );
   gpc1_1 gpc1381 (
      {stage0_46[119]},
      {stage1_46[71]}
   );
   gpc1_1 gpc1382 (
      {stage0_46[120]},
      {stage1_46[72]}
   );
   gpc1_1 gpc1383 (
      {stage0_46[121]},
      {stage1_46[73]}
   );
   gpc1_1 gpc1384 (
      {stage0_46[122]},
      {stage1_46[74]}
   );
   gpc1_1 gpc1385 (
      {stage0_46[123]},
      {stage1_46[75]}
   );
   gpc1_1 gpc1386 (
      {stage0_46[124]},
      {stage1_46[76]}
   );
   gpc1_1 gpc1387 (
      {stage0_46[125]},
      {stage1_46[77]}
   );
   gpc1_1 gpc1388 (
      {stage0_46[126]},
      {stage1_46[78]}
   );
   gpc1_1 gpc1389 (
      {stage0_46[127]},
      {stage1_46[79]}
   );
   gpc1_1 gpc1390 (
      {stage0_47[103]},
      {stage1_47[45]}
   );
   gpc1_1 gpc1391 (
      {stage0_47[104]},
      {stage1_47[46]}
   );
   gpc1_1 gpc1392 (
      {stage0_47[105]},
      {stage1_47[47]}
   );
   gpc1_1 gpc1393 (
      {stage0_47[106]},
      {stage1_47[48]}
   );
   gpc1_1 gpc1394 (
      {stage0_47[107]},
      {stage1_47[49]}
   );
   gpc1_1 gpc1395 (
      {stage0_47[108]},
      {stage1_47[50]}
   );
   gpc1_1 gpc1396 (
      {stage0_47[109]},
      {stage1_47[51]}
   );
   gpc1_1 gpc1397 (
      {stage0_47[110]},
      {stage1_47[52]}
   );
   gpc1_1 gpc1398 (
      {stage0_47[111]},
      {stage1_47[53]}
   );
   gpc1_1 gpc1399 (
      {stage0_47[112]},
      {stage1_47[54]}
   );
   gpc1_1 gpc1400 (
      {stage0_47[113]},
      {stage1_47[55]}
   );
   gpc1_1 gpc1401 (
      {stage0_47[114]},
      {stage1_47[56]}
   );
   gpc1_1 gpc1402 (
      {stage0_47[115]},
      {stage1_47[57]}
   );
   gpc1_1 gpc1403 (
      {stage0_47[116]},
      {stage1_47[58]}
   );
   gpc1_1 gpc1404 (
      {stage0_47[117]},
      {stage1_47[59]}
   );
   gpc1_1 gpc1405 (
      {stage0_47[118]},
      {stage1_47[60]}
   );
   gpc1_1 gpc1406 (
      {stage0_47[119]},
      {stage1_47[61]}
   );
   gpc1_1 gpc1407 (
      {stage0_47[120]},
      {stage1_47[62]}
   );
   gpc1_1 gpc1408 (
      {stage0_47[121]},
      {stage1_47[63]}
   );
   gpc1_1 gpc1409 (
      {stage0_47[122]},
      {stage1_47[64]}
   );
   gpc1_1 gpc1410 (
      {stage0_47[123]},
      {stage1_47[65]}
   );
   gpc1_1 gpc1411 (
      {stage0_47[124]},
      {stage1_47[66]}
   );
   gpc1_1 gpc1412 (
      {stage0_47[125]},
      {stage1_47[67]}
   );
   gpc1_1 gpc1413 (
      {stage0_47[126]},
      {stage1_47[68]}
   );
   gpc1_1 gpc1414 (
      {stage0_47[127]},
      {stage1_47[69]}
   );
   gpc1_1 gpc1415 (
      {stage0_48[127]},
      {stage1_48[45]}
   );
   gpc1_1 gpc1416 (
      {stage0_50[106]},
      {stage1_50[49]}
   );
   gpc1_1 gpc1417 (
      {stage0_50[107]},
      {stage1_50[50]}
   );
   gpc1_1 gpc1418 (
      {stage0_50[108]},
      {stage1_50[51]}
   );
   gpc1_1 gpc1419 (
      {stage0_50[109]},
      {stage1_50[52]}
   );
   gpc1_1 gpc1420 (
      {stage0_50[110]},
      {stage1_50[53]}
   );
   gpc1_1 gpc1421 (
      {stage0_50[111]},
      {stage1_50[54]}
   );
   gpc1_1 gpc1422 (
      {stage0_50[112]},
      {stage1_50[55]}
   );
   gpc1_1 gpc1423 (
      {stage0_50[113]},
      {stage1_50[56]}
   );
   gpc1_1 gpc1424 (
      {stage0_50[114]},
      {stage1_50[57]}
   );
   gpc1_1 gpc1425 (
      {stage0_50[115]},
      {stage1_50[58]}
   );
   gpc1_1 gpc1426 (
      {stage0_50[116]},
      {stage1_50[59]}
   );
   gpc1_1 gpc1427 (
      {stage0_50[117]},
      {stage1_50[60]}
   );
   gpc1_1 gpc1428 (
      {stage0_50[118]},
      {stage1_50[61]}
   );
   gpc1_1 gpc1429 (
      {stage0_50[119]},
      {stage1_50[62]}
   );
   gpc1_1 gpc1430 (
      {stage0_50[120]},
      {stage1_50[63]}
   );
   gpc1_1 gpc1431 (
      {stage0_50[121]},
      {stage1_50[64]}
   );
   gpc1_1 gpc1432 (
      {stage0_50[122]},
      {stage1_50[65]}
   );
   gpc1_1 gpc1433 (
      {stage0_50[123]},
      {stage1_50[66]}
   );
   gpc1_1 gpc1434 (
      {stage0_50[124]},
      {stage1_50[67]}
   );
   gpc1_1 gpc1435 (
      {stage0_50[125]},
      {stage1_50[68]}
   );
   gpc1_1 gpc1436 (
      {stage0_50[126]},
      {stage1_50[69]}
   );
   gpc1_1 gpc1437 (
      {stage0_50[127]},
      {stage1_50[70]}
   );
   gpc1_1 gpc1438 (
      {stage0_52[120]},
      {stage1_52[53]}
   );
   gpc1_1 gpc1439 (
      {stage0_52[121]},
      {stage1_52[54]}
   );
   gpc1_1 gpc1440 (
      {stage0_52[122]},
      {stage1_52[55]}
   );
   gpc1_1 gpc1441 (
      {stage0_52[123]},
      {stage1_52[56]}
   );
   gpc1_1 gpc1442 (
      {stage0_52[124]},
      {stage1_52[57]}
   );
   gpc1_1 gpc1443 (
      {stage0_52[125]},
      {stage1_52[58]}
   );
   gpc1_1 gpc1444 (
      {stage0_52[126]},
      {stage1_52[59]}
   );
   gpc1_1 gpc1445 (
      {stage0_52[127]},
      {stage1_52[60]}
   );
   gpc1_1 gpc1446 (
      {stage0_53[120]},
      {stage1_53[54]}
   );
   gpc1_1 gpc1447 (
      {stage0_53[121]},
      {stage1_53[55]}
   );
   gpc1_1 gpc1448 (
      {stage0_53[122]},
      {stage1_53[56]}
   );
   gpc1_1 gpc1449 (
      {stage0_53[123]},
      {stage1_53[57]}
   );
   gpc1_1 gpc1450 (
      {stage0_53[124]},
      {stage1_53[58]}
   );
   gpc1_1 gpc1451 (
      {stage0_53[125]},
      {stage1_53[59]}
   );
   gpc1_1 gpc1452 (
      {stage0_53[126]},
      {stage1_53[60]}
   );
   gpc1_1 gpc1453 (
      {stage0_53[127]},
      {stage1_53[61]}
   );
   gpc1_1 gpc1454 (
      {stage0_54[123]},
      {stage1_54[47]}
   );
   gpc1_1 gpc1455 (
      {stage0_54[124]},
      {stage1_54[48]}
   );
   gpc1_1 gpc1456 (
      {stage0_54[125]},
      {stage1_54[49]}
   );
   gpc1_1 gpc1457 (
      {stage0_54[126]},
      {stage1_54[50]}
   );
   gpc1_1 gpc1458 (
      {stage0_54[127]},
      {stage1_54[51]}
   );
   gpc1_1 gpc1459 (
      {stage0_55[108]},
      {stage1_55[48]}
   );
   gpc1_1 gpc1460 (
      {stage0_55[109]},
      {stage1_55[49]}
   );
   gpc1_1 gpc1461 (
      {stage0_55[110]},
      {stage1_55[50]}
   );
   gpc1_1 gpc1462 (
      {stage0_55[111]},
      {stage1_55[51]}
   );
   gpc1_1 gpc1463 (
      {stage0_55[112]},
      {stage1_55[52]}
   );
   gpc1_1 gpc1464 (
      {stage0_55[113]},
      {stage1_55[53]}
   );
   gpc1_1 gpc1465 (
      {stage0_55[114]},
      {stage1_55[54]}
   );
   gpc1_1 gpc1466 (
      {stage0_55[115]},
      {stage1_55[55]}
   );
   gpc1_1 gpc1467 (
      {stage0_55[116]},
      {stage1_55[56]}
   );
   gpc1_1 gpc1468 (
      {stage0_55[117]},
      {stage1_55[57]}
   );
   gpc1_1 gpc1469 (
      {stage0_55[118]},
      {stage1_55[58]}
   );
   gpc1_1 gpc1470 (
      {stage0_55[119]},
      {stage1_55[59]}
   );
   gpc1_1 gpc1471 (
      {stage0_55[120]},
      {stage1_55[60]}
   );
   gpc1_1 gpc1472 (
      {stage0_55[121]},
      {stage1_55[61]}
   );
   gpc1_1 gpc1473 (
      {stage0_55[122]},
      {stage1_55[62]}
   );
   gpc1_1 gpc1474 (
      {stage0_55[123]},
      {stage1_55[63]}
   );
   gpc1_1 gpc1475 (
      {stage0_55[124]},
      {stage1_55[64]}
   );
   gpc1_1 gpc1476 (
      {stage0_55[125]},
      {stage1_55[65]}
   );
   gpc1_1 gpc1477 (
      {stage0_55[126]},
      {stage1_55[66]}
   );
   gpc1_1 gpc1478 (
      {stage0_55[127]},
      {stage1_55[67]}
   );
   gpc1_1 gpc1479 (
      {stage0_56[122]},
      {stage1_56[51]}
   );
   gpc1_1 gpc1480 (
      {stage0_56[123]},
      {stage1_56[52]}
   );
   gpc1_1 gpc1481 (
      {stage0_56[124]},
      {stage1_56[53]}
   );
   gpc1_1 gpc1482 (
      {stage0_56[125]},
      {stage1_56[54]}
   );
   gpc1_1 gpc1483 (
      {stage0_56[126]},
      {stage1_56[55]}
   );
   gpc1_1 gpc1484 (
      {stage0_56[127]},
      {stage1_56[56]}
   );
   gpc1_1 gpc1485 (
      {stage0_57[122]},
      {stage1_57[52]}
   );
   gpc1_1 gpc1486 (
      {stage0_57[123]},
      {stage1_57[53]}
   );
   gpc1_1 gpc1487 (
      {stage0_57[124]},
      {stage1_57[54]}
   );
   gpc1_1 gpc1488 (
      {stage0_57[125]},
      {stage1_57[55]}
   );
   gpc1_1 gpc1489 (
      {stage0_57[126]},
      {stage1_57[56]}
   );
   gpc1_1 gpc1490 (
      {stage0_57[127]},
      {stage1_57[57]}
   );
   gpc1_1 gpc1491 (
      {stage0_58[117]},
      {stage1_58[49]}
   );
   gpc1_1 gpc1492 (
      {stage0_58[118]},
      {stage1_58[50]}
   );
   gpc1_1 gpc1493 (
      {stage0_58[119]},
      {stage1_58[51]}
   );
   gpc1_1 gpc1494 (
      {stage0_58[120]},
      {stage1_58[52]}
   );
   gpc1_1 gpc1495 (
      {stage0_58[121]},
      {stage1_58[53]}
   );
   gpc1_1 gpc1496 (
      {stage0_58[122]},
      {stage1_58[54]}
   );
   gpc1_1 gpc1497 (
      {stage0_58[123]},
      {stage1_58[55]}
   );
   gpc1_1 gpc1498 (
      {stage0_58[124]},
      {stage1_58[56]}
   );
   gpc1_1 gpc1499 (
      {stage0_58[125]},
      {stage1_58[57]}
   );
   gpc1_1 gpc1500 (
      {stage0_58[126]},
      {stage1_58[58]}
   );
   gpc1_1 gpc1501 (
      {stage0_58[127]},
      {stage1_58[59]}
   );
   gpc1_1 gpc1502 (
      {stage0_59[118]},
      {stage1_59[46]}
   );
   gpc1_1 gpc1503 (
      {stage0_59[119]},
      {stage1_59[47]}
   );
   gpc1_1 gpc1504 (
      {stage0_59[120]},
      {stage1_59[48]}
   );
   gpc1_1 gpc1505 (
      {stage0_59[121]},
      {stage1_59[49]}
   );
   gpc1_1 gpc1506 (
      {stage0_59[122]},
      {stage1_59[50]}
   );
   gpc1_1 gpc1507 (
      {stage0_59[123]},
      {stage1_59[51]}
   );
   gpc1_1 gpc1508 (
      {stage0_59[124]},
      {stage1_59[52]}
   );
   gpc1_1 gpc1509 (
      {stage0_59[125]},
      {stage1_59[53]}
   );
   gpc1_1 gpc1510 (
      {stage0_59[126]},
      {stage1_59[54]}
   );
   gpc1_1 gpc1511 (
      {stage0_59[127]},
      {stage1_59[55]}
   );
   gpc1_1 gpc1512 (
      {stage0_60[126]},
      {stage1_60[51]}
   );
   gpc1_1 gpc1513 (
      {stage0_60[127]},
      {stage1_60[52]}
   );
   gpc1_1 gpc1514 (
      {stage0_61[126]},
      {stage1_61[57]}
   );
   gpc1_1 gpc1515 (
      {stage0_61[127]},
      {stage1_61[58]}
   );
   gpc1_1 gpc1516 (
      {stage0_62[72]},
      {stage1_62[42]}
   );
   gpc1_1 gpc1517 (
      {stage0_62[73]},
      {stage1_62[43]}
   );
   gpc1_1 gpc1518 (
      {stage0_62[74]},
      {stage1_62[44]}
   );
   gpc1_1 gpc1519 (
      {stage0_62[75]},
      {stage1_62[45]}
   );
   gpc1_1 gpc1520 (
      {stage0_62[76]},
      {stage1_62[46]}
   );
   gpc1_1 gpc1521 (
      {stage0_62[77]},
      {stage1_62[47]}
   );
   gpc1_1 gpc1522 (
      {stage0_62[78]},
      {stage1_62[48]}
   );
   gpc1_1 gpc1523 (
      {stage0_62[79]},
      {stage1_62[49]}
   );
   gpc1_1 gpc1524 (
      {stage0_62[80]},
      {stage1_62[50]}
   );
   gpc1_1 gpc1525 (
      {stage0_62[81]},
      {stage1_62[51]}
   );
   gpc1_1 gpc1526 (
      {stage0_62[82]},
      {stage1_62[52]}
   );
   gpc1_1 gpc1527 (
      {stage0_62[83]},
      {stage1_62[53]}
   );
   gpc1_1 gpc1528 (
      {stage0_62[84]},
      {stage1_62[54]}
   );
   gpc1_1 gpc1529 (
      {stage0_62[85]},
      {stage1_62[55]}
   );
   gpc1_1 gpc1530 (
      {stage0_62[86]},
      {stage1_62[56]}
   );
   gpc1_1 gpc1531 (
      {stage0_62[87]},
      {stage1_62[57]}
   );
   gpc1_1 gpc1532 (
      {stage0_62[88]},
      {stage1_62[58]}
   );
   gpc1_1 gpc1533 (
      {stage0_62[89]},
      {stage1_62[59]}
   );
   gpc1_1 gpc1534 (
      {stage0_62[90]},
      {stage1_62[60]}
   );
   gpc1_1 gpc1535 (
      {stage0_62[91]},
      {stage1_62[61]}
   );
   gpc1_1 gpc1536 (
      {stage0_62[92]},
      {stage1_62[62]}
   );
   gpc1_1 gpc1537 (
      {stage0_62[93]},
      {stage1_62[63]}
   );
   gpc1_1 gpc1538 (
      {stage0_62[94]},
      {stage1_62[64]}
   );
   gpc1_1 gpc1539 (
      {stage0_62[95]},
      {stage1_62[65]}
   );
   gpc1_1 gpc1540 (
      {stage0_62[96]},
      {stage1_62[66]}
   );
   gpc1_1 gpc1541 (
      {stage0_62[97]},
      {stage1_62[67]}
   );
   gpc1_1 gpc1542 (
      {stage0_62[98]},
      {stage1_62[68]}
   );
   gpc1_1 gpc1543 (
      {stage0_62[99]},
      {stage1_62[69]}
   );
   gpc1_1 gpc1544 (
      {stage0_62[100]},
      {stage1_62[70]}
   );
   gpc1_1 gpc1545 (
      {stage0_62[101]},
      {stage1_62[71]}
   );
   gpc1_1 gpc1546 (
      {stage0_62[102]},
      {stage1_62[72]}
   );
   gpc1_1 gpc1547 (
      {stage0_62[103]},
      {stage1_62[73]}
   );
   gpc1_1 gpc1548 (
      {stage0_62[104]},
      {stage1_62[74]}
   );
   gpc1_1 gpc1549 (
      {stage0_62[105]},
      {stage1_62[75]}
   );
   gpc1_1 gpc1550 (
      {stage0_62[106]},
      {stage1_62[76]}
   );
   gpc1_1 gpc1551 (
      {stage0_62[107]},
      {stage1_62[77]}
   );
   gpc1_1 gpc1552 (
      {stage0_62[108]},
      {stage1_62[78]}
   );
   gpc1_1 gpc1553 (
      {stage0_62[109]},
      {stage1_62[79]}
   );
   gpc1_1 gpc1554 (
      {stage0_62[110]},
      {stage1_62[80]}
   );
   gpc1_1 gpc1555 (
      {stage0_62[111]},
      {stage1_62[81]}
   );
   gpc1_1 gpc1556 (
      {stage0_62[112]},
      {stage1_62[82]}
   );
   gpc1_1 gpc1557 (
      {stage0_62[113]},
      {stage1_62[83]}
   );
   gpc1_1 gpc1558 (
      {stage0_62[114]},
      {stage1_62[84]}
   );
   gpc1_1 gpc1559 (
      {stage0_62[115]},
      {stage1_62[85]}
   );
   gpc1_1 gpc1560 (
      {stage0_62[116]},
      {stage1_62[86]}
   );
   gpc1_1 gpc1561 (
      {stage0_62[117]},
      {stage1_62[87]}
   );
   gpc1_1 gpc1562 (
      {stage0_62[118]},
      {stage1_62[88]}
   );
   gpc1_1 gpc1563 (
      {stage0_62[119]},
      {stage1_62[89]}
   );
   gpc1_1 gpc1564 (
      {stage0_62[120]},
      {stage1_62[90]}
   );
   gpc1_1 gpc1565 (
      {stage0_62[121]},
      {stage1_62[91]}
   );
   gpc1_1 gpc1566 (
      {stage0_62[122]},
      {stage1_62[92]}
   );
   gpc1_1 gpc1567 (
      {stage0_62[123]},
      {stage1_62[93]}
   );
   gpc1_1 gpc1568 (
      {stage0_62[124]},
      {stage1_62[94]}
   );
   gpc1_1 gpc1569 (
      {stage0_62[125]},
      {stage1_62[95]}
   );
   gpc1_1 gpc1570 (
      {stage0_62[126]},
      {stage1_62[96]}
   );
   gpc1_1 gpc1571 (
      {stage0_62[127]},
      {stage1_62[97]}
   );
   gpc1_1 gpc1572 (
      {stage0_63[108]},
      {stage1_63[33]}
   );
   gpc1_1 gpc1573 (
      {stage0_63[109]},
      {stage1_63[34]}
   );
   gpc1_1 gpc1574 (
      {stage0_63[110]},
      {stage1_63[35]}
   );
   gpc1_1 gpc1575 (
      {stage0_63[111]},
      {stage1_63[36]}
   );
   gpc1_1 gpc1576 (
      {stage0_63[112]},
      {stage1_63[37]}
   );
   gpc1_1 gpc1577 (
      {stage0_63[113]},
      {stage1_63[38]}
   );
   gpc1_1 gpc1578 (
      {stage0_63[114]},
      {stage1_63[39]}
   );
   gpc1_1 gpc1579 (
      {stage0_63[115]},
      {stage1_63[40]}
   );
   gpc1_1 gpc1580 (
      {stage0_63[116]},
      {stage1_63[41]}
   );
   gpc1_1 gpc1581 (
      {stage0_63[117]},
      {stage1_63[42]}
   );
   gpc1_1 gpc1582 (
      {stage0_63[118]},
      {stage1_63[43]}
   );
   gpc1_1 gpc1583 (
      {stage0_63[119]},
      {stage1_63[44]}
   );
   gpc1_1 gpc1584 (
      {stage0_63[120]},
      {stage1_63[45]}
   );
   gpc1_1 gpc1585 (
      {stage0_63[121]},
      {stage1_63[46]}
   );
   gpc1_1 gpc1586 (
      {stage0_63[122]},
      {stage1_63[47]}
   );
   gpc1_1 gpc1587 (
      {stage0_63[123]},
      {stage1_63[48]}
   );
   gpc1_1 gpc1588 (
      {stage0_63[124]},
      {stage1_63[49]}
   );
   gpc1_1 gpc1589 (
      {stage0_63[125]},
      {stage1_63[50]}
   );
   gpc1_1 gpc1590 (
      {stage0_63[126]},
      {stage1_63[51]}
   );
   gpc1_1 gpc1591 (
      {stage0_63[127]},
      {stage1_63[52]}
   );
   gpc1163_5 gpc1592 (
      {stage1_0[0], stage1_0[1], stage1_0[2]},
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_2[0]},
      {stage1_3[0]},
      {stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0],stage2_0[0]}
   );
   gpc615_5 gpc1593 (
      {stage1_0[3], stage1_0[4], stage1_0[5], stage1_0[6], stage1_0[7]},
      {stage1_1[6]},
      {stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5], stage1_2[6]},
      {stage2_4[1],stage2_3[1],stage2_2[1],stage2_1[1],stage2_0[1]}
   );
   gpc615_5 gpc1594 (
      {stage1_0[8], stage1_0[9], stage1_0[10], stage1_0[11], stage1_0[12]},
      {stage1_1[7]},
      {stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10], stage1_2[11], stage1_2[12]},
      {stage2_4[2],stage2_3[2],stage2_2[2],stage2_1[2],stage2_0[2]}
   );
   gpc606_5 gpc1595 (
      {stage1_1[8], stage1_1[9], stage1_1[10], stage1_1[11], stage1_1[12], stage1_1[13]},
      {stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5], stage1_3[6]},
      {stage2_5[0],stage2_4[3],stage2_3[3],stage2_2[3],stage2_1[3]}
   );
   gpc606_5 gpc1596 (
      {stage1_1[14], stage1_1[15], stage1_1[16], stage1_1[17], stage1_1[18], stage1_1[19]},
      {stage1_3[7], stage1_3[8], stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12]},
      {stage2_5[1],stage2_4[4],stage2_3[4],stage2_2[4],stage2_1[4]}
   );
   gpc606_5 gpc1597 (
      {stage1_1[20], stage1_1[21], stage1_1[22], stage1_1[23], stage1_1[24], stage1_1[25]},
      {stage1_3[13], stage1_3[14], stage1_3[15], stage1_3[16], stage1_3[17], stage1_3[18]},
      {stage2_5[2],stage2_4[5],stage2_3[5],stage2_2[5],stage2_1[5]}
   );
   gpc606_5 gpc1598 (
      {stage1_2[13], stage1_2[14], stage1_2[15], stage1_2[16], stage1_2[17], stage1_2[18]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[3],stage2_4[6],stage2_3[6],stage2_2[6]}
   );
   gpc606_5 gpc1599 (
      {stage1_2[19], stage1_2[20], stage1_2[21], stage1_2[22], stage1_2[23], stage1_2[24]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[4],stage2_4[7],stage2_3[7],stage2_2[7]}
   );
   gpc606_5 gpc1600 (
      {stage1_2[25], stage1_2[26], stage1_2[27], stage1_2[28], stage1_2[29], stage1_2[30]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[5],stage2_4[8],stage2_3[8],stage2_2[8]}
   );
   gpc1163_5 gpc1601 (
      {stage1_3[19], stage1_3[20], stage1_3[21]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage1_5[0]},
      {stage1_6[0]},
      {stage2_7[0],stage2_6[3],stage2_5[6],stage2_4[9],stage2_3[9]}
   );
   gpc606_5 gpc1602 (
      {stage1_3[22], stage1_3[23], stage1_3[24], stage1_3[25], stage1_3[26], stage1_3[27]},
      {stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5], stage1_5[6]},
      {stage2_7[1],stage2_6[4],stage2_5[7],stage2_4[10],stage2_3[10]}
   );
   gpc606_5 gpc1603 (
      {stage1_3[28], stage1_3[29], stage1_3[30], stage1_3[31], stage1_3[32], stage1_3[33]},
      {stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11], stage1_5[12]},
      {stage2_7[2],stage2_6[5],stage2_5[8],stage2_4[11],stage2_3[11]}
   );
   gpc606_5 gpc1604 (
      {stage1_3[34], stage1_3[35], stage1_3[36], stage1_3[37], stage1_3[38], stage1_3[39]},
      {stage1_5[13], stage1_5[14], stage1_5[15], stage1_5[16], stage1_5[17], stage1_5[18]},
      {stage2_7[3],stage2_6[6],stage2_5[9],stage2_4[12],stage2_3[12]}
   );
   gpc615_5 gpc1605 (
      {stage1_3[40], stage1_3[41], stage1_3[42], stage1_3[43], stage1_3[44]},
      {stage1_4[24]},
      {stage1_5[19], stage1_5[20], stage1_5[21], stage1_5[22], stage1_5[23], stage1_5[24]},
      {stage2_7[4],stage2_6[7],stage2_5[10],stage2_4[13],stage2_3[13]}
   );
   gpc615_5 gpc1606 (
      {stage1_3[45], stage1_3[46], stage1_3[47], stage1_3[48], stage1_3[49]},
      {stage1_4[25]},
      {stage1_5[25], stage1_5[26], stage1_5[27], stage1_5[28], stage1_5[29], stage1_5[30]},
      {stage2_7[5],stage2_6[8],stage2_5[11],stage2_4[14],stage2_3[14]}
   );
   gpc615_5 gpc1607 (
      {stage1_3[50], stage1_3[51], stage1_3[52], stage1_3[53], stage1_3[54]},
      {stage1_4[26]},
      {stage1_5[31], stage1_5[32], stage1_5[33], stage1_5[34], stage1_5[35], stage1_5[36]},
      {stage2_7[6],stage2_6[9],stage2_5[12],stage2_4[15],stage2_3[15]}
   );
   gpc606_5 gpc1608 (
      {stage1_4[27], stage1_4[28], stage1_4[29], stage1_4[30], stage1_4[31], stage1_4[32]},
      {stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5], stage1_6[6]},
      {stage2_8[0],stage2_7[7],stage2_6[10],stage2_5[13],stage2_4[16]}
   );
   gpc615_5 gpc1609 (
      {stage1_4[33], stage1_4[34], stage1_4[35], stage1_4[36], stage1_4[37]},
      {stage1_5[37]},
      {stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10], stage1_6[11], stage1_6[12]},
      {stage2_8[1],stage2_7[8],stage2_6[11],stage2_5[14],stage2_4[17]}
   );
   gpc615_5 gpc1610 (
      {stage1_4[38], stage1_4[39], stage1_4[40], stage1_4[41], stage1_4[42]},
      {stage1_5[38]},
      {stage1_6[13], stage1_6[14], stage1_6[15], stage1_6[16], stage1_6[17], stage1_6[18]},
      {stage2_8[2],stage2_7[9],stage2_6[12],stage2_5[15],stage2_4[18]}
   );
   gpc615_5 gpc1611 (
      {stage1_4[43], stage1_4[44], stage1_4[45], stage1_4[46], stage1_4[47]},
      {stage1_5[39]},
      {stage1_6[19], stage1_6[20], stage1_6[21], stage1_6[22], stage1_6[23], stage1_6[24]},
      {stage2_8[3],stage2_7[10],stage2_6[13],stage2_5[16],stage2_4[19]}
   );
   gpc615_5 gpc1612 (
      {stage1_4[48], stage1_4[49], stage1_4[50], stage1_4[51], stage1_4[52]},
      {stage1_5[40]},
      {stage1_6[25], stage1_6[26], stage1_6[27], stage1_6[28], stage1_6[29], stage1_6[30]},
      {stage2_8[4],stage2_7[11],stage2_6[14],stage2_5[17],stage2_4[20]}
   );
   gpc615_5 gpc1613 (
      {stage1_4[53], stage1_4[54], stage1_4[55], stage1_4[56], stage1_4[57]},
      {stage1_5[41]},
      {stage1_6[31], stage1_6[32], stage1_6[33], stage1_6[34], stage1_6[35], stage1_6[36]},
      {stage2_8[5],stage2_7[12],stage2_6[15],stage2_5[18],stage2_4[21]}
   );
   gpc615_5 gpc1614 (
      {stage1_4[58], stage1_4[59], stage1_4[60], stage1_4[61], stage1_4[62]},
      {stage1_5[42]},
      {stage1_6[37], stage1_6[38], stage1_6[39], stage1_6[40], stage1_6[41], stage1_6[42]},
      {stage2_8[6],stage2_7[13],stage2_6[16],stage2_5[19],stage2_4[22]}
   );
   gpc606_5 gpc1615 (
      {stage1_6[43], stage1_6[44], stage1_6[45], stage1_6[46], stage1_6[47], stage1_6[48]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[0],stage2_8[7],stage2_7[14],stage2_6[17]}
   );
   gpc606_5 gpc1616 (
      {stage1_6[49], stage1_6[50], stage1_6[51], stage1_6[52], stage1_6[53], stage1_6[54]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[1],stage2_8[8],stage2_7[15],stage2_6[18]}
   );
   gpc615_5 gpc1617 (
      {stage1_6[55], stage1_6[56], stage1_6[57], stage1_6[58], stage1_6[59]},
      {stage1_7[0]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[2],stage2_8[9],stage2_7[16],stage2_6[19]}
   );
   gpc615_5 gpc1618 (
      {stage1_6[60], stage1_6[61], stage1_6[62], stage1_6[63], stage1_6[64]},
      {stage1_7[1]},
      {stage1_8[18], stage1_8[19], stage1_8[20], stage1_8[21], stage1_8[22], stage1_8[23]},
      {stage2_10[3],stage2_9[3],stage2_8[10],stage2_7[17],stage2_6[20]}
   );
   gpc615_5 gpc1619 (
      {stage1_6[65], stage1_6[66], stage1_6[67], stage1_6[68], stage1_6[69]},
      {stage1_7[2]},
      {stage1_8[24], stage1_8[25], stage1_8[26], stage1_8[27], stage1_8[28], stage1_8[29]},
      {stage2_10[4],stage2_9[4],stage2_8[11],stage2_7[18],stage2_6[21]}
   );
   gpc615_5 gpc1620 (
      {stage1_6[70], stage1_6[71], stage1_6[72], stage1_6[73], stage1_6[74]},
      {stage1_7[3]},
      {stage1_8[30], stage1_8[31], stage1_8[32], stage1_8[33], stage1_8[34], stage1_8[35]},
      {stage2_10[5],stage2_9[5],stage2_8[12],stage2_7[19],stage2_6[22]}
   );
   gpc615_5 gpc1621 (
      {stage1_6[75], stage1_6[76], stage1_6[77], stage1_6[78], stage1_6[79]},
      {stage1_7[4]},
      {stage1_8[36], stage1_8[37], stage1_8[38], stage1_8[39], stage1_8[40], stage1_8[41]},
      {stage2_10[6],stage2_9[6],stage2_8[13],stage2_7[20],stage2_6[23]}
   );
   gpc615_5 gpc1622 (
      {stage1_6[80], stage1_6[81], stage1_6[82], stage1_6[83], stage1_6[84]},
      {stage1_7[5]},
      {stage1_8[42], stage1_8[43], stage1_8[44], stage1_8[45], stage1_8[46], stage1_8[47]},
      {stage2_10[7],stage2_9[7],stage2_8[14],stage2_7[21],stage2_6[24]}
   );
   gpc615_5 gpc1623 (
      {stage1_6[85], stage1_6[86], stage1_6[87], stage1_6[88], 1'b0},
      {stage1_7[6]},
      {stage1_8[48], stage1_8[49], stage1_8[50], stage1_8[51], stage1_8[52], stage1_8[53]},
      {stage2_10[8],stage2_9[8],stage2_8[15],stage2_7[22],stage2_6[25]}
   );
   gpc1406_5 gpc1624 (
      {stage1_7[7], stage1_7[8], stage1_7[9], stage1_7[10], stage1_7[11], stage1_7[12]},
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3]},
      {stage1_10[0]},
      {stage2_11[0],stage2_10[9],stage2_9[9],stage2_8[16],stage2_7[23]}
   );
   gpc117_4 gpc1625 (
      {stage1_7[13], stage1_7[14], stage1_7[15], stage1_7[16], stage1_7[17], stage1_7[18], stage1_7[19]},
      {stage1_8[54]},
      {stage1_9[4]},
      {stage2_10[10],stage2_9[10],stage2_8[17],stage2_7[24]}
   );
   gpc117_4 gpc1626 (
      {stage1_7[20], stage1_7[21], stage1_7[22], stage1_7[23], stage1_7[24], stage1_7[25], stage1_7[26]},
      {stage1_8[55]},
      {stage1_9[5]},
      {stage2_10[11],stage2_9[11],stage2_8[18],stage2_7[25]}
   );
   gpc117_4 gpc1627 (
      {stage1_7[27], stage1_7[28], stage1_7[29], stage1_7[30], stage1_7[31], stage1_7[32], stage1_7[33]},
      {stage1_8[56]},
      {stage1_9[6]},
      {stage2_10[12],stage2_9[12],stage2_8[19],stage2_7[26]}
   );
   gpc117_4 gpc1628 (
      {stage1_7[34], stage1_7[35], stage1_7[36], stage1_7[37], stage1_7[38], stage1_7[39], stage1_7[40]},
      {stage1_8[57]},
      {stage1_9[7]},
      {stage2_10[13],stage2_9[13],stage2_8[20],stage2_7[27]}
   );
   gpc606_5 gpc1629 (
      {stage1_7[41], stage1_7[42], stage1_7[43], stage1_7[44], stage1_7[45], stage1_7[46]},
      {stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11], stage1_9[12], stage1_9[13]},
      {stage2_11[1],stage2_10[14],stage2_9[14],stage2_8[21],stage2_7[28]}
   );
   gpc606_5 gpc1630 (
      {stage1_7[47], stage1_7[48], stage1_7[49], stage1_7[50], stage1_7[51], stage1_7[52]},
      {stage1_9[14], stage1_9[15], stage1_9[16], stage1_9[17], stage1_9[18], stage1_9[19]},
      {stage2_11[2],stage2_10[15],stage2_9[15],stage2_8[22],stage2_7[29]}
   );
   gpc606_5 gpc1631 (
      {stage1_7[53], stage1_7[54], stage1_7[55], stage1_7[56], stage1_7[57], stage1_7[58]},
      {stage1_9[20], stage1_9[21], stage1_9[22], stage1_9[23], stage1_9[24], stage1_9[25]},
      {stage2_11[3],stage2_10[16],stage2_9[16],stage2_8[23],stage2_7[30]}
   );
   gpc615_5 gpc1632 (
      {stage1_7[59], stage1_7[60], stage1_7[61], stage1_7[62], stage1_7[63]},
      {stage1_8[58]},
      {stage1_9[26], stage1_9[27], stage1_9[28], stage1_9[29], stage1_9[30], stage1_9[31]},
      {stage2_11[4],stage2_10[17],stage2_9[17],stage2_8[24],stage2_7[31]}
   );
   gpc606_5 gpc1633 (
      {stage1_9[32], stage1_9[33], stage1_9[34], stage1_9[35], stage1_9[36], stage1_9[37]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[0],stage2_11[5],stage2_10[18],stage2_9[18]}
   );
   gpc615_5 gpc1634 (
      {stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage1_11[6]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[1],stage2_12[1],stage2_11[6],stage2_10[19]}
   );
   gpc615_5 gpc1635 (
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10]},
      {stage1_11[7]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[2],stage2_12[2],stage2_11[7],stage2_10[20]}
   );
   gpc615_5 gpc1636 (
      {stage1_10[11], stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15]},
      {stage1_11[8]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[3],stage2_12[3],stage2_11[8],stage2_10[21]}
   );
   gpc615_5 gpc1637 (
      {stage1_10[16], stage1_10[17], stage1_10[18], stage1_10[19], stage1_10[20]},
      {stage1_11[9]},
      {stage1_12[18], stage1_12[19], stage1_12[20], stage1_12[21], stage1_12[22], stage1_12[23]},
      {stage2_14[3],stage2_13[4],stage2_12[4],stage2_11[9],stage2_10[22]}
   );
   gpc615_5 gpc1638 (
      {stage1_10[21], stage1_10[22], stage1_10[23], stage1_10[24], stage1_10[25]},
      {stage1_11[10]},
      {stage1_12[24], stage1_12[25], stage1_12[26], stage1_12[27], stage1_12[28], stage1_12[29]},
      {stage2_14[4],stage2_13[5],stage2_12[5],stage2_11[10],stage2_10[23]}
   );
   gpc615_5 gpc1639 (
      {stage1_10[26], stage1_10[27], stage1_10[28], stage1_10[29], stage1_10[30]},
      {stage1_11[11]},
      {stage1_12[30], stage1_12[31], stage1_12[32], stage1_12[33], stage1_12[34], stage1_12[35]},
      {stage2_14[5],stage2_13[6],stage2_12[6],stage2_11[11],stage2_10[24]}
   );
   gpc615_5 gpc1640 (
      {stage1_10[31], stage1_10[32], stage1_10[33], stage1_10[34], stage1_10[35]},
      {stage1_11[12]},
      {stage1_12[36], stage1_12[37], stage1_12[38], stage1_12[39], stage1_12[40], stage1_12[41]},
      {stage2_14[6],stage2_13[7],stage2_12[7],stage2_11[12],stage2_10[25]}
   );
   gpc606_5 gpc1641 (
      {stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16], stage1_11[17], stage1_11[18]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[7],stage2_13[8],stage2_12[8],stage2_11[13]}
   );
   gpc606_5 gpc1642 (
      {stage1_11[19], stage1_11[20], stage1_11[21], stage1_11[22], stage1_11[23], stage1_11[24]},
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage2_15[1],stage2_14[8],stage2_13[9],stage2_12[9],stage2_11[14]}
   );
   gpc606_5 gpc1643 (
      {stage1_11[25], stage1_11[26], stage1_11[27], stage1_11[28], stage1_11[29], stage1_11[30]},
      {stage1_13[12], stage1_13[13], stage1_13[14], stage1_13[15], stage1_13[16], stage1_13[17]},
      {stage2_15[2],stage2_14[9],stage2_13[10],stage2_12[10],stage2_11[15]}
   );
   gpc606_5 gpc1644 (
      {stage1_11[31], stage1_11[32], stage1_11[33], stage1_11[34], stage1_11[35], stage1_11[36]},
      {stage1_13[18], stage1_13[19], stage1_13[20], stage1_13[21], stage1_13[22], stage1_13[23]},
      {stage2_15[3],stage2_14[10],stage2_13[11],stage2_12[11],stage2_11[16]}
   );
   gpc606_5 gpc1645 (
      {stage1_11[37], stage1_11[38], stage1_11[39], stage1_11[40], stage1_11[41], stage1_11[42]},
      {stage1_13[24], stage1_13[25], stage1_13[26], stage1_13[27], stage1_13[28], stage1_13[29]},
      {stage2_15[4],stage2_14[11],stage2_13[12],stage2_12[12],stage2_11[17]}
   );
   gpc606_5 gpc1646 (
      {stage1_11[43], stage1_11[44], stage1_11[45], stage1_11[46], stage1_11[47], stage1_11[48]},
      {stage1_13[30], stage1_13[31], stage1_13[32], stage1_13[33], stage1_13[34], stage1_13[35]},
      {stage2_15[5],stage2_14[12],stage2_13[13],stage2_12[13],stage2_11[18]}
   );
   gpc615_5 gpc1647 (
      {stage1_11[49], stage1_11[50], stage1_11[51], stage1_11[52], stage1_11[53]},
      {stage1_12[42]},
      {stage1_13[36], stage1_13[37], stage1_13[38], stage1_13[39], stage1_13[40], stage1_13[41]},
      {stage2_15[6],stage2_14[13],stage2_13[14],stage2_12[14],stage2_11[19]}
   );
   gpc615_5 gpc1648 (
      {stage1_11[54], stage1_11[55], stage1_11[56], stage1_11[57], stage1_11[58]},
      {stage1_12[43]},
      {stage1_13[42], stage1_13[43], stage1_13[44], stage1_13[45], stage1_13[46], stage1_13[47]},
      {stage2_15[7],stage2_14[14],stage2_13[15],stage2_12[15],stage2_11[20]}
   );
   gpc615_5 gpc1649 (
      {stage1_11[59], stage1_11[60], stage1_11[61], stage1_11[62], stage1_11[63]},
      {stage1_12[44]},
      {stage1_13[48], stage1_13[49], stage1_13[50], stage1_13[51], stage1_13[52], stage1_13[53]},
      {stage2_15[8],stage2_14[15],stage2_13[16],stage2_12[16],stage2_11[21]}
   );
   gpc606_5 gpc1650 (
      {stage1_14[0], stage1_14[1], stage1_14[2], stage1_14[3], stage1_14[4], stage1_14[5]},
      {stage1_16[0], stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5]},
      {stage2_18[0],stage2_17[0],stage2_16[0],stage2_15[9],stage2_14[16]}
   );
   gpc606_5 gpc1651 (
      {stage1_14[6], stage1_14[7], stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11]},
      {stage1_16[6], stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11]},
      {stage2_18[1],stage2_17[1],stage2_16[1],stage2_15[10],stage2_14[17]}
   );
   gpc606_5 gpc1652 (
      {stage1_14[12], stage1_14[13], stage1_14[14], stage1_14[15], stage1_14[16], stage1_14[17]},
      {stage1_16[12], stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17]},
      {stage2_18[2],stage2_17[2],stage2_16[2],stage2_15[11],stage2_14[18]}
   );
   gpc615_5 gpc1653 (
      {stage1_14[18], stage1_14[19], stage1_14[20], stage1_14[21], stage1_14[22]},
      {stage1_15[0]},
      {stage1_16[18], stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23]},
      {stage2_18[3],stage2_17[3],stage2_16[3],stage2_15[12],stage2_14[19]}
   );
   gpc615_5 gpc1654 (
      {stage1_14[23], stage1_14[24], stage1_14[25], stage1_14[26], stage1_14[27]},
      {stage1_15[1]},
      {stage1_16[24], stage1_16[25], stage1_16[26], stage1_16[27], stage1_16[28], stage1_16[29]},
      {stage2_18[4],stage2_17[4],stage2_16[4],stage2_15[13],stage2_14[20]}
   );
   gpc615_5 gpc1655 (
      {stage1_14[28], stage1_14[29], stage1_14[30], stage1_14[31], stage1_14[32]},
      {stage1_15[2]},
      {stage1_16[30], stage1_16[31], stage1_16[32], stage1_16[33], stage1_16[34], stage1_16[35]},
      {stage2_18[5],stage2_17[5],stage2_16[5],stage2_15[14],stage2_14[21]}
   );
   gpc615_5 gpc1656 (
      {stage1_14[33], stage1_14[34], stage1_14[35], stage1_14[36], stage1_14[37]},
      {stage1_15[3]},
      {stage1_16[36], stage1_16[37], stage1_16[38], stage1_16[39], stage1_16[40], stage1_16[41]},
      {stage2_18[6],stage2_17[6],stage2_16[6],stage2_15[15],stage2_14[22]}
   );
   gpc615_5 gpc1657 (
      {stage1_14[38], stage1_14[39], stage1_14[40], stage1_14[41], stage1_14[42]},
      {stage1_15[4]},
      {stage1_16[42], stage1_16[43], stage1_16[44], stage1_16[45], stage1_16[46], stage1_16[47]},
      {stage2_18[7],stage2_17[7],stage2_16[7],stage2_15[16],stage2_14[23]}
   );
   gpc615_5 gpc1658 (
      {stage1_14[43], stage1_14[44], stage1_14[45], stage1_14[46], stage1_14[47]},
      {stage1_15[5]},
      {stage1_16[48], stage1_16[49], stage1_16[50], stage1_16[51], stage1_16[52], stage1_16[53]},
      {stage2_18[8],stage2_17[8],stage2_16[8],stage2_15[17],stage2_14[24]}
   );
   gpc615_5 gpc1659 (
      {stage1_14[48], stage1_14[49], stage1_14[50], stage1_14[51], stage1_14[52]},
      {stage1_15[6]},
      {stage1_16[54], stage1_16[55], stage1_16[56], stage1_16[57], stage1_16[58], stage1_16[59]},
      {stage2_18[9],stage2_17[9],stage2_16[9],stage2_15[18],stage2_14[25]}
   );
   gpc1415_5 gpc1660 (
      {stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage1_16[60]},
      {stage1_17[0], stage1_17[1], stage1_17[2], stage1_17[3]},
      {stage1_18[0]},
      {stage2_19[0],stage2_18[10],stage2_17[10],stage2_16[10],stage2_15[19]}
   );
   gpc2116_5 gpc1661 (
      {stage1_15[12], stage1_15[13], stage1_15[14], stage1_15[15], stage1_15[16], stage1_15[17]},
      {stage1_16[61]},
      {stage1_17[4]},
      {stage1_18[1], stage1_18[2]},
      {stage2_19[1],stage2_18[11],stage2_17[11],stage2_16[11],stage2_15[20]}
   );
   gpc2116_5 gpc1662 (
      {stage1_15[18], stage1_15[19], stage1_15[20], stage1_15[21], stage1_15[22], stage1_15[23]},
      {stage1_16[62]},
      {stage1_17[5]},
      {stage1_18[3], stage1_18[4]},
      {stage2_19[2],stage2_18[12],stage2_17[12],stage2_16[12],stage2_15[21]}
   );
   gpc2116_5 gpc1663 (
      {stage1_15[24], stage1_15[25], stage1_15[26], stage1_15[27], stage1_15[28], stage1_15[29]},
      {stage1_16[63]},
      {stage1_17[6]},
      {stage1_18[5], stage1_18[6]},
      {stage2_19[3],stage2_18[13],stage2_17[13],stage2_16[13],stage2_15[22]}
   );
   gpc2116_5 gpc1664 (
      {stage1_15[30], stage1_15[31], stage1_15[32], stage1_15[33], stage1_15[34], stage1_15[35]},
      {stage1_16[64]},
      {stage1_17[7]},
      {stage1_18[7], stage1_18[8]},
      {stage2_19[4],stage2_18[14],stage2_17[14],stage2_16[14],stage2_15[23]}
   );
   gpc2116_5 gpc1665 (
      {stage1_15[36], stage1_15[37], stage1_15[38], stage1_15[39], stage1_15[40], stage1_15[41]},
      {stage1_16[65]},
      {stage1_17[8]},
      {stage1_18[9], stage1_18[10]},
      {stage2_19[5],stage2_18[15],stage2_17[15],stage2_16[15],stage2_15[24]}
   );
   gpc615_5 gpc1666 (
      {stage1_15[42], stage1_15[43], stage1_15[44], stage1_15[45], stage1_15[46]},
      {stage1_16[66]},
      {stage1_17[9], stage1_17[10], stage1_17[11], stage1_17[12], stage1_17[13], stage1_17[14]},
      {stage2_19[6],stage2_18[16],stage2_17[16],stage2_16[16],stage2_15[25]}
   );
   gpc615_5 gpc1667 (
      {stage1_15[47], stage1_15[48], stage1_15[49], stage1_15[50], stage1_15[51]},
      {stage1_16[67]},
      {stage1_17[15], stage1_17[16], stage1_17[17], stage1_17[18], stage1_17[19], stage1_17[20]},
      {stage2_19[7],stage2_18[17],stage2_17[17],stage2_16[17],stage2_15[26]}
   );
   gpc615_5 gpc1668 (
      {stage1_15[52], stage1_15[53], stage1_15[54], stage1_15[55], stage1_15[56]},
      {stage1_16[68]},
      {stage1_17[21], stage1_17[22], stage1_17[23], stage1_17[24], stage1_17[25], stage1_17[26]},
      {stage2_19[8],stage2_18[18],stage2_17[18],stage2_16[18],stage2_15[27]}
   );
   gpc615_5 gpc1669 (
      {stage1_15[57], stage1_15[58], stage1_15[59], stage1_15[60], stage1_15[61]},
      {stage1_16[69]},
      {stage1_17[27], stage1_17[28], stage1_17[29], stage1_17[30], stage1_17[31], stage1_17[32]},
      {stage2_19[9],stage2_18[19],stage2_17[19],stage2_16[19],stage2_15[28]}
   );
   gpc615_5 gpc1670 (
      {stage1_15[62], stage1_15[63], stage1_15[64], stage1_15[65], stage1_15[66]},
      {stage1_16[70]},
      {stage1_17[33], stage1_17[34], stage1_17[35], stage1_17[36], stage1_17[37], stage1_17[38]},
      {stage2_19[10],stage2_18[20],stage2_17[20],stage2_16[20],stage2_15[29]}
   );
   gpc606_5 gpc1671 (
      {stage1_16[71], stage1_16[72], stage1_16[73], stage1_16[74], stage1_16[75], stage1_16[76]},
      {stage1_18[11], stage1_18[12], stage1_18[13], stage1_18[14], stage1_18[15], stage1_18[16]},
      {stage2_20[0],stage2_19[11],stage2_18[21],stage2_17[21],stage2_16[21]}
   );
   gpc606_5 gpc1672 (
      {stage1_16[77], stage1_16[78], stage1_16[79], stage1_16[80], stage1_16[81], stage1_16[82]},
      {stage1_18[17], stage1_18[18], stage1_18[19], stage1_18[20], stage1_18[21], stage1_18[22]},
      {stage2_20[1],stage2_19[12],stage2_18[22],stage2_17[22],stage2_16[22]}
   );
   gpc606_5 gpc1673 (
      {stage1_16[83], stage1_16[84], stage1_16[85], stage1_16[86], stage1_16[87], stage1_16[88]},
      {stage1_18[23], stage1_18[24], stage1_18[25], stage1_18[26], stage1_18[27], stage1_18[28]},
      {stage2_20[2],stage2_19[13],stage2_18[23],stage2_17[23],stage2_16[23]}
   );
   gpc135_4 gpc1674 (
      {stage1_17[39], stage1_17[40], stage1_17[41], stage1_17[42], stage1_17[43]},
      {stage1_18[29], stage1_18[30], stage1_18[31]},
      {stage1_19[0]},
      {stage2_20[3],stage2_19[14],stage2_18[24],stage2_17[24]}
   );
   gpc1343_5 gpc1675 (
      {stage1_17[44], stage1_17[45], stage1_17[46]},
      {stage1_18[32], stage1_18[33], stage1_18[34], stage1_18[35]},
      {stage1_19[1], stage1_19[2], stage1_19[3]},
      {stage1_20[0]},
      {stage2_21[0],stage2_20[4],stage2_19[15],stage2_18[25],stage2_17[25]}
   );
   gpc1343_5 gpc1676 (
      {stage1_17[47], stage1_17[48], stage1_17[49]},
      {stage1_18[36], stage1_18[37], stage1_18[38], stage1_18[39]},
      {stage1_19[4], stage1_19[5], stage1_19[6]},
      {stage1_20[1]},
      {stage2_21[1],stage2_20[5],stage2_19[16],stage2_18[26],stage2_17[26]}
   );
   gpc606_5 gpc1677 (
      {stage1_17[50], stage1_17[51], stage1_17[52], stage1_17[53], stage1_17[54], stage1_17[55]},
      {stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11], stage1_19[12]},
      {stage2_21[2],stage2_20[6],stage2_19[17],stage2_18[27],stage2_17[27]}
   );
   gpc606_5 gpc1678 (
      {stage1_17[56], stage1_17[57], stage1_17[58], stage1_17[59], stage1_17[60], stage1_17[61]},
      {stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17], stage1_19[18]},
      {stage2_21[3],stage2_20[7],stage2_19[18],stage2_18[28],stage2_17[28]}
   );
   gpc615_5 gpc1679 (
      {stage1_19[19], stage1_19[20], stage1_19[21], stage1_19[22], stage1_19[23]},
      {stage1_20[2]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage2_23[0],stage2_22[0],stage2_21[4],stage2_20[8],stage2_19[19]}
   );
   gpc615_5 gpc1680 (
      {stage1_19[24], stage1_19[25], stage1_19[26], stage1_19[27], stage1_19[28]},
      {stage1_20[3]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage2_23[1],stage2_22[1],stage2_21[5],stage2_20[9],stage2_19[20]}
   );
   gpc615_5 gpc1681 (
      {stage1_19[29], stage1_19[30], stage1_19[31], stage1_19[32], stage1_19[33]},
      {stage1_20[4]},
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage2_23[2],stage2_22[2],stage2_21[6],stage2_20[10],stage2_19[21]}
   );
   gpc615_5 gpc1682 (
      {stage1_19[34], stage1_19[35], stage1_19[36], stage1_19[37], stage1_19[38]},
      {stage1_20[5]},
      {stage1_21[18], stage1_21[19], stage1_21[20], stage1_21[21], stage1_21[22], stage1_21[23]},
      {stage2_23[3],stage2_22[3],stage2_21[7],stage2_20[11],stage2_19[22]}
   );
   gpc615_5 gpc1683 (
      {stage1_19[39], stage1_19[40], stage1_19[41], stage1_19[42], stage1_19[43]},
      {stage1_20[6]},
      {stage1_21[24], stage1_21[25], stage1_21[26], stage1_21[27], stage1_21[28], stage1_21[29]},
      {stage2_23[4],stage2_22[4],stage2_21[8],stage2_20[12],stage2_19[23]}
   );
   gpc615_5 gpc1684 (
      {stage1_19[44], stage1_19[45], stage1_19[46], stage1_19[47], stage1_19[48]},
      {stage1_20[7]},
      {stage1_21[30], stage1_21[31], stage1_21[32], stage1_21[33], stage1_21[34], stage1_21[35]},
      {stage2_23[5],stage2_22[5],stage2_21[9],stage2_20[13],stage2_19[24]}
   );
   gpc615_5 gpc1685 (
      {stage1_19[49], stage1_19[50], stage1_19[51], stage1_19[52], stage1_19[53]},
      {stage1_20[8]},
      {stage1_21[36], stage1_21[37], stage1_21[38], stage1_21[39], stage1_21[40], stage1_21[41]},
      {stage2_23[6],stage2_22[6],stage2_21[10],stage2_20[14],stage2_19[25]}
   );
   gpc606_5 gpc1686 (
      {stage1_20[9], stage1_20[10], stage1_20[11], stage1_20[12], stage1_20[13], stage1_20[14]},
      {stage1_22[0], stage1_22[1], stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5]},
      {stage2_24[0],stage2_23[7],stage2_22[7],stage2_21[11],stage2_20[15]}
   );
   gpc606_5 gpc1687 (
      {stage1_20[15], stage1_20[16], stage1_20[17], stage1_20[18], stage1_20[19], stage1_20[20]},
      {stage1_22[6], stage1_22[7], stage1_22[8], stage1_22[9], stage1_22[10], stage1_22[11]},
      {stage2_24[1],stage2_23[8],stage2_22[8],stage2_21[12],stage2_20[16]}
   );
   gpc606_5 gpc1688 (
      {stage1_20[21], stage1_20[22], stage1_20[23], stage1_20[24], stage1_20[25], stage1_20[26]},
      {stage1_22[12], stage1_22[13], stage1_22[14], stage1_22[15], stage1_22[16], stage1_22[17]},
      {stage2_24[2],stage2_23[9],stage2_22[9],stage2_21[13],stage2_20[17]}
   );
   gpc606_5 gpc1689 (
      {stage1_20[27], stage1_20[28], stage1_20[29], stage1_20[30], stage1_20[31], stage1_20[32]},
      {stage1_22[18], stage1_22[19], stage1_22[20], stage1_22[21], stage1_22[22], stage1_22[23]},
      {stage2_24[3],stage2_23[10],stage2_22[10],stage2_21[14],stage2_20[18]}
   );
   gpc606_5 gpc1690 (
      {stage1_20[33], stage1_20[34], stage1_20[35], stage1_20[36], stage1_20[37], stage1_20[38]},
      {stage1_22[24], stage1_22[25], stage1_22[26], stage1_22[27], stage1_22[28], stage1_22[29]},
      {stage2_24[4],stage2_23[11],stage2_22[11],stage2_21[15],stage2_20[19]}
   );
   gpc606_5 gpc1691 (
      {stage1_20[39], stage1_20[40], stage1_20[41], stage1_20[42], stage1_20[43], stage1_20[44]},
      {stage1_22[30], stage1_22[31], stage1_22[32], stage1_22[33], stage1_22[34], stage1_22[35]},
      {stage2_24[5],stage2_23[12],stage2_22[12],stage2_21[16],stage2_20[20]}
   );
   gpc606_5 gpc1692 (
      {stage1_20[45], stage1_20[46], stage1_20[47], stage1_20[48], stage1_20[49], stage1_20[50]},
      {stage1_22[36], stage1_22[37], stage1_22[38], stage1_22[39], stage1_22[40], stage1_22[41]},
      {stage2_24[6],stage2_23[13],stage2_22[13],stage2_21[17],stage2_20[21]}
   );
   gpc606_5 gpc1693 (
      {stage1_20[51], stage1_20[52], stage1_20[53], stage1_20[54], stage1_20[55], stage1_20[56]},
      {stage1_22[42], stage1_22[43], stage1_22[44], stage1_22[45], stage1_22[46], stage1_22[47]},
      {stage2_24[7],stage2_23[14],stage2_22[14],stage2_21[18],stage2_20[22]}
   );
   gpc615_5 gpc1694 (
      {stage1_20[57], stage1_20[58], stage1_20[59], stage1_20[60], stage1_20[61]},
      {stage1_21[42]},
      {stage1_22[48], stage1_22[49], stage1_22[50], stage1_22[51], stage1_22[52], stage1_22[53]},
      {stage2_24[8],stage2_23[15],stage2_22[15],stage2_21[19],stage2_20[23]}
   );
   gpc606_5 gpc1695 (
      {stage1_21[43], stage1_21[44], stage1_21[45], stage1_21[46], stage1_21[47], stage1_21[48]},
      {stage1_23[0], stage1_23[1], stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5]},
      {stage2_25[0],stage2_24[9],stage2_23[16],stage2_22[16],stage2_21[20]}
   );
   gpc606_5 gpc1696 (
      {stage1_21[49], stage1_21[50], stage1_21[51], stage1_21[52], stage1_21[53], stage1_21[54]},
      {stage1_23[6], stage1_23[7], stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11]},
      {stage2_25[1],stage2_24[10],stage2_23[17],stage2_22[17],stage2_21[21]}
   );
   gpc615_5 gpc1697 (
      {stage1_23[12], stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16]},
      {stage1_24[0]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[0],stage2_25[2],stage2_24[11],stage2_23[18]}
   );
   gpc615_5 gpc1698 (
      {stage1_23[17], stage1_23[18], stage1_23[19], stage1_23[20], stage1_23[21]},
      {stage1_24[1]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[1],stage2_25[3],stage2_24[12],stage2_23[19]}
   );
   gpc615_5 gpc1699 (
      {stage1_23[22], stage1_23[23], stage1_23[24], stage1_23[25], stage1_23[26]},
      {stage1_24[2]},
      {stage1_25[12], stage1_25[13], stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17]},
      {stage2_27[2],stage2_26[2],stage2_25[4],stage2_24[13],stage2_23[20]}
   );
   gpc615_5 gpc1700 (
      {stage1_23[27], stage1_23[28], stage1_23[29], stage1_23[30], stage1_23[31]},
      {stage1_24[3]},
      {stage1_25[18], stage1_25[19], stage1_25[20], stage1_25[21], stage1_25[22], stage1_25[23]},
      {stage2_27[3],stage2_26[3],stage2_25[5],stage2_24[14],stage2_23[21]}
   );
   gpc615_5 gpc1701 (
      {stage1_23[32], stage1_23[33], stage1_23[34], stage1_23[35], stage1_23[36]},
      {stage1_24[4]},
      {stage1_25[24], stage1_25[25], stage1_25[26], stage1_25[27], stage1_25[28], stage1_25[29]},
      {stage2_27[4],stage2_26[4],stage2_25[6],stage2_24[15],stage2_23[22]}
   );
   gpc615_5 gpc1702 (
      {stage1_23[37], stage1_23[38], stage1_23[39], stage1_23[40], stage1_23[41]},
      {stage1_24[5]},
      {stage1_25[30], stage1_25[31], stage1_25[32], stage1_25[33], stage1_25[34], stage1_25[35]},
      {stage2_27[5],stage2_26[5],stage2_25[7],stage2_24[16],stage2_23[23]}
   );
   gpc615_5 gpc1703 (
      {stage1_23[42], stage1_23[43], stage1_23[44], stage1_23[45], stage1_23[46]},
      {stage1_24[6]},
      {stage1_25[36], stage1_25[37], stage1_25[38], stage1_25[39], stage1_25[40], stage1_25[41]},
      {stage2_27[6],stage2_26[6],stage2_25[8],stage2_24[17],stage2_23[24]}
   );
   gpc615_5 gpc1704 (
      {stage1_23[47], stage1_23[48], stage1_23[49], stage1_23[50], stage1_23[51]},
      {stage1_24[7]},
      {stage1_25[42], stage1_25[43], stage1_25[44], stage1_25[45], stage1_25[46], stage1_25[47]},
      {stage2_27[7],stage2_26[7],stage2_25[9],stage2_24[18],stage2_23[25]}
   );
   gpc606_5 gpc1705 (
      {stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11], stage1_24[12], stage1_24[13]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[8],stage2_26[8],stage2_25[10],stage2_24[19]}
   );
   gpc606_5 gpc1706 (
      {stage1_24[14], stage1_24[15], stage1_24[16], stage1_24[17], stage1_24[18], stage1_24[19]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[9],stage2_26[9],stage2_25[11],stage2_24[20]}
   );
   gpc606_5 gpc1707 (
      {stage1_24[20], stage1_24[21], stage1_24[22], stage1_24[23], stage1_24[24], stage1_24[25]},
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16], stage1_26[17]},
      {stage2_28[2],stage2_27[10],stage2_26[10],stage2_25[12],stage2_24[21]}
   );
   gpc606_5 gpc1708 (
      {stage1_24[26], stage1_24[27], stage1_24[28], stage1_24[29], stage1_24[30], stage1_24[31]},
      {stage1_26[18], stage1_26[19], stage1_26[20], stage1_26[21], stage1_26[22], stage1_26[23]},
      {stage2_28[3],stage2_27[11],stage2_26[11],stage2_25[13],stage2_24[22]}
   );
   gpc606_5 gpc1709 (
      {stage1_24[32], stage1_24[33], stage1_24[34], stage1_24[35], stage1_24[36], stage1_24[37]},
      {stage1_26[24], stage1_26[25], stage1_26[26], stage1_26[27], stage1_26[28], stage1_26[29]},
      {stage2_28[4],stage2_27[12],stage2_26[12],stage2_25[14],stage2_24[23]}
   );
   gpc606_5 gpc1710 (
      {stage1_24[38], stage1_24[39], stage1_24[40], stage1_24[41], stage1_24[42], stage1_24[43]},
      {stage1_26[30], stage1_26[31], stage1_26[32], stage1_26[33], stage1_26[34], stage1_26[35]},
      {stage2_28[5],stage2_27[13],stage2_26[13],stage2_25[15],stage2_24[24]}
   );
   gpc606_5 gpc1711 (
      {stage1_24[44], stage1_24[45], stage1_24[46], stage1_24[47], stage1_24[48], stage1_24[49]},
      {stage1_26[36], stage1_26[37], stage1_26[38], stage1_26[39], stage1_26[40], stage1_26[41]},
      {stage2_28[6],stage2_27[14],stage2_26[14],stage2_25[16],stage2_24[25]}
   );
   gpc606_5 gpc1712 (
      {stage1_24[50], stage1_24[51], stage1_24[52], stage1_24[53], stage1_24[54], stage1_24[55]},
      {stage1_26[42], stage1_26[43], stage1_26[44], stage1_26[45], stage1_26[46], stage1_26[47]},
      {stage2_28[7],stage2_27[15],stage2_26[15],stage2_25[17],stage2_24[26]}
   );
   gpc606_5 gpc1713 (
      {stage1_24[56], stage1_24[57], stage1_24[58], stage1_24[59], stage1_24[60], stage1_24[61]},
      {stage1_26[48], stage1_26[49], stage1_26[50], stage1_26[51], stage1_26[52], stage1_26[53]},
      {stage2_28[8],stage2_27[16],stage2_26[16],stage2_25[18],stage2_24[27]}
   );
   gpc615_5 gpc1714 (
      {stage1_26[54], stage1_26[55], stage1_26[56], stage1_26[57], stage1_26[58]},
      {stage1_27[0]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[0],stage2_28[9],stage2_27[17],stage2_26[17]}
   );
   gpc615_5 gpc1715 (
      {stage1_26[59], stage1_26[60], stage1_26[61], stage1_26[62], stage1_26[63]},
      {stage1_27[1]},
      {stage1_28[6], stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11]},
      {stage2_30[1],stage2_29[1],stage2_28[10],stage2_27[18],stage2_26[18]}
   );
   gpc615_5 gpc1716 (
      {stage1_26[64], stage1_26[65], stage1_26[66], stage1_26[67], stage1_26[68]},
      {stage1_27[2]},
      {stage1_28[12], stage1_28[13], stage1_28[14], stage1_28[15], stage1_28[16], stage1_28[17]},
      {stage2_30[2],stage2_29[2],stage2_28[11],stage2_27[19],stage2_26[19]}
   );
   gpc615_5 gpc1717 (
      {stage1_26[69], stage1_26[70], stage1_26[71], stage1_26[72], stage1_26[73]},
      {stage1_27[3]},
      {stage1_28[18], stage1_28[19], stage1_28[20], stage1_28[21], stage1_28[22], stage1_28[23]},
      {stage2_30[3],stage2_29[3],stage2_28[12],stage2_27[20],stage2_26[20]}
   );
   gpc615_5 gpc1718 (
      {stage1_26[74], stage1_26[75], stage1_26[76], stage1_26[77], stage1_26[78]},
      {stage1_27[4]},
      {stage1_28[24], stage1_28[25], stage1_28[26], stage1_28[27], stage1_28[28], stage1_28[29]},
      {stage2_30[4],stage2_29[4],stage2_28[13],stage2_27[21],stage2_26[21]}
   );
   gpc615_5 gpc1719 (
      {stage1_27[5], stage1_27[6], stage1_27[7], stage1_27[8], stage1_27[9]},
      {stage1_28[30]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[5],stage2_29[5],stage2_28[14],stage2_27[22]}
   );
   gpc615_5 gpc1720 (
      {stage1_27[10], stage1_27[11], stage1_27[12], stage1_27[13], stage1_27[14]},
      {stage1_28[31]},
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage2_31[1],stage2_30[6],stage2_29[6],stage2_28[15],stage2_27[23]}
   );
   gpc615_5 gpc1721 (
      {stage1_27[15], stage1_27[16], stage1_27[17], stage1_27[18], stage1_27[19]},
      {stage1_28[32]},
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage2_31[2],stage2_30[7],stage2_29[7],stage2_28[16],stage2_27[24]}
   );
   gpc615_5 gpc1722 (
      {stage1_27[20], stage1_27[21], stage1_27[22], stage1_27[23], stage1_27[24]},
      {stage1_28[33]},
      {stage1_29[18], stage1_29[19], stage1_29[20], stage1_29[21], stage1_29[22], stage1_29[23]},
      {stage2_31[3],stage2_30[8],stage2_29[8],stage2_28[17],stage2_27[25]}
   );
   gpc615_5 gpc1723 (
      {stage1_27[25], stage1_27[26], stage1_27[27], stage1_27[28], stage1_27[29]},
      {stage1_28[34]},
      {stage1_29[24], stage1_29[25], stage1_29[26], stage1_29[27], stage1_29[28], stage1_29[29]},
      {stage2_31[4],stage2_30[9],stage2_29[9],stage2_28[18],stage2_27[26]}
   );
   gpc615_5 gpc1724 (
      {stage1_27[30], stage1_27[31], stage1_27[32], stage1_27[33], stage1_27[34]},
      {stage1_28[35]},
      {stage1_29[30], stage1_29[31], stage1_29[32], stage1_29[33], stage1_29[34], stage1_29[35]},
      {stage2_31[5],stage2_30[10],stage2_29[10],stage2_28[19],stage2_27[27]}
   );
   gpc615_5 gpc1725 (
      {stage1_27[35], stage1_27[36], stage1_27[37], stage1_27[38], stage1_27[39]},
      {stage1_28[36]},
      {stage1_29[36], stage1_29[37], stage1_29[38], stage1_29[39], stage1_29[40], stage1_29[41]},
      {stage2_31[6],stage2_30[11],stage2_29[11],stage2_28[20],stage2_27[28]}
   );
   gpc615_5 gpc1726 (
      {stage1_27[40], stage1_27[41], stage1_27[42], stage1_27[43], stage1_27[44]},
      {stage1_28[37]},
      {stage1_29[42], stage1_29[43], stage1_29[44], stage1_29[45], stage1_29[46], stage1_29[47]},
      {stage2_31[7],stage2_30[12],stage2_29[12],stage2_28[21],stage2_27[29]}
   );
   gpc615_5 gpc1727 (
      {stage1_27[45], stage1_27[46], stage1_27[47], stage1_27[48], stage1_27[49]},
      {stage1_28[38]},
      {stage1_29[48], stage1_29[49], stage1_29[50], stage1_29[51], stage1_29[52], stage1_29[53]},
      {stage2_31[8],stage2_30[13],stage2_29[13],stage2_28[22],stage2_27[30]}
   );
   gpc615_5 gpc1728 (
      {stage1_27[50], stage1_27[51], stage1_27[52], stage1_27[53], stage1_27[54]},
      {stage1_28[39]},
      {stage1_29[54], stage1_29[55], stage1_29[56], stage1_29[57], stage1_29[58], stage1_29[59]},
      {stage2_31[9],stage2_30[14],stage2_29[14],stage2_28[23],stage2_27[31]}
   );
   gpc606_5 gpc1729 (
      {stage1_28[40], stage1_28[41], stage1_28[42], stage1_28[43], stage1_28[44], stage1_28[45]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[10],stage2_30[15],stage2_29[15],stage2_28[24]}
   );
   gpc606_5 gpc1730 (
      {stage1_29[60], stage1_29[61], stage1_29[62], stage1_29[63], stage1_29[64], stage1_29[65]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[1],stage2_31[11],stage2_30[16],stage2_29[16]}
   );
   gpc606_5 gpc1731 (
      {stage1_29[66], stage1_29[67], stage1_29[68], stage1_29[69], stage1_29[70], stage1_29[71]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[2],stage2_31[12],stage2_30[17],stage2_29[17]}
   );
   gpc606_5 gpc1732 (
      {stage1_29[72], stage1_29[73], stage1_29[74], stage1_29[75], stage1_29[76], stage1_29[77]},
      {stage1_31[12], stage1_31[13], stage1_31[14], stage1_31[15], stage1_31[16], stage1_31[17]},
      {stage2_33[2],stage2_32[3],stage2_31[13],stage2_30[18],stage2_29[18]}
   );
   gpc1406_5 gpc1733 (
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10], stage1_30[11]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3]},
      {stage1_33[0]},
      {stage2_34[0],stage2_33[3],stage2_32[4],stage2_31[14],stage2_30[19]}
   );
   gpc615_5 gpc1734 (
      {stage1_30[12], stage1_30[13], stage1_30[14], stage1_30[15], stage1_30[16]},
      {stage1_31[18]},
      {stage1_32[4], stage1_32[5], stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9]},
      {stage2_34[1],stage2_33[4],stage2_32[5],stage2_31[15],stage2_30[20]}
   );
   gpc615_5 gpc1735 (
      {stage1_30[17], stage1_30[18], stage1_30[19], stage1_30[20], stage1_30[21]},
      {stage1_31[19]},
      {stage1_32[10], stage1_32[11], stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15]},
      {stage2_34[2],stage2_33[5],stage2_32[6],stage2_31[16],stage2_30[21]}
   );
   gpc615_5 gpc1736 (
      {stage1_30[22], stage1_30[23], stage1_30[24], stage1_30[25], stage1_30[26]},
      {stage1_31[20]},
      {stage1_32[16], stage1_32[17], stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21]},
      {stage2_34[3],stage2_33[6],stage2_32[7],stage2_31[17],stage2_30[22]}
   );
   gpc615_5 gpc1737 (
      {stage1_30[27], stage1_30[28], stage1_30[29], stage1_30[30], stage1_30[31]},
      {stage1_31[21]},
      {stage1_32[22], stage1_32[23], stage1_32[24], stage1_32[25], stage1_32[26], stage1_32[27]},
      {stage2_34[4],stage2_33[7],stage2_32[8],stage2_31[18],stage2_30[23]}
   );
   gpc615_5 gpc1738 (
      {stage1_30[32], stage1_30[33], stage1_30[34], stage1_30[35], stage1_30[36]},
      {stage1_31[22]},
      {stage1_32[28], stage1_32[29], stage1_32[30], stage1_32[31], stage1_32[32], stage1_32[33]},
      {stage2_34[5],stage2_33[8],stage2_32[9],stage2_31[19],stage2_30[24]}
   );
   gpc615_5 gpc1739 (
      {stage1_30[37], stage1_30[38], stage1_30[39], stage1_30[40], stage1_30[41]},
      {stage1_31[23]},
      {stage1_32[34], stage1_32[35], stage1_32[36], stage1_32[37], stage1_32[38], stage1_32[39]},
      {stage2_34[6],stage2_33[9],stage2_32[10],stage2_31[20],stage2_30[25]}
   );
   gpc615_5 gpc1740 (
      {stage1_30[42], stage1_30[43], stage1_30[44], stage1_30[45], stage1_30[46]},
      {stage1_31[24]},
      {stage1_32[40], stage1_32[41], stage1_32[42], stage1_32[43], stage1_32[44], stage1_32[45]},
      {stage2_34[7],stage2_33[10],stage2_32[11],stage2_31[21],stage2_30[26]}
   );
   gpc606_5 gpc1741 (
      {stage1_31[25], stage1_31[26], stage1_31[27], stage1_31[28], stage1_31[29], stage1_31[30]},
      {stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4], stage1_33[5], stage1_33[6]},
      {stage2_35[0],stage2_34[8],stage2_33[11],stage2_32[12],stage2_31[22]}
   );
   gpc606_5 gpc1742 (
      {stage1_31[31], stage1_31[32], stage1_31[33], stage1_31[34], stage1_31[35], stage1_31[36]},
      {stage1_33[7], stage1_33[8], stage1_33[9], stage1_33[10], stage1_33[11], stage1_33[12]},
      {stage2_35[1],stage2_34[9],stage2_33[12],stage2_32[13],stage2_31[23]}
   );
   gpc606_5 gpc1743 (
      {stage1_31[37], stage1_31[38], stage1_31[39], stage1_31[40], stage1_31[41], stage1_31[42]},
      {stage1_33[13], stage1_33[14], stage1_33[15], stage1_33[16], stage1_33[17], stage1_33[18]},
      {stage2_35[2],stage2_34[10],stage2_33[13],stage2_32[14],stage2_31[24]}
   );
   gpc606_5 gpc1744 (
      {stage1_31[43], stage1_31[44], stage1_31[45], stage1_31[46], stage1_31[47], stage1_31[48]},
      {stage1_33[19], stage1_33[20], stage1_33[21], stage1_33[22], stage1_33[23], stage1_33[24]},
      {stage2_35[3],stage2_34[11],stage2_33[14],stage2_32[15],stage2_31[25]}
   );
   gpc606_5 gpc1745 (
      {stage1_31[49], stage1_31[50], stage1_31[51], stage1_31[52], stage1_31[53], stage1_31[54]},
      {stage1_33[25], stage1_33[26], stage1_33[27], stage1_33[28], stage1_33[29], stage1_33[30]},
      {stage2_35[4],stage2_34[12],stage2_33[15],stage2_32[16],stage2_31[26]}
   );
   gpc606_5 gpc1746 (
      {stage1_31[55], stage1_31[56], stage1_31[57], stage1_31[58], stage1_31[59], 1'b0},
      {stage1_33[31], stage1_33[32], stage1_33[33], stage1_33[34], stage1_33[35], stage1_33[36]},
      {stage2_35[5],stage2_34[13],stage2_33[16],stage2_32[17],stage2_31[27]}
   );
   gpc606_5 gpc1747 (
      {stage1_32[46], stage1_32[47], stage1_32[48], stage1_32[49], stage1_32[50], stage1_32[51]},
      {stage1_34[0], stage1_34[1], stage1_34[2], stage1_34[3], stage1_34[4], stage1_34[5]},
      {stage2_36[0],stage2_35[6],stage2_34[14],stage2_33[17],stage2_32[18]}
   );
   gpc606_5 gpc1748 (
      {stage1_32[52], stage1_32[53], stage1_32[54], stage1_32[55], stage1_32[56], stage1_32[57]},
      {stage1_34[6], stage1_34[7], stage1_34[8], stage1_34[9], stage1_34[10], stage1_34[11]},
      {stage2_36[1],stage2_35[7],stage2_34[15],stage2_33[18],stage2_32[19]}
   );
   gpc606_5 gpc1749 (
      {stage1_32[58], stage1_32[59], stage1_32[60], stage1_32[61], stage1_32[62], stage1_32[63]},
      {stage1_34[12], stage1_34[13], stage1_34[14], stage1_34[15], stage1_34[16], stage1_34[17]},
      {stage2_36[2],stage2_35[8],stage2_34[16],stage2_33[19],stage2_32[20]}
   );
   gpc606_5 gpc1750 (
      {stage1_32[64], stage1_32[65], stage1_32[66], stage1_32[67], stage1_32[68], stage1_32[69]},
      {stage1_34[18], stage1_34[19], stage1_34[20], stage1_34[21], stage1_34[22], stage1_34[23]},
      {stage2_36[3],stage2_35[9],stage2_34[17],stage2_33[20],stage2_32[21]}
   );
   gpc606_5 gpc1751 (
      {stage1_32[70], stage1_32[71], stage1_32[72], stage1_32[73], stage1_32[74], stage1_32[75]},
      {stage1_34[24], stage1_34[25], stage1_34[26], stage1_34[27], stage1_34[28], stage1_34[29]},
      {stage2_36[4],stage2_35[10],stage2_34[18],stage2_33[21],stage2_32[22]}
   );
   gpc606_5 gpc1752 (
      {stage1_32[76], stage1_32[77], stage1_32[78], stage1_32[79], stage1_32[80], stage1_32[81]},
      {stage1_34[30], stage1_34[31], stage1_34[32], stage1_34[33], stage1_34[34], stage1_34[35]},
      {stage2_36[5],stage2_35[11],stage2_34[19],stage2_33[22],stage2_32[23]}
   );
   gpc606_5 gpc1753 (
      {stage1_33[37], stage1_33[38], stage1_33[39], stage1_33[40], stage1_33[41], stage1_33[42]},
      {stage1_35[0], stage1_35[1], stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5]},
      {stage2_37[0],stage2_36[6],stage2_35[12],stage2_34[20],stage2_33[23]}
   );
   gpc606_5 gpc1754 (
      {stage1_33[43], stage1_33[44], stage1_33[45], stage1_33[46], stage1_33[47], stage1_33[48]},
      {stage1_35[6], stage1_35[7], stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11]},
      {stage2_37[1],stage2_36[7],stage2_35[13],stage2_34[21],stage2_33[24]}
   );
   gpc606_5 gpc1755 (
      {stage1_33[49], stage1_33[50], stage1_33[51], stage1_33[52], stage1_33[53], stage1_33[54]},
      {stage1_35[12], stage1_35[13], stage1_35[14], stage1_35[15], stage1_35[16], stage1_35[17]},
      {stage2_37[2],stage2_36[8],stage2_35[14],stage2_34[22],stage2_33[25]}
   );
   gpc606_5 gpc1756 (
      {stage1_33[55], stage1_33[56], stage1_33[57], stage1_33[58], stage1_33[59], stage1_33[60]},
      {stage1_35[18], stage1_35[19], stage1_35[20], stage1_35[21], stage1_35[22], stage1_35[23]},
      {stage2_37[3],stage2_36[9],stage2_35[15],stage2_34[23],stage2_33[26]}
   );
   gpc615_5 gpc1757 (
      {stage1_34[36], stage1_34[37], stage1_34[38], stage1_34[39], stage1_34[40]},
      {stage1_35[24]},
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5]},
      {stage2_38[0],stage2_37[4],stage2_36[10],stage2_35[16],stage2_34[24]}
   );
   gpc615_5 gpc1758 (
      {stage1_34[41], stage1_34[42], stage1_34[43], stage1_34[44], stage1_34[45]},
      {stage1_35[25]},
      {stage1_36[6], stage1_36[7], stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11]},
      {stage2_38[1],stage2_37[5],stage2_36[11],stage2_35[17],stage2_34[25]}
   );
   gpc615_5 gpc1759 (
      {stage1_34[46], stage1_34[47], stage1_34[48], stage1_34[49], stage1_34[50]},
      {stage1_35[26]},
      {stage1_36[12], stage1_36[13], stage1_36[14], stage1_36[15], stage1_36[16], stage1_36[17]},
      {stage2_38[2],stage2_37[6],stage2_36[12],stage2_35[18],stage2_34[26]}
   );
   gpc615_5 gpc1760 (
      {stage1_34[51], stage1_34[52], stage1_34[53], stage1_34[54], stage1_34[55]},
      {stage1_35[27]},
      {stage1_36[18], stage1_36[19], stage1_36[20], stage1_36[21], stage1_36[22], stage1_36[23]},
      {stage2_38[3],stage2_37[7],stage2_36[13],stage2_35[19],stage2_34[27]}
   );
   gpc615_5 gpc1761 (
      {stage1_34[56], stage1_34[57], stage1_34[58], stage1_34[59], stage1_34[60]},
      {stage1_35[28]},
      {stage1_36[24], stage1_36[25], stage1_36[26], stage1_36[27], stage1_36[28], stage1_36[29]},
      {stage2_38[4],stage2_37[8],stage2_36[14],stage2_35[20],stage2_34[28]}
   );
   gpc615_5 gpc1762 (
      {stage1_34[61], stage1_34[62], stage1_34[63], stage1_34[64], stage1_34[65]},
      {stage1_35[29]},
      {stage1_36[30], stage1_36[31], stage1_36[32], stage1_36[33], stage1_36[34], stage1_36[35]},
      {stage2_38[5],stage2_37[9],stage2_36[15],stage2_35[21],stage2_34[29]}
   );
   gpc606_5 gpc1763 (
      {stage1_35[30], stage1_35[31], stage1_35[32], stage1_35[33], stage1_35[34], stage1_35[35]},
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4], stage1_37[5]},
      {stage2_39[0],stage2_38[6],stage2_37[10],stage2_36[16],stage2_35[22]}
   );
   gpc606_5 gpc1764 (
      {stage1_35[36], stage1_35[37], stage1_35[38], stage1_35[39], stage1_35[40], stage1_35[41]},
      {stage1_37[6], stage1_37[7], stage1_37[8], stage1_37[9], stage1_37[10], stage1_37[11]},
      {stage2_39[1],stage2_38[7],stage2_37[11],stage2_36[17],stage2_35[23]}
   );
   gpc606_5 gpc1765 (
      {stage1_36[36], stage1_36[37], stage1_36[38], stage1_36[39], stage1_36[40], stage1_36[41]},
      {stage1_38[0], stage1_38[1], stage1_38[2], stage1_38[3], stage1_38[4], stage1_38[5]},
      {stage2_40[0],stage2_39[2],stage2_38[8],stage2_37[12],stage2_36[18]}
   );
   gpc606_5 gpc1766 (
      {stage1_36[42], stage1_36[43], stage1_36[44], stage1_36[45], stage1_36[46], stage1_36[47]},
      {stage1_38[6], stage1_38[7], stage1_38[8], stage1_38[9], stage1_38[10], stage1_38[11]},
      {stage2_40[1],stage2_39[3],stage2_38[9],stage2_37[13],stage2_36[19]}
   );
   gpc606_5 gpc1767 (
      {stage1_37[12], stage1_37[13], stage1_37[14], stage1_37[15], stage1_37[16], stage1_37[17]},
      {stage1_39[0], stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5]},
      {stage2_41[0],stage2_40[2],stage2_39[4],stage2_38[10],stage2_37[14]}
   );
   gpc606_5 gpc1768 (
      {stage1_37[18], stage1_37[19], stage1_37[20], stage1_37[21], stage1_37[22], stage1_37[23]},
      {stage1_39[6], stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11]},
      {stage2_41[1],stage2_40[3],stage2_39[5],stage2_38[11],stage2_37[15]}
   );
   gpc615_5 gpc1769 (
      {stage1_37[24], stage1_37[25], stage1_37[26], stage1_37[27], stage1_37[28]},
      {stage1_38[12]},
      {stage1_39[12], stage1_39[13], stage1_39[14], stage1_39[15], stage1_39[16], stage1_39[17]},
      {stage2_41[2],stage2_40[4],stage2_39[6],stage2_38[12],stage2_37[16]}
   );
   gpc615_5 gpc1770 (
      {stage1_37[29], stage1_37[30], stage1_37[31], stage1_37[32], stage1_37[33]},
      {stage1_38[13]},
      {stage1_39[18], stage1_39[19], stage1_39[20], stage1_39[21], stage1_39[22], stage1_39[23]},
      {stage2_41[3],stage2_40[5],stage2_39[7],stage2_38[13],stage2_37[17]}
   );
   gpc615_5 gpc1771 (
      {stage1_37[34], stage1_37[35], stage1_37[36], stage1_37[37], stage1_37[38]},
      {stage1_38[14]},
      {stage1_39[24], stage1_39[25], stage1_39[26], stage1_39[27], stage1_39[28], stage1_39[29]},
      {stage2_41[4],stage2_40[6],stage2_39[8],stage2_38[14],stage2_37[18]}
   );
   gpc615_5 gpc1772 (
      {stage1_37[39], stage1_37[40], stage1_37[41], stage1_37[42], stage1_37[43]},
      {stage1_38[15]},
      {stage1_39[30], stage1_39[31], stage1_39[32], stage1_39[33], stage1_39[34], stage1_39[35]},
      {stage2_41[5],stage2_40[7],stage2_39[9],stage2_38[15],stage2_37[19]}
   );
   gpc615_5 gpc1773 (
      {stage1_37[44], stage1_37[45], stage1_37[46], stage1_37[47], stage1_37[48]},
      {stage1_38[16]},
      {stage1_39[36], stage1_39[37], stage1_39[38], stage1_39[39], stage1_39[40], stage1_39[41]},
      {stage2_41[6],stage2_40[8],stage2_39[10],stage2_38[16],stage2_37[20]}
   );
   gpc615_5 gpc1774 (
      {stage1_37[49], stage1_37[50], stage1_37[51], stage1_37[52], stage1_37[53]},
      {stage1_38[17]},
      {stage1_39[42], stage1_39[43], stage1_39[44], stage1_39[45], stage1_39[46], stage1_39[47]},
      {stage2_41[7],stage2_40[9],stage2_39[11],stage2_38[17],stage2_37[21]}
   );
   gpc615_5 gpc1775 (
      {stage1_37[54], stage1_37[55], stage1_37[56], stage1_37[57], stage1_37[58]},
      {stage1_38[18]},
      {stage1_39[48], stage1_39[49], stage1_39[50], stage1_39[51], stage1_39[52], stage1_39[53]},
      {stage2_41[8],stage2_40[10],stage2_39[12],stage2_38[18],stage2_37[22]}
   );
   gpc615_5 gpc1776 (
      {stage1_37[59], stage1_37[60], stage1_37[61], stage1_37[62], stage1_37[63]},
      {stage1_38[19]},
      {stage1_39[54], stage1_39[55], stage1_39[56], stage1_39[57], stage1_39[58], stage1_39[59]},
      {stage2_41[9],stage2_40[11],stage2_39[13],stage2_38[19],stage2_37[23]}
   );
   gpc615_5 gpc1777 (
      {stage1_37[64], stage1_37[65], stage1_37[66], stage1_37[67], stage1_37[68]},
      {stage1_38[20]},
      {stage1_39[60], stage1_39[61], stage1_39[62], stage1_39[63], stage1_39[64], stage1_39[65]},
      {stage2_41[10],stage2_40[12],stage2_39[14],stage2_38[20],stage2_37[24]}
   );
   gpc615_5 gpc1778 (
      {stage1_37[69], stage1_37[70], stage1_37[71], stage1_37[72], stage1_37[73]},
      {stage1_38[21]},
      {stage1_39[66], stage1_39[67], stage1_39[68], stage1_39[69], stage1_39[70], stage1_39[71]},
      {stage2_41[11],stage2_40[13],stage2_39[15],stage2_38[21],stage2_37[25]}
   );
   gpc615_5 gpc1779 (
      {stage1_37[74], stage1_37[75], stage1_37[76], stage1_37[77], stage1_37[78]},
      {stage1_38[22]},
      {stage1_39[72], stage1_39[73], stage1_39[74], stage1_39[75], stage1_39[76], stage1_39[77]},
      {stage2_41[12],stage2_40[14],stage2_39[16],stage2_38[22],stage2_37[26]}
   );
   gpc615_5 gpc1780 (
      {stage1_37[79], stage1_37[80], stage1_37[81], stage1_37[82], stage1_37[83]},
      {stage1_38[23]},
      {stage1_39[78], stage1_39[79], stage1_39[80], stage1_39[81], stage1_39[82], stage1_39[83]},
      {stage2_41[13],stage2_40[15],stage2_39[17],stage2_38[23],stage2_37[27]}
   );
   gpc615_5 gpc1781 (
      {stage1_37[84], stage1_37[85], stage1_37[86], stage1_37[87], stage1_37[88]},
      {stage1_38[24]},
      {stage1_39[84], stage1_39[85], stage1_39[86], stage1_39[87], stage1_39[88], stage1_39[89]},
      {stage2_41[14],stage2_40[16],stage2_39[18],stage2_38[24],stage2_37[28]}
   );
   gpc615_5 gpc1782 (
      {stage1_38[25], stage1_38[26], stage1_38[27], stage1_38[28], stage1_38[29]},
      {stage1_39[90]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3], stage1_40[4], stage1_40[5]},
      {stage2_42[0],stage2_41[15],stage2_40[17],stage2_39[19],stage2_38[25]}
   );
   gpc615_5 gpc1783 (
      {stage1_38[30], stage1_38[31], stage1_38[32], stage1_38[33], stage1_38[34]},
      {stage1_39[91]},
      {stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10], stage1_40[11]},
      {stage2_42[1],stage2_41[16],stage2_40[18],stage2_39[20],stage2_38[26]}
   );
   gpc606_5 gpc1784 (
      {stage1_40[12], stage1_40[13], stage1_40[14], stage1_40[15], stage1_40[16], stage1_40[17]},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[0],stage2_42[2],stage2_41[17],stage2_40[19]}
   );
   gpc606_5 gpc1785 (
      {stage1_40[18], stage1_40[19], stage1_40[20], stage1_40[21], stage1_40[22], stage1_40[23]},
      {stage1_42[6], stage1_42[7], stage1_42[8], stage1_42[9], stage1_42[10], stage1_42[11]},
      {stage2_44[1],stage2_43[1],stage2_42[3],stage2_41[18],stage2_40[20]}
   );
   gpc606_5 gpc1786 (
      {stage1_40[24], stage1_40[25], stage1_40[26], stage1_40[27], stage1_40[28], stage1_40[29]},
      {stage1_42[12], stage1_42[13], stage1_42[14], stage1_42[15], stage1_42[16], stage1_42[17]},
      {stage2_44[2],stage2_43[2],stage2_42[4],stage2_41[19],stage2_40[21]}
   );
   gpc606_5 gpc1787 (
      {stage1_40[30], stage1_40[31], stage1_40[32], stage1_40[33], stage1_40[34], stage1_40[35]},
      {stage1_42[18], stage1_42[19], stage1_42[20], stage1_42[21], stage1_42[22], stage1_42[23]},
      {stage2_44[3],stage2_43[3],stage2_42[5],stage2_41[20],stage2_40[22]}
   );
   gpc606_5 gpc1788 (
      {stage1_40[36], stage1_40[37], stage1_40[38], stage1_40[39], stage1_40[40], stage1_40[41]},
      {stage1_42[24], stage1_42[25], stage1_42[26], stage1_42[27], stage1_42[28], stage1_42[29]},
      {stage2_44[4],stage2_43[4],stage2_42[6],stage2_41[21],stage2_40[23]}
   );
   gpc606_5 gpc1789 (
      {stage1_40[42], stage1_40[43], stage1_40[44], stage1_40[45], stage1_40[46], stage1_40[47]},
      {stage1_42[30], stage1_42[31], stage1_42[32], stage1_42[33], stage1_42[34], stage1_42[35]},
      {stage2_44[5],stage2_43[5],stage2_42[7],stage2_41[22],stage2_40[24]}
   );
   gpc606_5 gpc1790 (
      {stage1_40[48], stage1_40[49], stage1_40[50], stage1_40[51], stage1_40[52], stage1_40[53]},
      {stage1_42[36], stage1_42[37], stage1_42[38], stage1_42[39], stage1_42[40], stage1_42[41]},
      {stage2_44[6],stage2_43[6],stage2_42[8],stage2_41[23],stage2_40[25]}
   );
   gpc615_5 gpc1791 (
      {stage1_41[0], stage1_41[1], stage1_41[2], stage1_41[3], stage1_41[4]},
      {stage1_42[42]},
      {stage1_43[0], stage1_43[1], stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5]},
      {stage2_45[0],stage2_44[7],stage2_43[7],stage2_42[9],stage2_41[24]}
   );
   gpc615_5 gpc1792 (
      {stage1_41[5], stage1_41[6], stage1_41[7], stage1_41[8], stage1_41[9]},
      {stage1_42[43]},
      {stage1_43[6], stage1_43[7], stage1_43[8], stage1_43[9], stage1_43[10], stage1_43[11]},
      {stage2_45[1],stage2_44[8],stage2_43[8],stage2_42[10],stage2_41[25]}
   );
   gpc615_5 gpc1793 (
      {stage1_41[10], stage1_41[11], stage1_41[12], stage1_41[13], stage1_41[14]},
      {stage1_42[44]},
      {stage1_43[12], stage1_43[13], stage1_43[14], stage1_43[15], stage1_43[16], stage1_43[17]},
      {stage2_45[2],stage2_44[9],stage2_43[9],stage2_42[11],stage2_41[26]}
   );
   gpc615_5 gpc1794 (
      {stage1_41[15], stage1_41[16], stage1_41[17], stage1_41[18], stage1_41[19]},
      {stage1_42[45]},
      {stage1_43[18], stage1_43[19], stage1_43[20], stage1_43[21], stage1_43[22], stage1_43[23]},
      {stage2_45[3],stage2_44[10],stage2_43[10],stage2_42[12],stage2_41[27]}
   );
   gpc615_5 gpc1795 (
      {stage1_41[20], stage1_41[21], stage1_41[22], stage1_41[23], stage1_41[24]},
      {stage1_42[46]},
      {stage1_43[24], stage1_43[25], stage1_43[26], stage1_43[27], stage1_43[28], stage1_43[29]},
      {stage2_45[4],stage2_44[11],stage2_43[11],stage2_42[13],stage2_41[28]}
   );
   gpc615_5 gpc1796 (
      {stage1_41[25], stage1_41[26], stage1_41[27], stage1_41[28], stage1_41[29]},
      {stage1_42[47]},
      {stage1_43[30], stage1_43[31], stage1_43[32], stage1_43[33], stage1_43[34], stage1_43[35]},
      {stage2_45[5],stage2_44[12],stage2_43[12],stage2_42[14],stage2_41[29]}
   );
   gpc615_5 gpc1797 (
      {stage1_41[30], stage1_41[31], stage1_41[32], stage1_41[33], stage1_41[34]},
      {stage1_42[48]},
      {stage1_43[36], stage1_43[37], stage1_43[38], stage1_43[39], stage1_43[40], stage1_43[41]},
      {stage2_45[6],stage2_44[13],stage2_43[13],stage2_42[15],stage2_41[30]}
   );
   gpc615_5 gpc1798 (
      {stage1_41[35], stage1_41[36], stage1_41[37], stage1_41[38], stage1_41[39]},
      {stage1_42[49]},
      {stage1_43[42], stage1_43[43], stage1_43[44], stage1_43[45], stage1_43[46], stage1_43[47]},
      {stage2_45[7],stage2_44[14],stage2_43[14],stage2_42[16],stage2_41[31]}
   );
   gpc606_5 gpc1799 (
      {stage1_43[48], stage1_43[49], stage1_43[50], stage1_43[51], stage1_43[52], stage1_43[53]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5]},
      {stage2_47[0],stage2_46[0],stage2_45[8],stage2_44[15],stage2_43[15]}
   );
   gpc606_5 gpc1800 (
      {stage1_43[54], stage1_43[55], stage1_43[56], stage1_43[57], stage1_43[58], stage1_43[59]},
      {stage1_45[6], stage1_45[7], stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage2_47[1],stage2_46[1],stage2_45[9],stage2_44[16],stage2_43[16]}
   );
   gpc606_5 gpc1801 (
      {stage1_43[60], stage1_43[61], stage1_43[62], stage1_43[63], stage1_43[64], stage1_43[65]},
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15], stage1_45[16], stage1_45[17]},
      {stage2_47[2],stage2_46[2],stage2_45[10],stage2_44[17],stage2_43[17]}
   );
   gpc606_5 gpc1802 (
      {stage1_43[66], stage1_43[67], stage1_43[68], stage1_43[69], stage1_43[70], stage1_43[71]},
      {stage1_45[18], stage1_45[19], stage1_45[20], stage1_45[21], stage1_45[22], stage1_45[23]},
      {stage2_47[3],stage2_46[3],stage2_45[11],stage2_44[18],stage2_43[18]}
   );
   gpc606_5 gpc1803 (
      {stage1_43[72], stage1_43[73], stage1_43[74], stage1_43[75], stage1_43[76], stage1_43[77]},
      {stage1_45[24], stage1_45[25], stage1_45[26], stage1_45[27], stage1_45[28], stage1_45[29]},
      {stage2_47[4],stage2_46[4],stage2_45[12],stage2_44[19],stage2_43[19]}
   );
   gpc615_5 gpc1804 (
      {stage1_44[0], stage1_44[1], stage1_44[2], stage1_44[3], stage1_44[4]},
      {stage1_45[30]},
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4], stage1_46[5]},
      {stage2_48[0],stage2_47[5],stage2_46[5],stage2_45[13],stage2_44[20]}
   );
   gpc615_5 gpc1805 (
      {stage1_44[5], stage1_44[6], stage1_44[7], stage1_44[8], stage1_44[9]},
      {stage1_45[31]},
      {stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9], stage1_46[10], stage1_46[11]},
      {stage2_48[1],stage2_47[6],stage2_46[6],stage2_45[14],stage2_44[21]}
   );
   gpc615_5 gpc1806 (
      {stage1_44[10], stage1_44[11], stage1_44[12], stage1_44[13], stage1_44[14]},
      {stage1_45[32]},
      {stage1_46[12], stage1_46[13], stage1_46[14], stage1_46[15], stage1_46[16], stage1_46[17]},
      {stage2_48[2],stage2_47[7],stage2_46[7],stage2_45[15],stage2_44[22]}
   );
   gpc615_5 gpc1807 (
      {stage1_44[15], stage1_44[16], stage1_44[17], stage1_44[18], stage1_44[19]},
      {stage1_45[33]},
      {stage1_46[18], stage1_46[19], stage1_46[20], stage1_46[21], stage1_46[22], stage1_46[23]},
      {stage2_48[3],stage2_47[8],stage2_46[8],stage2_45[16],stage2_44[23]}
   );
   gpc615_5 gpc1808 (
      {stage1_44[20], stage1_44[21], stage1_44[22], stage1_44[23], stage1_44[24]},
      {stage1_45[34]},
      {stage1_46[24], stage1_46[25], stage1_46[26], stage1_46[27], stage1_46[28], stage1_46[29]},
      {stage2_48[4],stage2_47[9],stage2_46[9],stage2_45[17],stage2_44[24]}
   );
   gpc615_5 gpc1809 (
      {stage1_44[25], stage1_44[26], stage1_44[27], stage1_44[28], stage1_44[29]},
      {stage1_45[35]},
      {stage1_46[30], stage1_46[31], stage1_46[32], stage1_46[33], stage1_46[34], stage1_46[35]},
      {stage2_48[5],stage2_47[10],stage2_46[10],stage2_45[18],stage2_44[25]}
   );
   gpc615_5 gpc1810 (
      {stage1_44[30], stage1_44[31], stage1_44[32], stage1_44[33], stage1_44[34]},
      {stage1_45[36]},
      {stage1_46[36], stage1_46[37], stage1_46[38], stage1_46[39], stage1_46[40], stage1_46[41]},
      {stage2_48[6],stage2_47[11],stage2_46[11],stage2_45[19],stage2_44[26]}
   );
   gpc615_5 gpc1811 (
      {stage1_44[35], stage1_44[36], stage1_44[37], stage1_44[38], stage1_44[39]},
      {stage1_45[37]},
      {stage1_46[42], stage1_46[43], stage1_46[44], stage1_46[45], stage1_46[46], stage1_46[47]},
      {stage2_48[7],stage2_47[12],stage2_46[12],stage2_45[20],stage2_44[27]}
   );
   gpc615_5 gpc1812 (
      {stage1_44[40], stage1_44[41], stage1_44[42], stage1_44[43], stage1_44[44]},
      {stage1_45[38]},
      {stage1_46[48], stage1_46[49], stage1_46[50], stage1_46[51], stage1_46[52], stage1_46[53]},
      {stage2_48[8],stage2_47[13],stage2_46[13],stage2_45[21],stage2_44[28]}
   );
   gpc615_5 gpc1813 (
      {stage1_44[45], stage1_44[46], stage1_44[47], stage1_44[48], stage1_44[49]},
      {stage1_45[39]},
      {stage1_46[54], stage1_46[55], stage1_46[56], stage1_46[57], stage1_46[58], stage1_46[59]},
      {stage2_48[9],stage2_47[14],stage2_46[14],stage2_45[22],stage2_44[29]}
   );
   gpc117_4 gpc1814 (
      {stage1_45[40], stage1_45[41], stage1_45[42], stage1_45[43], stage1_45[44], stage1_45[45], stage1_45[46]},
      {stage1_46[60]},
      {stage1_47[0]},
      {stage2_48[10],stage2_47[15],stage2_46[15],stage2_45[23]}
   );
   gpc615_5 gpc1815 (
      {stage1_46[61], stage1_46[62], stage1_46[63], stage1_46[64], stage1_46[65]},
      {stage1_47[1]},
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5]},
      {stage2_50[0],stage2_49[0],stage2_48[11],stage2_47[16],stage2_46[16]}
   );
   gpc615_5 gpc1816 (
      {stage1_46[66], stage1_46[67], stage1_46[68], stage1_46[69], stage1_46[70]},
      {stage1_47[2]},
      {stage1_48[6], stage1_48[7], stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11]},
      {stage2_50[1],stage2_49[1],stage2_48[12],stage2_47[17],stage2_46[17]}
   );
   gpc615_5 gpc1817 (
      {stage1_46[71], stage1_46[72], stage1_46[73], stage1_46[74], stage1_46[75]},
      {stage1_47[3]},
      {stage1_48[12], stage1_48[13], stage1_48[14], stage1_48[15], stage1_48[16], stage1_48[17]},
      {stage2_50[2],stage2_49[2],stage2_48[13],stage2_47[18],stage2_46[18]}
   );
   gpc2135_5 gpc1818 (
      {stage1_47[4], stage1_47[5], stage1_47[6], stage1_47[7], stage1_47[8]},
      {stage1_48[18], stage1_48[19], stage1_48[20]},
      {stage1_49[0]},
      {stage1_50[0], stage1_50[1]},
      {stage2_51[0],stage2_50[3],stage2_49[3],stage2_48[14],stage2_47[19]}
   );
   gpc2135_5 gpc1819 (
      {stage1_47[9], stage1_47[10], stage1_47[11], stage1_47[12], stage1_47[13]},
      {stage1_48[21], stage1_48[22], stage1_48[23]},
      {stage1_49[1]},
      {stage1_50[2], stage1_50[3]},
      {stage2_51[1],stage2_50[4],stage2_49[4],stage2_48[15],stage2_47[20]}
   );
   gpc2135_5 gpc1820 (
      {stage1_47[14], stage1_47[15], stage1_47[16], stage1_47[17], stage1_47[18]},
      {stage1_48[24], stage1_48[25], stage1_48[26]},
      {stage1_49[2]},
      {stage1_50[4], stage1_50[5]},
      {stage2_51[2],stage2_50[5],stage2_49[5],stage2_48[16],stage2_47[21]}
   );
   gpc606_5 gpc1821 (
      {stage1_47[19], stage1_47[20], stage1_47[21], stage1_47[22], stage1_47[23], stage1_47[24]},
      {stage1_49[3], stage1_49[4], stage1_49[5], stage1_49[6], stage1_49[7], stage1_49[8]},
      {stage2_51[3],stage2_50[6],stage2_49[6],stage2_48[17],stage2_47[22]}
   );
   gpc606_5 gpc1822 (
      {stage1_47[25], stage1_47[26], stage1_47[27], stage1_47[28], stage1_47[29], stage1_47[30]},
      {stage1_49[9], stage1_49[10], stage1_49[11], stage1_49[12], stage1_49[13], stage1_49[14]},
      {stage2_51[4],stage2_50[7],stage2_49[7],stage2_48[18],stage2_47[23]}
   );
   gpc606_5 gpc1823 (
      {stage1_47[31], stage1_47[32], stage1_47[33], stage1_47[34], stage1_47[35], stage1_47[36]},
      {stage1_49[15], stage1_49[16], stage1_49[17], stage1_49[18], stage1_49[19], stage1_49[20]},
      {stage2_51[5],stage2_50[8],stage2_49[8],stage2_48[19],stage2_47[24]}
   );
   gpc606_5 gpc1824 (
      {stage1_47[37], stage1_47[38], stage1_47[39], stage1_47[40], stage1_47[41], stage1_47[42]},
      {stage1_49[21], stage1_49[22], stage1_49[23], stage1_49[24], stage1_49[25], stage1_49[26]},
      {stage2_51[6],stage2_50[9],stage2_49[9],stage2_48[20],stage2_47[25]}
   );
   gpc606_5 gpc1825 (
      {stage1_47[43], stage1_47[44], stage1_47[45], stage1_47[46], stage1_47[47], stage1_47[48]},
      {stage1_49[27], stage1_49[28], stage1_49[29], stage1_49[30], stage1_49[31], stage1_49[32]},
      {stage2_51[7],stage2_50[10],stage2_49[10],stage2_48[21],stage2_47[26]}
   );
   gpc615_5 gpc1826 (
      {stage1_47[49], stage1_47[50], stage1_47[51], stage1_47[52], stage1_47[53]},
      {stage1_48[27]},
      {stage1_49[33], stage1_49[34], stage1_49[35], stage1_49[36], stage1_49[37], stage1_49[38]},
      {stage2_51[8],stage2_50[11],stage2_49[11],stage2_48[22],stage2_47[27]}
   );
   gpc615_5 gpc1827 (
      {stage1_47[54], stage1_47[55], stage1_47[56], stage1_47[57], stage1_47[58]},
      {stage1_48[28]},
      {stage1_49[39], stage1_49[40], stage1_49[41], stage1_49[42], stage1_49[43], stage1_49[44]},
      {stage2_51[9],stage2_50[12],stage2_49[12],stage2_48[23],stage2_47[28]}
   );
   gpc615_5 gpc1828 (
      {stage1_47[59], stage1_47[60], stage1_47[61], stage1_47[62], stage1_47[63]},
      {stage1_48[29]},
      {stage1_49[45], stage1_49[46], stage1_49[47], stage1_49[48], stage1_49[49], stage1_49[50]},
      {stage2_51[10],stage2_50[13],stage2_49[13],stage2_48[24],stage2_47[29]}
   );
   gpc606_5 gpc1829 (
      {stage1_48[30], stage1_48[31], stage1_48[32], stage1_48[33], stage1_48[34], stage1_48[35]},
      {stage1_50[6], stage1_50[7], stage1_50[8], stage1_50[9], stage1_50[10], stage1_50[11]},
      {stage2_52[0],stage2_51[11],stage2_50[14],stage2_49[14],stage2_48[25]}
   );
   gpc606_5 gpc1830 (
      {stage1_48[36], stage1_48[37], stage1_48[38], stage1_48[39], stage1_48[40], stage1_48[41]},
      {stage1_50[12], stage1_50[13], stage1_50[14], stage1_50[15], stage1_50[16], stage1_50[17]},
      {stage2_52[1],stage2_51[12],stage2_50[15],stage2_49[15],stage2_48[26]}
   );
   gpc1163_5 gpc1831 (
      {stage1_50[18], stage1_50[19], stage1_50[20]},
      {stage1_51[0], stage1_51[1], stage1_51[2], stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage1_52[0]},
      {stage1_53[0]},
      {stage2_54[0],stage2_53[0],stage2_52[2],stage2_51[13],stage2_50[16]}
   );
   gpc1163_5 gpc1832 (
      {stage1_50[21], stage1_50[22], stage1_50[23]},
      {stage1_51[6], stage1_51[7], stage1_51[8], stage1_51[9], stage1_51[10], stage1_51[11]},
      {stage1_52[1]},
      {stage1_53[1]},
      {stage2_54[1],stage2_53[1],stage2_52[3],stage2_51[14],stage2_50[17]}
   );
   gpc1163_5 gpc1833 (
      {stage1_50[24], stage1_50[25], stage1_50[26]},
      {stage1_51[12], stage1_51[13], stage1_51[14], stage1_51[15], stage1_51[16], stage1_51[17]},
      {stage1_52[2]},
      {stage1_53[2]},
      {stage2_54[2],stage2_53[2],stage2_52[4],stage2_51[15],stage2_50[18]}
   );
   gpc1163_5 gpc1834 (
      {stage1_50[27], stage1_50[28], stage1_50[29]},
      {stage1_51[18], stage1_51[19], stage1_51[20], stage1_51[21], stage1_51[22], stage1_51[23]},
      {stage1_52[3]},
      {stage1_53[3]},
      {stage2_54[3],stage2_53[3],stage2_52[5],stage2_51[16],stage2_50[19]}
   );
   gpc1163_5 gpc1835 (
      {stage1_50[30], stage1_50[31], stage1_50[32]},
      {stage1_51[24], stage1_51[25], stage1_51[26], stage1_51[27], stage1_51[28], stage1_51[29]},
      {stage1_52[4]},
      {stage1_53[4]},
      {stage2_54[4],stage2_53[4],stage2_52[6],stage2_51[17],stage2_50[20]}
   );
   gpc1163_5 gpc1836 (
      {stage1_50[33], stage1_50[34], stage1_50[35]},
      {stage1_51[30], stage1_51[31], stage1_51[32], stage1_51[33], stage1_51[34], stage1_51[35]},
      {stage1_52[5]},
      {stage1_53[5]},
      {stage2_54[5],stage2_53[5],stage2_52[7],stage2_51[18],stage2_50[21]}
   );
   gpc615_5 gpc1837 (
      {stage1_50[36], stage1_50[37], stage1_50[38], stage1_50[39], stage1_50[40]},
      {stage1_51[36]},
      {stage1_52[6], stage1_52[7], stage1_52[8], stage1_52[9], stage1_52[10], stage1_52[11]},
      {stage2_54[6],stage2_53[6],stage2_52[8],stage2_51[19],stage2_50[22]}
   );
   gpc615_5 gpc1838 (
      {stage1_50[41], stage1_50[42], stage1_50[43], stage1_50[44], stage1_50[45]},
      {stage1_51[37]},
      {stage1_52[12], stage1_52[13], stage1_52[14], stage1_52[15], stage1_52[16], stage1_52[17]},
      {stage2_54[7],stage2_53[7],stage2_52[9],stage2_51[20],stage2_50[23]}
   );
   gpc615_5 gpc1839 (
      {stage1_50[46], stage1_50[47], stage1_50[48], stage1_50[49], stage1_50[50]},
      {stage1_51[38]},
      {stage1_52[18], stage1_52[19], stage1_52[20], stage1_52[21], stage1_52[22], stage1_52[23]},
      {stage2_54[8],stage2_53[8],stage2_52[10],stage2_51[21],stage2_50[24]}
   );
   gpc615_5 gpc1840 (
      {stage1_50[51], stage1_50[52], stage1_50[53], stage1_50[54], stage1_50[55]},
      {stage1_51[39]},
      {stage1_52[24], stage1_52[25], stage1_52[26], stage1_52[27], stage1_52[28], stage1_52[29]},
      {stage2_54[9],stage2_53[9],stage2_52[11],stage2_51[22],stage2_50[25]}
   );
   gpc615_5 gpc1841 (
      {stage1_50[56], stage1_50[57], stage1_50[58], stage1_50[59], stage1_50[60]},
      {stage1_51[40]},
      {stage1_52[30], stage1_52[31], stage1_52[32], stage1_52[33], stage1_52[34], stage1_52[35]},
      {stage2_54[10],stage2_53[10],stage2_52[12],stage2_51[23],stage2_50[26]}
   );
   gpc615_5 gpc1842 (
      {stage1_50[61], stage1_50[62], stage1_50[63], stage1_50[64], stage1_50[65]},
      {stage1_51[41]},
      {stage1_52[36], stage1_52[37], stage1_52[38], stage1_52[39], stage1_52[40], stage1_52[41]},
      {stage2_54[11],stage2_53[11],stage2_52[13],stage2_51[24],stage2_50[27]}
   );
   gpc606_5 gpc1843 (
      {stage1_52[42], stage1_52[43], stage1_52[44], stage1_52[45], stage1_52[46], stage1_52[47]},
      {stage1_54[0], stage1_54[1], stage1_54[2], stage1_54[3], stage1_54[4], stage1_54[5]},
      {stage2_56[0],stage2_55[0],stage2_54[12],stage2_53[12],stage2_52[14]}
   );
   gpc606_5 gpc1844 (
      {stage1_52[48], stage1_52[49], stage1_52[50], stage1_52[51], stage1_52[52], stage1_52[53]},
      {stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9], stage1_54[10], stage1_54[11]},
      {stage2_56[1],stage2_55[1],stage2_54[13],stage2_53[13],stage2_52[15]}
   );
   gpc606_5 gpc1845 (
      {stage1_52[54], stage1_52[55], stage1_52[56], stage1_52[57], stage1_52[58], stage1_52[59]},
      {stage1_54[12], stage1_54[13], stage1_54[14], stage1_54[15], stage1_54[16], stage1_54[17]},
      {stage2_56[2],stage2_55[2],stage2_54[14],stage2_53[14],stage2_52[16]}
   );
   gpc606_5 gpc1846 (
      {stage1_53[6], stage1_53[7], stage1_53[8], stage1_53[9], stage1_53[10], stage1_53[11]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5]},
      {stage2_57[0],stage2_56[3],stage2_55[3],stage2_54[15],stage2_53[15]}
   );
   gpc606_5 gpc1847 (
      {stage1_53[12], stage1_53[13], stage1_53[14], stage1_53[15], stage1_53[16], stage1_53[17]},
      {stage1_55[6], stage1_55[7], stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11]},
      {stage2_57[1],stage2_56[4],stage2_55[4],stage2_54[16],stage2_53[16]}
   );
   gpc606_5 gpc1848 (
      {stage1_53[18], stage1_53[19], stage1_53[20], stage1_53[21], stage1_53[22], stage1_53[23]},
      {stage1_55[12], stage1_55[13], stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17]},
      {stage2_57[2],stage2_56[5],stage2_55[5],stage2_54[17],stage2_53[17]}
   );
   gpc606_5 gpc1849 (
      {stage1_53[24], stage1_53[25], stage1_53[26], stage1_53[27], stage1_53[28], stage1_53[29]},
      {stage1_55[18], stage1_55[19], stage1_55[20], stage1_55[21], stage1_55[22], stage1_55[23]},
      {stage2_57[3],stage2_56[6],stage2_55[6],stage2_54[18],stage2_53[18]}
   );
   gpc615_5 gpc1850 (
      {stage1_53[30], stage1_53[31], stage1_53[32], stage1_53[33], stage1_53[34]},
      {stage1_54[18]},
      {stage1_55[24], stage1_55[25], stage1_55[26], stage1_55[27], stage1_55[28], stage1_55[29]},
      {stage2_57[4],stage2_56[7],stage2_55[7],stage2_54[19],stage2_53[19]}
   );
   gpc615_5 gpc1851 (
      {stage1_53[35], stage1_53[36], stage1_53[37], stage1_53[38], stage1_53[39]},
      {stage1_54[19]},
      {stage1_55[30], stage1_55[31], stage1_55[32], stage1_55[33], stage1_55[34], stage1_55[35]},
      {stage2_57[5],stage2_56[8],stage2_55[8],stage2_54[20],stage2_53[20]}
   );
   gpc615_5 gpc1852 (
      {stage1_53[40], stage1_53[41], stage1_53[42], stage1_53[43], stage1_53[44]},
      {stage1_54[20]},
      {stage1_55[36], stage1_55[37], stage1_55[38], stage1_55[39], stage1_55[40], stage1_55[41]},
      {stage2_57[6],stage2_56[9],stage2_55[9],stage2_54[21],stage2_53[21]}
   );
   gpc615_5 gpc1853 (
      {stage1_54[21], stage1_54[22], stage1_54[23], stage1_54[24], stage1_54[25]},
      {stage1_55[42]},
      {stage1_56[0], stage1_56[1], stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage2_58[0],stage2_57[7],stage2_56[10],stage2_55[10],stage2_54[22]}
   );
   gpc615_5 gpc1854 (
      {stage1_54[26], stage1_54[27], stage1_54[28], stage1_54[29], stage1_54[30]},
      {stage1_55[43]},
      {stage1_56[6], stage1_56[7], stage1_56[8], stage1_56[9], stage1_56[10], stage1_56[11]},
      {stage2_58[1],stage2_57[8],stage2_56[11],stage2_55[11],stage2_54[23]}
   );
   gpc615_5 gpc1855 (
      {stage1_54[31], stage1_54[32], stage1_54[33], stage1_54[34], stage1_54[35]},
      {stage1_55[44]},
      {stage1_56[12], stage1_56[13], stage1_56[14], stage1_56[15], stage1_56[16], stage1_56[17]},
      {stage2_58[2],stage2_57[9],stage2_56[12],stage2_55[12],stage2_54[24]}
   );
   gpc615_5 gpc1856 (
      {stage1_54[36], stage1_54[37], stage1_54[38], stage1_54[39], stage1_54[40]},
      {stage1_55[45]},
      {stage1_56[18], stage1_56[19], stage1_56[20], stage1_56[21], stage1_56[22], stage1_56[23]},
      {stage2_58[3],stage2_57[10],stage2_56[13],stage2_55[13],stage2_54[25]}
   );
   gpc615_5 gpc1857 (
      {stage1_54[41], stage1_54[42], stage1_54[43], stage1_54[44], stage1_54[45]},
      {stage1_55[46]},
      {stage1_56[24], stage1_56[25], stage1_56[26], stage1_56[27], stage1_56[28], stage1_56[29]},
      {stage2_58[4],stage2_57[11],stage2_56[14],stage2_55[14],stage2_54[26]}
   );
   gpc615_5 gpc1858 (
      {stage1_54[46], stage1_54[47], stage1_54[48], stage1_54[49], stage1_54[50]},
      {stage1_55[47]},
      {stage1_56[30], stage1_56[31], stage1_56[32], stage1_56[33], stage1_56[34], stage1_56[35]},
      {stage2_58[5],stage2_57[12],stage2_56[15],stage2_55[15],stage2_54[27]}
   );
   gpc615_5 gpc1859 (
      {stage1_55[48], stage1_55[49], stage1_55[50], stage1_55[51], stage1_55[52]},
      {stage1_56[36]},
      {stage1_57[0], stage1_57[1], stage1_57[2], stage1_57[3], stage1_57[4], stage1_57[5]},
      {stage2_59[0],stage2_58[6],stage2_57[13],stage2_56[16],stage2_55[16]}
   );
   gpc615_5 gpc1860 (
      {stage1_55[53], stage1_55[54], stage1_55[55], stage1_55[56], stage1_55[57]},
      {stage1_56[37]},
      {stage1_57[6], stage1_57[7], stage1_57[8], stage1_57[9], stage1_57[10], stage1_57[11]},
      {stage2_59[1],stage2_58[7],stage2_57[14],stage2_56[17],stage2_55[17]}
   );
   gpc615_5 gpc1861 (
      {stage1_55[58], stage1_55[59], stage1_55[60], stage1_55[61], stage1_55[62]},
      {stage1_56[38]},
      {stage1_57[12], stage1_57[13], stage1_57[14], stage1_57[15], stage1_57[16], stage1_57[17]},
      {stage2_59[2],stage2_58[8],stage2_57[15],stage2_56[18],stage2_55[18]}
   );
   gpc615_5 gpc1862 (
      {stage1_55[63], stage1_55[64], stage1_55[65], stage1_55[66], stage1_55[67]},
      {stage1_56[39]},
      {stage1_57[18], stage1_57[19], stage1_57[20], stage1_57[21], stage1_57[22], stage1_57[23]},
      {stage2_59[3],stage2_58[9],stage2_57[16],stage2_56[19],stage2_55[19]}
   );
   gpc606_5 gpc1863 (
      {stage1_56[40], stage1_56[41], stage1_56[42], stage1_56[43], stage1_56[44], stage1_56[45]},
      {stage1_58[0], stage1_58[1], stage1_58[2], stage1_58[3], stage1_58[4], stage1_58[5]},
      {stage2_60[0],stage2_59[4],stage2_58[10],stage2_57[17],stage2_56[20]}
   );
   gpc606_5 gpc1864 (
      {stage1_56[46], stage1_56[47], stage1_56[48], stage1_56[49], stage1_56[50], stage1_56[51]},
      {stage1_58[6], stage1_58[7], stage1_58[8], stage1_58[9], stage1_58[10], stage1_58[11]},
      {stage2_60[1],stage2_59[5],stage2_58[11],stage2_57[18],stage2_56[21]}
   );
   gpc606_5 gpc1865 (
      {stage1_57[24], stage1_57[25], stage1_57[26], stage1_57[27], stage1_57[28], stage1_57[29]},
      {stage1_59[0], stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5]},
      {stage2_61[0],stage2_60[2],stage2_59[6],stage2_58[12],stage2_57[19]}
   );
   gpc606_5 gpc1866 (
      {stage1_57[30], stage1_57[31], stage1_57[32], stage1_57[33], stage1_57[34], stage1_57[35]},
      {stage1_59[6], stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10], stage1_59[11]},
      {stage2_61[1],stage2_60[3],stage2_59[7],stage2_58[13],stage2_57[20]}
   );
   gpc606_5 gpc1867 (
      {stage1_57[36], stage1_57[37], stage1_57[38], stage1_57[39], stage1_57[40], stage1_57[41]},
      {stage1_59[12], stage1_59[13], stage1_59[14], stage1_59[15], stage1_59[16], stage1_59[17]},
      {stage2_61[2],stage2_60[4],stage2_59[8],stage2_58[14],stage2_57[21]}
   );
   gpc606_5 gpc1868 (
      {stage1_57[42], stage1_57[43], stage1_57[44], stage1_57[45], stage1_57[46], stage1_57[47]},
      {stage1_59[18], stage1_59[19], stage1_59[20], stage1_59[21], stage1_59[22], stage1_59[23]},
      {stage2_61[3],stage2_60[5],stage2_59[9],stage2_58[15],stage2_57[22]}
   );
   gpc606_5 gpc1869 (
      {stage1_58[12], stage1_58[13], stage1_58[14], stage1_58[15], stage1_58[16], stage1_58[17]},
      {stage1_60[0], stage1_60[1], stage1_60[2], stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage2_62[0],stage2_61[4],stage2_60[6],stage2_59[10],stage2_58[16]}
   );
   gpc606_5 gpc1870 (
      {stage1_58[18], stage1_58[19], stage1_58[20], stage1_58[21], stage1_58[22], stage1_58[23]},
      {stage1_60[6], stage1_60[7], stage1_60[8], stage1_60[9], stage1_60[10], stage1_60[11]},
      {stage2_62[1],stage2_61[5],stage2_60[7],stage2_59[11],stage2_58[17]}
   );
   gpc606_5 gpc1871 (
      {stage1_58[24], stage1_58[25], stage1_58[26], stage1_58[27], stage1_58[28], stage1_58[29]},
      {stage1_60[12], stage1_60[13], stage1_60[14], stage1_60[15], stage1_60[16], stage1_60[17]},
      {stage2_62[2],stage2_61[6],stage2_60[8],stage2_59[12],stage2_58[18]}
   );
   gpc606_5 gpc1872 (
      {stage1_58[30], stage1_58[31], stage1_58[32], stage1_58[33], stage1_58[34], stage1_58[35]},
      {stage1_60[18], stage1_60[19], stage1_60[20], stage1_60[21], stage1_60[22], stage1_60[23]},
      {stage2_62[3],stage2_61[7],stage2_60[9],stage2_59[13],stage2_58[19]}
   );
   gpc606_5 gpc1873 (
      {stage1_58[36], stage1_58[37], stage1_58[38], stage1_58[39], stage1_58[40], stage1_58[41]},
      {stage1_60[24], stage1_60[25], stage1_60[26], stage1_60[27], stage1_60[28], stage1_60[29]},
      {stage2_62[4],stage2_61[8],stage2_60[10],stage2_59[14],stage2_58[20]}
   );
   gpc606_5 gpc1874 (
      {stage1_58[42], stage1_58[43], stage1_58[44], stage1_58[45], stage1_58[46], stage1_58[47]},
      {stage1_60[30], stage1_60[31], stage1_60[32], stage1_60[33], stage1_60[34], stage1_60[35]},
      {stage2_62[5],stage2_61[9],stage2_60[11],stage2_59[15],stage2_58[21]}
   );
   gpc606_5 gpc1875 (
      {stage1_58[48], stage1_58[49], stage1_58[50], stage1_58[51], stage1_58[52], stage1_58[53]},
      {stage1_60[36], stage1_60[37], stage1_60[38], stage1_60[39], stage1_60[40], stage1_60[41]},
      {stage2_62[6],stage2_61[10],stage2_60[12],stage2_59[16],stage2_58[22]}
   );
   gpc606_5 gpc1876 (
      {stage1_58[54], stage1_58[55], stage1_58[56], stage1_58[57], stage1_58[58], stage1_58[59]},
      {stage1_60[42], stage1_60[43], stage1_60[44], stage1_60[45], stage1_60[46], stage1_60[47]},
      {stage2_62[7],stage2_61[11],stage2_60[13],stage2_59[17],stage2_58[23]}
   );
   gpc606_5 gpc1877 (
      {stage1_59[24], stage1_59[25], stage1_59[26], stage1_59[27], stage1_59[28], stage1_59[29]},
      {stage1_61[0], stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5]},
      {stage2_63[0],stage2_62[8],stage2_61[12],stage2_60[14],stage2_59[18]}
   );
   gpc606_5 gpc1878 (
      {stage1_59[30], stage1_59[31], stage1_59[32], stage1_59[33], stage1_59[34], stage1_59[35]},
      {stage1_61[6], stage1_61[7], stage1_61[8], stage1_61[9], stage1_61[10], stage1_61[11]},
      {stage2_63[1],stage2_62[9],stage2_61[13],stage2_60[15],stage2_59[19]}
   );
   gpc606_5 gpc1879 (
      {stage1_59[36], stage1_59[37], stage1_59[38], stage1_59[39], stage1_59[40], stage1_59[41]},
      {stage1_61[12], stage1_61[13], stage1_61[14], stage1_61[15], stage1_61[16], stage1_61[17]},
      {stage2_63[2],stage2_62[10],stage2_61[14],stage2_60[16],stage2_59[20]}
   );
   gpc1163_5 gpc1880 (
      {stage1_61[18], stage1_61[19], stage1_61[20]},
      {stage1_62[0], stage1_62[1], stage1_62[2], stage1_62[3], stage1_62[4], stage1_62[5]},
      {stage1_63[0]},
      {stage1_64[0]},
      {stage2_65[0],stage2_64[0],stage2_63[3],stage2_62[11],stage2_61[15]}
   );
   gpc1163_5 gpc1881 (
      {stage1_61[21], stage1_61[22], stage1_61[23]},
      {stage1_62[6], stage1_62[7], stage1_62[8], stage1_62[9], stage1_62[10], stage1_62[11]},
      {stage1_63[1]},
      {stage1_64[1]},
      {stage2_65[1],stage2_64[1],stage2_63[4],stage2_62[12],stage2_61[16]}
   );
   gpc1163_5 gpc1882 (
      {stage1_61[24], stage1_61[25], stage1_61[26]},
      {stage1_62[12], stage1_62[13], stage1_62[14], stage1_62[15], stage1_62[16], stage1_62[17]},
      {stage1_63[2]},
      {stage1_64[2]},
      {stage2_65[2],stage2_64[2],stage2_63[5],stage2_62[13],stage2_61[17]}
   );
   gpc1163_5 gpc1883 (
      {stage1_61[27], stage1_61[28], stage1_61[29]},
      {stage1_62[18], stage1_62[19], stage1_62[20], stage1_62[21], stage1_62[22], stage1_62[23]},
      {stage1_63[3]},
      {stage1_64[3]},
      {stage2_65[3],stage2_64[3],stage2_63[6],stage2_62[14],stage2_61[18]}
   );
   gpc1163_5 gpc1884 (
      {stage1_61[30], stage1_61[31], stage1_61[32]},
      {stage1_62[24], stage1_62[25], stage1_62[26], stage1_62[27], stage1_62[28], stage1_62[29]},
      {stage1_63[4]},
      {stage1_64[4]},
      {stage2_65[4],stage2_64[4],stage2_63[7],stage2_62[15],stage2_61[19]}
   );
   gpc1163_5 gpc1885 (
      {stage1_61[33], stage1_61[34], stage1_61[35]},
      {stage1_62[30], stage1_62[31], stage1_62[32], stage1_62[33], stage1_62[34], stage1_62[35]},
      {stage1_63[5]},
      {stage1_64[5]},
      {stage2_65[5],stage2_64[5],stage2_63[8],stage2_62[16],stage2_61[20]}
   );
   gpc1163_5 gpc1886 (
      {stage1_61[36], stage1_61[37], stage1_61[38]},
      {stage1_62[36], stage1_62[37], stage1_62[38], stage1_62[39], stage1_62[40], stage1_62[41]},
      {stage1_63[6]},
      {stage1_64[6]},
      {stage2_65[6],stage2_64[6],stage2_63[9],stage2_62[17],stage2_61[21]}
   );
   gpc1163_5 gpc1887 (
      {stage1_61[39], stage1_61[40], stage1_61[41]},
      {stage1_62[42], stage1_62[43], stage1_62[44], stage1_62[45], stage1_62[46], stage1_62[47]},
      {stage1_63[7]},
      {stage1_64[7]},
      {stage2_65[7],stage2_64[7],stage2_63[10],stage2_62[18],stage2_61[22]}
   );
   gpc1163_5 gpc1888 (
      {stage1_61[42], stage1_61[43], stage1_61[44]},
      {stage1_62[48], stage1_62[49], stage1_62[50], stage1_62[51], stage1_62[52], stage1_62[53]},
      {stage1_63[8]},
      {stage1_64[8]},
      {stage2_65[8],stage2_64[8],stage2_63[11],stage2_62[19],stage2_61[23]}
   );
   gpc1163_5 gpc1889 (
      {stage1_61[45], stage1_61[46], stage1_61[47]},
      {stage1_62[54], stage1_62[55], stage1_62[56], stage1_62[57], stage1_62[58], stage1_62[59]},
      {stage1_63[9]},
      {stage1_64[9]},
      {stage2_65[9],stage2_64[9],stage2_63[12],stage2_62[20],stage2_61[24]}
   );
   gpc1163_5 gpc1890 (
      {stage1_61[48], stage1_61[49], stage1_61[50]},
      {stage1_62[60], stage1_62[61], stage1_62[62], stage1_62[63], stage1_62[64], stage1_62[65]},
      {stage1_63[10]},
      {stage1_64[10]},
      {stage2_65[10],stage2_64[10],stage2_63[13],stage2_62[21],stage2_61[25]}
   );
   gpc606_5 gpc1891 (
      {stage1_61[51], stage1_61[52], stage1_61[53], stage1_61[54], stage1_61[55], stage1_61[56]},
      {stage1_63[11], stage1_63[12], stage1_63[13], stage1_63[14], stage1_63[15], stage1_63[16]},
      {stage2_65[11],stage2_64[11],stage2_63[14],stage2_62[22],stage2_61[26]}
   );
   gpc2135_5 gpc1892 (
      {stage1_62[66], stage1_62[67], stage1_62[68], stage1_62[69], stage1_62[70]},
      {stage1_63[17], stage1_63[18], stage1_63[19]},
      {stage1_64[11]},
      {stage1_65[0], stage1_65[1]},
      {stage2_66[0],stage2_65[12],stage2_64[12],stage2_63[15],stage2_62[23]}
   );
   gpc2135_5 gpc1893 (
      {stage1_62[71], stage1_62[72], stage1_62[73], stage1_62[74], stage1_62[75]},
      {stage1_63[20], stage1_63[21], stage1_63[22]},
      {stage1_64[12]},
      {stage1_65[2], stage1_65[3]},
      {stage2_66[1],stage2_65[13],stage2_64[13],stage2_63[16],stage2_62[24]}
   );
   gpc2135_5 gpc1894 (
      {stage1_62[76], stage1_62[77], stage1_62[78], stage1_62[79], stage1_62[80]},
      {stage1_63[23], stage1_63[24], stage1_63[25]},
      {stage1_64[13]},
      {stage1_65[4], stage1_65[5]},
      {stage2_66[2],stage2_65[14],stage2_64[14],stage2_63[17],stage2_62[25]}
   );
   gpc606_5 gpc1895 (
      {stage1_62[81], stage1_62[82], stage1_62[83], stage1_62[84], stage1_62[85], stage1_62[86]},
      {stage1_64[14], stage1_64[15], stage1_64[16], stage1_64[17], stage1_64[18], stage1_64[19]},
      {stage2_66[3],stage2_65[15],stage2_64[15],stage2_63[18],stage2_62[26]}
   );
   gpc615_5 gpc1896 (
      {stage1_63[26], stage1_63[27], stage1_63[28], stage1_63[29], stage1_63[30]},
      {stage1_64[20]},
      {stage1_65[6], stage1_65[7], stage1_65[8], stage1_65[9], stage1_65[10], stage1_65[11]},
      {stage2_67[0],stage2_66[4],stage2_65[16],stage2_64[16],stage2_63[19]}
   );
   gpc615_5 gpc1897 (
      {stage1_63[31], stage1_63[32], stage1_63[33], stage1_63[34], stage1_63[35]},
      {stage1_64[21]},
      {stage1_65[12], stage1_65[13], stage1_65[14], stage1_65[15], stage1_65[16], stage1_65[17]},
      {stage2_67[1],stage2_66[5],stage2_65[17],stage2_64[17],stage2_63[20]}
   );
   gpc1_1 gpc1898 (
      {stage1_0[13]},
      {stage2_0[3]}
   );
   gpc1_1 gpc1899 (
      {stage1_0[14]},
      {stage2_0[4]}
   );
   gpc1_1 gpc1900 (
      {stage1_0[15]},
      {stage2_0[5]}
   );
   gpc1_1 gpc1901 (
      {stage1_0[16]},
      {stage2_0[6]}
   );
   gpc1_1 gpc1902 (
      {stage1_0[17]},
      {stage2_0[7]}
   );
   gpc1_1 gpc1903 (
      {stage1_0[18]},
      {stage2_0[8]}
   );
   gpc1_1 gpc1904 (
      {stage1_0[19]},
      {stage2_0[9]}
   );
   gpc1_1 gpc1905 (
      {stage1_0[20]},
      {stage2_0[10]}
   );
   gpc1_1 gpc1906 (
      {stage1_0[21]},
      {stage2_0[11]}
   );
   gpc1_1 gpc1907 (
      {stage1_0[22]},
      {stage2_0[12]}
   );
   gpc1_1 gpc1908 (
      {stage1_0[23]},
      {stage2_0[13]}
   );
   gpc1_1 gpc1909 (
      {stage1_0[24]},
      {stage2_0[14]}
   );
   gpc1_1 gpc1910 (
      {stage1_0[25]},
      {stage2_0[15]}
   );
   gpc1_1 gpc1911 (
      {stage1_0[26]},
      {stage2_0[16]}
   );
   gpc1_1 gpc1912 (
      {stage1_0[27]},
      {stage2_0[17]}
   );
   gpc1_1 gpc1913 (
      {stage1_0[28]},
      {stage2_0[18]}
   );
   gpc1_1 gpc1914 (
      {stage1_0[29]},
      {stage2_0[19]}
   );
   gpc1_1 gpc1915 (
      {stage1_1[26]},
      {stage2_1[6]}
   );
   gpc1_1 gpc1916 (
      {stage1_1[27]},
      {stage2_1[7]}
   );
   gpc1_1 gpc1917 (
      {stage1_1[28]},
      {stage2_1[8]}
   );
   gpc1_1 gpc1918 (
      {stage1_1[29]},
      {stage2_1[9]}
   );
   gpc1_1 gpc1919 (
      {stage1_1[30]},
      {stage2_1[10]}
   );
   gpc1_1 gpc1920 (
      {stage1_1[31]},
      {stage2_1[11]}
   );
   gpc1_1 gpc1921 (
      {stage1_1[32]},
      {stage2_1[12]}
   );
   gpc1_1 gpc1922 (
      {stage1_2[31]},
      {stage2_2[9]}
   );
   gpc1_1 gpc1923 (
      {stage1_2[32]},
      {stage2_2[10]}
   );
   gpc1_1 gpc1924 (
      {stage1_2[33]},
      {stage2_2[11]}
   );
   gpc1_1 gpc1925 (
      {stage1_2[34]},
      {stage2_2[12]}
   );
   gpc1_1 gpc1926 (
      {stage1_2[35]},
      {stage2_2[13]}
   );
   gpc1_1 gpc1927 (
      {stage1_2[36]},
      {stage2_2[14]}
   );
   gpc1_1 gpc1928 (
      {stage1_2[37]},
      {stage2_2[15]}
   );
   gpc1_1 gpc1929 (
      {stage1_2[38]},
      {stage2_2[16]}
   );
   gpc1_1 gpc1930 (
      {stage1_2[39]},
      {stage2_2[17]}
   );
   gpc1_1 gpc1931 (
      {stage1_2[40]},
      {stage2_2[18]}
   );
   gpc1_1 gpc1932 (
      {stage1_2[41]},
      {stage2_2[19]}
   );
   gpc1_1 gpc1933 (
      {stage1_2[42]},
      {stage2_2[20]}
   );
   gpc1_1 gpc1934 (
      {stage1_2[43]},
      {stage2_2[21]}
   );
   gpc1_1 gpc1935 (
      {stage1_2[44]},
      {stage2_2[22]}
   );
   gpc1_1 gpc1936 (
      {stage1_2[45]},
      {stage2_2[23]}
   );
   gpc1_1 gpc1937 (
      {stage1_2[46]},
      {stage2_2[24]}
   );
   gpc1_1 gpc1938 (
      {stage1_3[55]},
      {stage2_3[16]}
   );
   gpc1_1 gpc1939 (
      {stage1_3[56]},
      {stage2_3[17]}
   );
   gpc1_1 gpc1940 (
      {stage1_3[57]},
      {stage2_3[18]}
   );
   gpc1_1 gpc1941 (
      {stage1_3[58]},
      {stage2_3[19]}
   );
   gpc1_1 gpc1942 (
      {stage1_3[59]},
      {stage2_3[20]}
   );
   gpc1_1 gpc1943 (
      {stage1_3[60]},
      {stage2_3[21]}
   );
   gpc1_1 gpc1944 (
      {stage1_3[61]},
      {stage2_3[22]}
   );
   gpc1_1 gpc1945 (
      {stage1_3[62]},
      {stage2_3[23]}
   );
   gpc1_1 gpc1946 (
      {stage1_3[63]},
      {stage2_3[24]}
   );
   gpc1_1 gpc1947 (
      {stage1_3[64]},
      {stage2_3[25]}
   );
   gpc1_1 gpc1948 (
      {stage1_3[65]},
      {stage2_3[26]}
   );
   gpc1_1 gpc1949 (
      {stage1_3[66]},
      {stage2_3[27]}
   );
   gpc1_1 gpc1950 (
      {stage1_4[63]},
      {stage2_4[23]}
   );
   gpc1_1 gpc1951 (
      {stage1_4[64]},
      {stage2_4[24]}
   );
   gpc1_1 gpc1952 (
      {stage1_4[65]},
      {stage2_4[25]}
   );
   gpc1_1 gpc1953 (
      {stage1_5[43]},
      {stage2_5[20]}
   );
   gpc1_1 gpc1954 (
      {stage1_5[44]},
      {stage2_5[21]}
   );
   gpc1_1 gpc1955 (
      {stage1_5[45]},
      {stage2_5[22]}
   );
   gpc1_1 gpc1956 (
      {stage1_5[46]},
      {stage2_5[23]}
   );
   gpc1_1 gpc1957 (
      {stage1_5[47]},
      {stage2_5[24]}
   );
   gpc1_1 gpc1958 (
      {stage1_5[48]},
      {stage2_5[25]}
   );
   gpc1_1 gpc1959 (
      {stage1_5[49]},
      {stage2_5[26]}
   );
   gpc1_1 gpc1960 (
      {stage1_5[50]},
      {stage2_5[27]}
   );
   gpc1_1 gpc1961 (
      {stage1_5[51]},
      {stage2_5[28]}
   );
   gpc1_1 gpc1962 (
      {stage1_7[64]},
      {stage2_7[32]}
   );
   gpc1_1 gpc1963 (
      {stage1_7[65]},
      {stage2_7[33]}
   );
   gpc1_1 gpc1964 (
      {stage1_7[66]},
      {stage2_7[34]}
   );
   gpc1_1 gpc1965 (
      {stage1_7[67]},
      {stage2_7[35]}
   );
   gpc1_1 gpc1966 (
      {stage1_7[68]},
      {stage2_7[36]}
   );
   gpc1_1 gpc1967 (
      {stage1_7[69]},
      {stage2_7[37]}
   );
   gpc1_1 gpc1968 (
      {stage1_7[70]},
      {stage2_7[38]}
   );
   gpc1_1 gpc1969 (
      {stage1_8[59]},
      {stage2_8[25]}
   );
   gpc1_1 gpc1970 (
      {stage1_8[60]},
      {stage2_8[26]}
   );
   gpc1_1 gpc1971 (
      {stage1_8[61]},
      {stage2_8[27]}
   );
   gpc1_1 gpc1972 (
      {stage1_8[62]},
      {stage2_8[28]}
   );
   gpc1_1 gpc1973 (
      {stage1_8[63]},
      {stage2_8[29]}
   );
   gpc1_1 gpc1974 (
      {stage1_8[64]},
      {stage2_8[30]}
   );
   gpc1_1 gpc1975 (
      {stage1_8[65]},
      {stage2_8[31]}
   );
   gpc1_1 gpc1976 (
      {stage1_9[38]},
      {stage2_9[19]}
   );
   gpc1_1 gpc1977 (
      {stage1_9[39]},
      {stage2_9[20]}
   );
   gpc1_1 gpc1978 (
      {stage1_9[40]},
      {stage2_9[21]}
   );
   gpc1_1 gpc1979 (
      {stage1_9[41]},
      {stage2_9[22]}
   );
   gpc1_1 gpc1980 (
      {stage1_9[42]},
      {stage2_9[23]}
   );
   gpc1_1 gpc1981 (
      {stage1_9[43]},
      {stage2_9[24]}
   );
   gpc1_1 gpc1982 (
      {stage1_9[44]},
      {stage2_9[25]}
   );
   gpc1_1 gpc1983 (
      {stage1_9[45]},
      {stage2_9[26]}
   );
   gpc1_1 gpc1984 (
      {stage1_9[46]},
      {stage2_9[27]}
   );
   gpc1_1 gpc1985 (
      {stage1_9[47]},
      {stage2_9[28]}
   );
   gpc1_1 gpc1986 (
      {stage1_9[48]},
      {stage2_9[29]}
   );
   gpc1_1 gpc1987 (
      {stage1_9[49]},
      {stage2_9[30]}
   );
   gpc1_1 gpc1988 (
      {stage1_9[50]},
      {stage2_9[31]}
   );
   gpc1_1 gpc1989 (
      {stage1_9[51]},
      {stage2_9[32]}
   );
   gpc1_1 gpc1990 (
      {stage1_9[52]},
      {stage2_9[33]}
   );
   gpc1_1 gpc1991 (
      {stage1_9[53]},
      {stage2_9[34]}
   );
   gpc1_1 gpc1992 (
      {stage1_9[54]},
      {stage2_9[35]}
   );
   gpc1_1 gpc1993 (
      {stage1_9[55]},
      {stage2_9[36]}
   );
   gpc1_1 gpc1994 (
      {stage1_9[56]},
      {stage2_9[37]}
   );
   gpc1_1 gpc1995 (
      {stage1_9[57]},
      {stage2_9[38]}
   );
   gpc1_1 gpc1996 (
      {stage1_9[58]},
      {stage2_9[39]}
   );
   gpc1_1 gpc1997 (
      {stage1_9[59]},
      {stage2_9[40]}
   );
   gpc1_1 gpc1998 (
      {stage1_9[60]},
      {stage2_9[41]}
   );
   gpc1_1 gpc1999 (
      {stage1_10[36]},
      {stage2_10[26]}
   );
   gpc1_1 gpc2000 (
      {stage1_10[37]},
      {stage2_10[27]}
   );
   gpc1_1 gpc2001 (
      {stage1_10[38]},
      {stage2_10[28]}
   );
   gpc1_1 gpc2002 (
      {stage1_10[39]},
      {stage2_10[29]}
   );
   gpc1_1 gpc2003 (
      {stage1_10[40]},
      {stage2_10[30]}
   );
   gpc1_1 gpc2004 (
      {stage1_12[45]},
      {stage2_12[17]}
   );
   gpc1_1 gpc2005 (
      {stage1_12[46]},
      {stage2_12[18]}
   );
   gpc1_1 gpc2006 (
      {stage1_12[47]},
      {stage2_12[19]}
   );
   gpc1_1 gpc2007 (
      {stage1_12[48]},
      {stage2_12[20]}
   );
   gpc1_1 gpc2008 (
      {stage1_12[49]},
      {stage2_12[21]}
   );
   gpc1_1 gpc2009 (
      {stage1_12[50]},
      {stage2_12[22]}
   );
   gpc1_1 gpc2010 (
      {stage1_12[51]},
      {stage2_12[23]}
   );
   gpc1_1 gpc2011 (
      {stage1_12[52]},
      {stage2_12[24]}
   );
   gpc1_1 gpc2012 (
      {stage1_12[53]},
      {stage2_12[25]}
   );
   gpc1_1 gpc2013 (
      {stage1_12[54]},
      {stage2_12[26]}
   );
   gpc1_1 gpc2014 (
      {stage1_12[55]},
      {stage2_12[27]}
   );
   gpc1_1 gpc2015 (
      {stage1_14[53]},
      {stage2_14[26]}
   );
   gpc1_1 gpc2016 (
      {stage1_14[54]},
      {stage2_14[27]}
   );
   gpc1_1 gpc2017 (
      {stage1_14[55]},
      {stage2_14[28]}
   );
   gpc1_1 gpc2018 (
      {stage1_14[56]},
      {stage2_14[29]}
   );
   gpc1_1 gpc2019 (
      {stage1_14[57]},
      {stage2_14[30]}
   );
   gpc1_1 gpc2020 (
      {stage1_14[58]},
      {stage2_14[31]}
   );
   gpc1_1 gpc2021 (
      {stage1_14[59]},
      {stage2_14[32]}
   );
   gpc1_1 gpc2022 (
      {stage1_14[60]},
      {stage2_14[33]}
   );
   gpc1_1 gpc2023 (
      {stage1_14[61]},
      {stage2_14[34]}
   );
   gpc1_1 gpc2024 (
      {stage1_14[62]},
      {stage2_14[35]}
   );
   gpc1_1 gpc2025 (
      {stage1_14[63]},
      {stage2_14[36]}
   );
   gpc1_1 gpc2026 (
      {stage1_14[64]},
      {stage2_14[37]}
   );
   gpc1_1 gpc2027 (
      {stage1_14[65]},
      {stage2_14[38]}
   );
   gpc1_1 gpc2028 (
      {stage1_15[67]},
      {stage2_15[30]}
   );
   gpc1_1 gpc2029 (
      {stage1_17[62]},
      {stage2_17[29]}
   );
   gpc1_1 gpc2030 (
      {stage1_17[63]},
      {stage2_17[30]}
   );
   gpc1_1 gpc2031 (
      {stage1_17[64]},
      {stage2_17[31]}
   );
   gpc1_1 gpc2032 (
      {stage1_17[65]},
      {stage2_17[32]}
   );
   gpc1_1 gpc2033 (
      {stage1_17[66]},
      {stage2_17[33]}
   );
   gpc1_1 gpc2034 (
      {stage1_18[40]},
      {stage2_18[29]}
   );
   gpc1_1 gpc2035 (
      {stage1_18[41]},
      {stage2_18[30]}
   );
   gpc1_1 gpc2036 (
      {stage1_19[54]},
      {stage2_19[26]}
   );
   gpc1_1 gpc2037 (
      {stage1_20[62]},
      {stage2_20[24]}
   );
   gpc1_1 gpc2038 (
      {stage1_20[63]},
      {stage2_20[25]}
   );
   gpc1_1 gpc2039 (
      {stage1_20[64]},
      {stage2_20[26]}
   );
   gpc1_1 gpc2040 (
      {stage1_20[65]},
      {stage2_20[27]}
   );
   gpc1_1 gpc2041 (
      {stage1_20[66]},
      {stage2_20[28]}
   );
   gpc1_1 gpc2042 (
      {stage1_20[67]},
      {stage2_20[29]}
   );
   gpc1_1 gpc2043 (
      {stage1_20[68]},
      {stage2_20[30]}
   );
   gpc1_1 gpc2044 (
      {stage1_20[69]},
      {stage2_20[31]}
   );
   gpc1_1 gpc2045 (
      {stage1_20[70]},
      {stage2_20[32]}
   );
   gpc1_1 gpc2046 (
      {stage1_20[71]},
      {stage2_20[33]}
   );
   gpc1_1 gpc2047 (
      {stage1_22[54]},
      {stage2_22[18]}
   );
   gpc1_1 gpc2048 (
      {stage1_22[55]},
      {stage2_22[19]}
   );
   gpc1_1 gpc2049 (
      {stage1_22[56]},
      {stage2_22[20]}
   );
   gpc1_1 gpc2050 (
      {stage1_22[57]},
      {stage2_22[21]}
   );
   gpc1_1 gpc2051 (
      {stage1_22[58]},
      {stage2_22[22]}
   );
   gpc1_1 gpc2052 (
      {stage1_22[59]},
      {stage2_22[23]}
   );
   gpc1_1 gpc2053 (
      {stage1_22[60]},
      {stage2_22[24]}
   );
   gpc1_1 gpc2054 (
      {stage1_22[61]},
      {stage2_22[25]}
   );
   gpc1_1 gpc2055 (
      {stage1_22[62]},
      {stage2_22[26]}
   );
   gpc1_1 gpc2056 (
      {stage1_22[63]},
      {stage2_22[27]}
   );
   gpc1_1 gpc2057 (
      {stage1_22[64]},
      {stage2_22[28]}
   );
   gpc1_1 gpc2058 (
      {stage1_22[65]},
      {stage2_22[29]}
   );
   gpc1_1 gpc2059 (
      {stage1_22[66]},
      {stage2_22[30]}
   );
   gpc1_1 gpc2060 (
      {stage1_22[67]},
      {stage2_22[31]}
   );
   gpc1_1 gpc2061 (
      {stage1_22[68]},
      {stage2_22[32]}
   );
   gpc1_1 gpc2062 (
      {stage1_22[69]},
      {stage2_22[33]}
   );
   gpc1_1 gpc2063 (
      {stage1_22[70]},
      {stage2_22[34]}
   );
   gpc1_1 gpc2064 (
      {stage1_23[52]},
      {stage2_23[26]}
   );
   gpc1_1 gpc2065 (
      {stage1_23[53]},
      {stage2_23[27]}
   );
   gpc1_1 gpc2066 (
      {stage1_25[48]},
      {stage2_25[19]}
   );
   gpc1_1 gpc2067 (
      {stage1_25[49]},
      {stage2_25[20]}
   );
   gpc1_1 gpc2068 (
      {stage1_25[50]},
      {stage2_25[21]}
   );
   gpc1_1 gpc2069 (
      {stage1_25[51]},
      {stage2_25[22]}
   );
   gpc1_1 gpc2070 (
      {stage1_25[52]},
      {stage2_25[23]}
   );
   gpc1_1 gpc2071 (
      {stage1_25[53]},
      {stage2_25[24]}
   );
   gpc1_1 gpc2072 (
      {stage1_25[54]},
      {stage2_25[25]}
   );
   gpc1_1 gpc2073 (
      {stage1_25[55]},
      {stage2_25[26]}
   );
   gpc1_1 gpc2074 (
      {stage1_25[56]},
      {stage2_25[27]}
   );
   gpc1_1 gpc2075 (
      {stage1_25[57]},
      {stage2_25[28]}
   );
   gpc1_1 gpc2076 (
      {stage1_25[58]},
      {stage2_25[29]}
   );
   gpc1_1 gpc2077 (
      {stage1_25[59]},
      {stage2_25[30]}
   );
   gpc1_1 gpc2078 (
      {stage1_25[60]},
      {stage2_25[31]}
   );
   gpc1_1 gpc2079 (
      {stage1_26[79]},
      {stage2_26[22]}
   );
   gpc1_1 gpc2080 (
      {stage1_26[80]},
      {stage2_26[23]}
   );
   gpc1_1 gpc2081 (
      {stage1_26[81]},
      {stage2_26[24]}
   );
   gpc1_1 gpc2082 (
      {stage1_26[82]},
      {stage2_26[25]}
   );
   gpc1_1 gpc2083 (
      {stage1_26[83]},
      {stage2_26[26]}
   );
   gpc1_1 gpc2084 (
      {stage1_27[55]},
      {stage2_27[32]}
   );
   gpc1_1 gpc2085 (
      {stage1_28[46]},
      {stage2_28[25]}
   );
   gpc1_1 gpc2086 (
      {stage1_28[47]},
      {stage2_28[26]}
   );
   gpc1_1 gpc2087 (
      {stage1_29[78]},
      {stage2_29[19]}
   );
   gpc1_1 gpc2088 (
      {stage1_29[79]},
      {stage2_29[20]}
   );
   gpc1_1 gpc2089 (
      {stage1_30[47]},
      {stage2_30[27]}
   );
   gpc1_1 gpc2090 (
      {stage1_30[48]},
      {stage2_30[28]}
   );
   gpc1_1 gpc2091 (
      {stage1_30[49]},
      {stage2_30[29]}
   );
   gpc1_1 gpc2092 (
      {stage1_30[50]},
      {stage2_30[30]}
   );
   gpc1_1 gpc2093 (
      {stage1_30[51]},
      {stage2_30[31]}
   );
   gpc1_1 gpc2094 (
      {stage1_30[52]},
      {stage2_30[32]}
   );
   gpc1_1 gpc2095 (
      {stage1_30[53]},
      {stage2_30[33]}
   );
   gpc1_1 gpc2096 (
      {stage1_30[54]},
      {stage2_30[34]}
   );
   gpc1_1 gpc2097 (
      {stage1_30[55]},
      {stage2_30[35]}
   );
   gpc1_1 gpc2098 (
      {stage1_30[56]},
      {stage2_30[36]}
   );
   gpc1_1 gpc2099 (
      {stage1_30[57]},
      {stage2_30[37]}
   );
   gpc1_1 gpc2100 (
      {stage1_30[58]},
      {stage2_30[38]}
   );
   gpc1_1 gpc2101 (
      {stage1_30[59]},
      {stage2_30[39]}
   );
   gpc1_1 gpc2102 (
      {stage1_30[60]},
      {stage2_30[40]}
   );
   gpc1_1 gpc2103 (
      {stage1_30[61]},
      {stage2_30[41]}
   );
   gpc1_1 gpc2104 (
      {stage1_30[62]},
      {stage2_30[42]}
   );
   gpc1_1 gpc2105 (
      {stage1_30[63]},
      {stage2_30[43]}
   );
   gpc1_1 gpc2106 (
      {stage1_30[64]},
      {stage2_30[44]}
   );
   gpc1_1 gpc2107 (
      {stage1_30[65]},
      {stage2_30[45]}
   );
   gpc1_1 gpc2108 (
      {stage1_30[66]},
      {stage2_30[46]}
   );
   gpc1_1 gpc2109 (
      {stage1_30[67]},
      {stage2_30[47]}
   );
   gpc1_1 gpc2110 (
      {stage1_30[68]},
      {stage2_30[48]}
   );
   gpc1_1 gpc2111 (
      {stage1_30[69]},
      {stage2_30[49]}
   );
   gpc1_1 gpc2112 (
      {stage1_30[70]},
      {stage2_30[50]}
   );
   gpc1_1 gpc2113 (
      {stage1_30[71]},
      {stage2_30[51]}
   );
   gpc1_1 gpc2114 (
      {stage1_32[82]},
      {stage2_32[24]}
   );
   gpc1_1 gpc2115 (
      {stage1_33[61]},
      {stage2_33[27]}
   );
   gpc1_1 gpc2116 (
      {stage1_33[62]},
      {stage2_33[28]}
   );
   gpc1_1 gpc2117 (
      {stage1_34[66]},
      {stage2_34[30]}
   );
   gpc1_1 gpc2118 (
      {stage1_34[67]},
      {stage2_34[31]}
   );
   gpc1_1 gpc2119 (
      {stage1_35[42]},
      {stage2_35[24]}
   );
   gpc1_1 gpc2120 (
      {stage1_35[43]},
      {stage2_35[25]}
   );
   gpc1_1 gpc2121 (
      {stage1_35[44]},
      {stage2_35[26]}
   );
   gpc1_1 gpc2122 (
      {stage1_35[45]},
      {stage2_35[27]}
   );
   gpc1_1 gpc2123 (
      {stage1_35[46]},
      {stage2_35[28]}
   );
   gpc1_1 gpc2124 (
      {stage1_35[47]},
      {stage2_35[29]}
   );
   gpc1_1 gpc2125 (
      {stage1_36[48]},
      {stage2_36[20]}
   );
   gpc1_1 gpc2126 (
      {stage1_36[49]},
      {stage2_36[21]}
   );
   gpc1_1 gpc2127 (
      {stage1_36[50]},
      {stage2_36[22]}
   );
   gpc1_1 gpc2128 (
      {stage1_36[51]},
      {stage2_36[23]}
   );
   gpc1_1 gpc2129 (
      {stage1_36[52]},
      {stage2_36[24]}
   );
   gpc1_1 gpc2130 (
      {stage1_36[53]},
      {stage2_36[25]}
   );
   gpc1_1 gpc2131 (
      {stage1_36[54]},
      {stage2_36[26]}
   );
   gpc1_1 gpc2132 (
      {stage1_36[55]},
      {stage2_36[27]}
   );
   gpc1_1 gpc2133 (
      {stage1_36[56]},
      {stage2_36[28]}
   );
   gpc1_1 gpc2134 (
      {stage1_36[57]},
      {stage2_36[29]}
   );
   gpc1_1 gpc2135 (
      {stage1_36[58]},
      {stage2_36[30]}
   );
   gpc1_1 gpc2136 (
      {stage1_36[59]},
      {stage2_36[31]}
   );
   gpc1_1 gpc2137 (
      {stage1_36[60]},
      {stage2_36[32]}
   );
   gpc1_1 gpc2138 (
      {stage1_37[89]},
      {stage2_37[29]}
   );
   gpc1_1 gpc2139 (
      {stage1_37[90]},
      {stage2_37[30]}
   );
   gpc1_1 gpc2140 (
      {stage1_37[91]},
      {stage2_37[31]}
   );
   gpc1_1 gpc2141 (
      {stage1_37[92]},
      {stage2_37[32]}
   );
   gpc1_1 gpc2142 (
      {stage1_37[93]},
      {stage2_37[33]}
   );
   gpc1_1 gpc2143 (
      {stage1_37[94]},
      {stage2_37[34]}
   );
   gpc1_1 gpc2144 (
      {stage1_37[95]},
      {stage2_37[35]}
   );
   gpc1_1 gpc2145 (
      {stage1_37[96]},
      {stage2_37[36]}
   );
   gpc1_1 gpc2146 (
      {stage1_38[35]},
      {stage2_38[27]}
   );
   gpc1_1 gpc2147 (
      {stage1_38[36]},
      {stage2_38[28]}
   );
   gpc1_1 gpc2148 (
      {stage1_38[37]},
      {stage2_38[29]}
   );
   gpc1_1 gpc2149 (
      {stage1_38[38]},
      {stage2_38[30]}
   );
   gpc1_1 gpc2150 (
      {stage1_38[39]},
      {stage2_38[31]}
   );
   gpc1_1 gpc2151 (
      {stage1_38[40]},
      {stage2_38[32]}
   );
   gpc1_1 gpc2152 (
      {stage1_38[41]},
      {stage2_38[33]}
   );
   gpc1_1 gpc2153 (
      {stage1_38[42]},
      {stage2_38[34]}
   );
   gpc1_1 gpc2154 (
      {stage1_38[43]},
      {stage2_38[35]}
   );
   gpc1_1 gpc2155 (
      {stage1_39[92]},
      {stage2_39[21]}
   );
   gpc1_1 gpc2156 (
      {stage1_40[54]},
      {stage2_40[26]}
   );
   gpc1_1 gpc2157 (
      {stage1_40[55]},
      {stage2_40[27]}
   );
   gpc1_1 gpc2158 (
      {stage1_40[56]},
      {stage2_40[28]}
   );
   gpc1_1 gpc2159 (
      {stage1_40[57]},
      {stage2_40[29]}
   );
   gpc1_1 gpc2160 (
      {stage1_40[58]},
      {stage2_40[30]}
   );
   gpc1_1 gpc2161 (
      {stage1_40[59]},
      {stage2_40[31]}
   );
   gpc1_1 gpc2162 (
      {stage1_40[60]},
      {stage2_40[32]}
   );
   gpc1_1 gpc2163 (
      {stage1_40[61]},
      {stage2_40[33]}
   );
   gpc1_1 gpc2164 (
      {stage1_40[62]},
      {stage2_40[34]}
   );
   gpc1_1 gpc2165 (
      {stage1_42[50]},
      {stage2_42[17]}
   );
   gpc1_1 gpc2166 (
      {stage1_43[78]},
      {stage2_43[20]}
   );
   gpc1_1 gpc2167 (
      {stage1_45[47]},
      {stage2_45[24]}
   );
   gpc1_1 gpc2168 (
      {stage1_45[48]},
      {stage2_45[25]}
   );
   gpc1_1 gpc2169 (
      {stage1_45[49]},
      {stage2_45[26]}
   );
   gpc1_1 gpc2170 (
      {stage1_45[50]},
      {stage2_45[27]}
   );
   gpc1_1 gpc2171 (
      {stage1_45[51]},
      {stage2_45[28]}
   );
   gpc1_1 gpc2172 (
      {stage1_45[52]},
      {stage2_45[29]}
   );
   gpc1_1 gpc2173 (
      {stage1_45[53]},
      {stage2_45[30]}
   );
   gpc1_1 gpc2174 (
      {stage1_45[54]},
      {stage2_45[31]}
   );
   gpc1_1 gpc2175 (
      {stage1_45[55]},
      {stage2_45[32]}
   );
   gpc1_1 gpc2176 (
      {stage1_45[56]},
      {stage2_45[33]}
   );
   gpc1_1 gpc2177 (
      {stage1_45[57]},
      {stage2_45[34]}
   );
   gpc1_1 gpc2178 (
      {stage1_46[76]},
      {stage2_46[19]}
   );
   gpc1_1 gpc2179 (
      {stage1_46[77]},
      {stage2_46[20]}
   );
   gpc1_1 gpc2180 (
      {stage1_46[78]},
      {stage2_46[21]}
   );
   gpc1_1 gpc2181 (
      {stage1_46[79]},
      {stage2_46[22]}
   );
   gpc1_1 gpc2182 (
      {stage1_47[64]},
      {stage2_47[30]}
   );
   gpc1_1 gpc2183 (
      {stage1_47[65]},
      {stage2_47[31]}
   );
   gpc1_1 gpc2184 (
      {stage1_47[66]},
      {stage2_47[32]}
   );
   gpc1_1 gpc2185 (
      {stage1_47[67]},
      {stage2_47[33]}
   );
   gpc1_1 gpc2186 (
      {stage1_47[68]},
      {stage2_47[34]}
   );
   gpc1_1 gpc2187 (
      {stage1_47[69]},
      {stage2_47[35]}
   );
   gpc1_1 gpc2188 (
      {stage1_48[42]},
      {stage2_48[27]}
   );
   gpc1_1 gpc2189 (
      {stage1_48[43]},
      {stage2_48[28]}
   );
   gpc1_1 gpc2190 (
      {stage1_48[44]},
      {stage2_48[29]}
   );
   gpc1_1 gpc2191 (
      {stage1_48[45]},
      {stage2_48[30]}
   );
   gpc1_1 gpc2192 (
      {stage1_50[66]},
      {stage2_50[28]}
   );
   gpc1_1 gpc2193 (
      {stage1_50[67]},
      {stage2_50[29]}
   );
   gpc1_1 gpc2194 (
      {stage1_50[68]},
      {stage2_50[30]}
   );
   gpc1_1 gpc2195 (
      {stage1_50[69]},
      {stage2_50[31]}
   );
   gpc1_1 gpc2196 (
      {stage1_50[70]},
      {stage2_50[32]}
   );
   gpc1_1 gpc2197 (
      {stage1_51[42]},
      {stage2_51[25]}
   );
   gpc1_1 gpc2198 (
      {stage1_51[43]},
      {stage2_51[26]}
   );
   gpc1_1 gpc2199 (
      {stage1_51[44]},
      {stage2_51[27]}
   );
   gpc1_1 gpc2200 (
      {stage1_51[45]},
      {stage2_51[28]}
   );
   gpc1_1 gpc2201 (
      {stage1_51[46]},
      {stage2_51[29]}
   );
   gpc1_1 gpc2202 (
      {stage1_51[47]},
      {stage2_51[30]}
   );
   gpc1_1 gpc2203 (
      {stage1_52[60]},
      {stage2_52[17]}
   );
   gpc1_1 gpc2204 (
      {stage1_53[45]},
      {stage2_53[22]}
   );
   gpc1_1 gpc2205 (
      {stage1_53[46]},
      {stage2_53[23]}
   );
   gpc1_1 gpc2206 (
      {stage1_53[47]},
      {stage2_53[24]}
   );
   gpc1_1 gpc2207 (
      {stage1_53[48]},
      {stage2_53[25]}
   );
   gpc1_1 gpc2208 (
      {stage1_53[49]},
      {stage2_53[26]}
   );
   gpc1_1 gpc2209 (
      {stage1_53[50]},
      {stage2_53[27]}
   );
   gpc1_1 gpc2210 (
      {stage1_53[51]},
      {stage2_53[28]}
   );
   gpc1_1 gpc2211 (
      {stage1_53[52]},
      {stage2_53[29]}
   );
   gpc1_1 gpc2212 (
      {stage1_53[53]},
      {stage2_53[30]}
   );
   gpc1_1 gpc2213 (
      {stage1_53[54]},
      {stage2_53[31]}
   );
   gpc1_1 gpc2214 (
      {stage1_53[55]},
      {stage2_53[32]}
   );
   gpc1_1 gpc2215 (
      {stage1_53[56]},
      {stage2_53[33]}
   );
   gpc1_1 gpc2216 (
      {stage1_53[57]},
      {stage2_53[34]}
   );
   gpc1_1 gpc2217 (
      {stage1_53[58]},
      {stage2_53[35]}
   );
   gpc1_1 gpc2218 (
      {stage1_53[59]},
      {stage2_53[36]}
   );
   gpc1_1 gpc2219 (
      {stage1_53[60]},
      {stage2_53[37]}
   );
   gpc1_1 gpc2220 (
      {stage1_53[61]},
      {stage2_53[38]}
   );
   gpc1_1 gpc2221 (
      {stage1_54[51]},
      {stage2_54[28]}
   );
   gpc1_1 gpc2222 (
      {stage1_56[52]},
      {stage2_56[22]}
   );
   gpc1_1 gpc2223 (
      {stage1_56[53]},
      {stage2_56[23]}
   );
   gpc1_1 gpc2224 (
      {stage1_56[54]},
      {stage2_56[24]}
   );
   gpc1_1 gpc2225 (
      {stage1_56[55]},
      {stage2_56[25]}
   );
   gpc1_1 gpc2226 (
      {stage1_56[56]},
      {stage2_56[26]}
   );
   gpc1_1 gpc2227 (
      {stage1_57[48]},
      {stage2_57[23]}
   );
   gpc1_1 gpc2228 (
      {stage1_57[49]},
      {stage2_57[24]}
   );
   gpc1_1 gpc2229 (
      {stage1_57[50]},
      {stage2_57[25]}
   );
   gpc1_1 gpc2230 (
      {stage1_57[51]},
      {stage2_57[26]}
   );
   gpc1_1 gpc2231 (
      {stage1_57[52]},
      {stage2_57[27]}
   );
   gpc1_1 gpc2232 (
      {stage1_57[53]},
      {stage2_57[28]}
   );
   gpc1_1 gpc2233 (
      {stage1_57[54]},
      {stage2_57[29]}
   );
   gpc1_1 gpc2234 (
      {stage1_57[55]},
      {stage2_57[30]}
   );
   gpc1_1 gpc2235 (
      {stage1_57[56]},
      {stage2_57[31]}
   );
   gpc1_1 gpc2236 (
      {stage1_57[57]},
      {stage2_57[32]}
   );
   gpc1_1 gpc2237 (
      {stage1_59[42]},
      {stage2_59[21]}
   );
   gpc1_1 gpc2238 (
      {stage1_59[43]},
      {stage2_59[22]}
   );
   gpc1_1 gpc2239 (
      {stage1_59[44]},
      {stage2_59[23]}
   );
   gpc1_1 gpc2240 (
      {stage1_59[45]},
      {stage2_59[24]}
   );
   gpc1_1 gpc2241 (
      {stage1_59[46]},
      {stage2_59[25]}
   );
   gpc1_1 gpc2242 (
      {stage1_59[47]},
      {stage2_59[26]}
   );
   gpc1_1 gpc2243 (
      {stage1_59[48]},
      {stage2_59[27]}
   );
   gpc1_1 gpc2244 (
      {stage1_59[49]},
      {stage2_59[28]}
   );
   gpc1_1 gpc2245 (
      {stage1_59[50]},
      {stage2_59[29]}
   );
   gpc1_1 gpc2246 (
      {stage1_59[51]},
      {stage2_59[30]}
   );
   gpc1_1 gpc2247 (
      {stage1_59[52]},
      {stage2_59[31]}
   );
   gpc1_1 gpc2248 (
      {stage1_59[53]},
      {stage2_59[32]}
   );
   gpc1_1 gpc2249 (
      {stage1_59[54]},
      {stage2_59[33]}
   );
   gpc1_1 gpc2250 (
      {stage1_59[55]},
      {stage2_59[34]}
   );
   gpc1_1 gpc2251 (
      {stage1_60[48]},
      {stage2_60[17]}
   );
   gpc1_1 gpc2252 (
      {stage1_60[49]},
      {stage2_60[18]}
   );
   gpc1_1 gpc2253 (
      {stage1_60[50]},
      {stage2_60[19]}
   );
   gpc1_1 gpc2254 (
      {stage1_60[51]},
      {stage2_60[20]}
   );
   gpc1_1 gpc2255 (
      {stage1_60[52]},
      {stage2_60[21]}
   );
   gpc1_1 gpc2256 (
      {stage1_61[57]},
      {stage2_61[27]}
   );
   gpc1_1 gpc2257 (
      {stage1_61[58]},
      {stage2_61[28]}
   );
   gpc1_1 gpc2258 (
      {stage1_62[87]},
      {stage2_62[27]}
   );
   gpc1_1 gpc2259 (
      {stage1_62[88]},
      {stage2_62[28]}
   );
   gpc1_1 gpc2260 (
      {stage1_62[89]},
      {stage2_62[29]}
   );
   gpc1_1 gpc2261 (
      {stage1_62[90]},
      {stage2_62[30]}
   );
   gpc1_1 gpc2262 (
      {stage1_62[91]},
      {stage2_62[31]}
   );
   gpc1_1 gpc2263 (
      {stage1_62[92]},
      {stage2_62[32]}
   );
   gpc1_1 gpc2264 (
      {stage1_62[93]},
      {stage2_62[33]}
   );
   gpc1_1 gpc2265 (
      {stage1_62[94]},
      {stage2_62[34]}
   );
   gpc1_1 gpc2266 (
      {stage1_62[95]},
      {stage2_62[35]}
   );
   gpc1_1 gpc2267 (
      {stage1_62[96]},
      {stage2_62[36]}
   );
   gpc1_1 gpc2268 (
      {stage1_62[97]},
      {stage2_62[37]}
   );
   gpc1_1 gpc2269 (
      {stage1_63[36]},
      {stage2_63[21]}
   );
   gpc1_1 gpc2270 (
      {stage1_63[37]},
      {stage2_63[22]}
   );
   gpc1_1 gpc2271 (
      {stage1_63[38]},
      {stage2_63[23]}
   );
   gpc1_1 gpc2272 (
      {stage1_63[39]},
      {stage2_63[24]}
   );
   gpc1_1 gpc2273 (
      {stage1_63[40]},
      {stage2_63[25]}
   );
   gpc1_1 gpc2274 (
      {stage1_63[41]},
      {stage2_63[26]}
   );
   gpc1_1 gpc2275 (
      {stage1_63[42]},
      {stage2_63[27]}
   );
   gpc1_1 gpc2276 (
      {stage1_63[43]},
      {stage2_63[28]}
   );
   gpc1_1 gpc2277 (
      {stage1_63[44]},
      {stage2_63[29]}
   );
   gpc1_1 gpc2278 (
      {stage1_63[45]},
      {stage2_63[30]}
   );
   gpc1_1 gpc2279 (
      {stage1_63[46]},
      {stage2_63[31]}
   );
   gpc1_1 gpc2280 (
      {stage1_63[47]},
      {stage2_63[32]}
   );
   gpc1_1 gpc2281 (
      {stage1_63[48]},
      {stage2_63[33]}
   );
   gpc1_1 gpc2282 (
      {stage1_63[49]},
      {stage2_63[34]}
   );
   gpc1_1 gpc2283 (
      {stage1_63[50]},
      {stage2_63[35]}
   );
   gpc1_1 gpc2284 (
      {stage1_63[51]},
      {stage2_63[36]}
   );
   gpc1_1 gpc2285 (
      {stage1_63[52]},
      {stage2_63[37]}
   );
   gpc1_1 gpc2286 (
      {stage1_64[22]},
      {stage2_64[18]}
   );
   gpc1_1 gpc2287 (
      {stage1_64[23]},
      {stage2_64[19]}
   );
   gpc1_1 gpc2288 (
      {stage1_64[24]},
      {stage2_64[20]}
   );
   gpc1_1 gpc2289 (
      {stage1_64[25]},
      {stage2_64[21]}
   );
   gpc1_1 gpc2290 (
      {stage1_64[26]},
      {stage2_64[22]}
   );
   gpc1_1 gpc2291 (
      {stage1_64[27]},
      {stage2_64[23]}
   );
   gpc1_1 gpc2292 (
      {stage1_64[28]},
      {stage2_64[24]}
   );
   gpc1_1 gpc2293 (
      {stage1_64[29]},
      {stage2_64[25]}
   );
   gpc606_5 gpc2294 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4], stage2_0[5]},
      {stage2_2[0], stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5]},
      {stage3_4[0],stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc2295 (
      {stage2_0[6], stage2_0[7], stage2_0[8], stage2_0[9], stage2_0[10], stage2_0[11]},
      {stage2_2[6], stage2_2[7], stage2_2[8], stage2_2[9], stage2_2[10], stage2_2[11]},
      {stage3_4[1],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc606_5 gpc2296 (
      {stage2_0[12], stage2_0[13], stage2_0[14], stage2_0[15], stage2_0[16], stage2_0[17]},
      {stage2_2[12], stage2_2[13], stage2_2[14], stage2_2[15], stage2_2[16], stage2_2[17]},
      {stage3_4[2],stage3_3[2],stage3_2[2],stage3_1[2],stage3_0[2]}
   );
   gpc615_5 gpc2297 (
      {stage2_1[0], stage2_1[1], stage2_1[2], stage2_1[3], stage2_1[4]},
      {stage2_2[18]},
      {stage2_3[0], stage2_3[1], stage2_3[2], stage2_3[3], stage2_3[4], stage2_3[5]},
      {stage3_5[0],stage3_4[3],stage3_3[3],stage3_2[3],stage3_1[3]}
   );
   gpc615_5 gpc2298 (
      {stage2_1[5], stage2_1[6], stage2_1[7], stage2_1[8], stage2_1[9]},
      {stage2_2[19]},
      {stage2_3[6], stage2_3[7], stage2_3[8], stage2_3[9], stage2_3[10], stage2_3[11]},
      {stage3_5[1],stage3_4[4],stage3_3[4],stage3_2[4],stage3_1[4]}
   );
   gpc606_5 gpc2299 (
      {stage2_2[20], stage2_2[21], stage2_2[22], stage2_2[23], stage2_2[24], 1'b0},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3], stage2_4[4], stage2_4[5]},
      {stage3_6[0],stage3_5[2],stage3_4[5],stage3_3[5],stage3_2[5]}
   );
   gpc606_5 gpc2300 (
      {stage2_4[6], stage2_4[7], stage2_4[8], stage2_4[9], stage2_4[10], stage2_4[11]},
      {stage2_6[0], stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage3_8[0],stage3_7[0],stage3_6[1],stage3_5[3],stage3_4[6]}
   );
   gpc606_5 gpc2301 (
      {stage2_4[12], stage2_4[13], stage2_4[14], stage2_4[15], stage2_4[16], stage2_4[17]},
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10], stage2_6[11]},
      {stage3_8[1],stage3_7[1],stage3_6[2],stage3_5[4],stage3_4[7]}
   );
   gpc615_5 gpc2302 (
      {stage2_4[18], stage2_4[19], stage2_4[20], stage2_4[21], stage2_4[22]},
      {stage2_5[0]},
      {stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16], stage2_6[17]},
      {stage3_8[2],stage3_7[2],stage3_6[3],stage3_5[5],stage3_4[8]}
   );
   gpc606_5 gpc2303 (
      {stage2_5[1], stage2_5[2], stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6]},
      {stage2_7[0], stage2_7[1], stage2_7[2], stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage3_9[0],stage3_8[3],stage3_7[3],stage3_6[4],stage3_5[6]}
   );
   gpc606_5 gpc2304 (
      {stage2_5[7], stage2_5[8], stage2_5[9], stage2_5[10], stage2_5[11], stage2_5[12]},
      {stage2_7[6], stage2_7[7], stage2_7[8], stage2_7[9], stage2_7[10], stage2_7[11]},
      {stage3_9[1],stage3_8[4],stage3_7[4],stage3_6[5],stage3_5[7]}
   );
   gpc615_5 gpc2305 (
      {stage2_6[18], stage2_6[19], stage2_6[20], stage2_6[21], stage2_6[22]},
      {stage2_7[12]},
      {stage2_8[0], stage2_8[1], stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage3_10[0],stage3_9[2],stage3_8[5],stage3_7[5],stage3_6[6]}
   );
   gpc606_5 gpc2306 (
      {stage2_7[13], stage2_7[14], stage2_7[15], stage2_7[16], stage2_7[17], stage2_7[18]},
      {stage2_9[0], stage2_9[1], stage2_9[2], stage2_9[3], stage2_9[4], stage2_9[5]},
      {stage3_11[0],stage3_10[1],stage3_9[3],stage3_8[6],stage3_7[6]}
   );
   gpc606_5 gpc2307 (
      {stage2_7[19], stage2_7[20], stage2_7[21], stage2_7[22], stage2_7[23], stage2_7[24]},
      {stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9], stage2_9[10], stage2_9[11]},
      {stage3_11[1],stage3_10[2],stage3_9[4],stage3_8[7],stage3_7[7]}
   );
   gpc606_5 gpc2308 (
      {stage2_7[25], stage2_7[26], stage2_7[27], stage2_7[28], stage2_7[29], stage2_7[30]},
      {stage2_9[12], stage2_9[13], stage2_9[14], stage2_9[15], stage2_9[16], stage2_9[17]},
      {stage3_11[2],stage3_10[3],stage3_9[5],stage3_8[8],stage3_7[8]}
   );
   gpc606_5 gpc2309 (
      {stage2_7[31], stage2_7[32], stage2_7[33], stage2_7[34], stage2_7[35], stage2_7[36]},
      {stage2_9[18], stage2_9[19], stage2_9[20], stage2_9[21], stage2_9[22], stage2_9[23]},
      {stage3_11[3],stage3_10[4],stage3_9[6],stage3_8[9],stage3_7[9]}
   );
   gpc615_5 gpc2310 (
      {stage2_8[6], stage2_8[7], stage2_8[8], stage2_8[9], stage2_8[10]},
      {stage2_9[24]},
      {stage2_10[0], stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5]},
      {stage3_12[0],stage3_11[4],stage3_10[5],stage3_9[7],stage3_8[10]}
   );
   gpc615_5 gpc2311 (
      {stage2_8[11], stage2_8[12], stage2_8[13], stage2_8[14], stage2_8[15]},
      {stage2_9[25]},
      {stage2_10[6], stage2_10[7], stage2_10[8], stage2_10[9], stage2_10[10], stage2_10[11]},
      {stage3_12[1],stage3_11[5],stage3_10[6],stage3_9[8],stage3_8[11]}
   );
   gpc615_5 gpc2312 (
      {stage2_8[16], stage2_8[17], stage2_8[18], stage2_8[19], stage2_8[20]},
      {stage2_9[26]},
      {stage2_10[12], stage2_10[13], stage2_10[14], stage2_10[15], stage2_10[16], stage2_10[17]},
      {stage3_12[2],stage3_11[6],stage3_10[7],stage3_9[9],stage3_8[12]}
   );
   gpc615_5 gpc2313 (
      {stage2_8[21], stage2_8[22], stage2_8[23], stage2_8[24], stage2_8[25]},
      {stage2_9[27]},
      {stage2_10[18], stage2_10[19], stage2_10[20], stage2_10[21], stage2_10[22], stage2_10[23]},
      {stage3_12[3],stage3_11[7],stage3_10[8],stage3_9[10],stage3_8[13]}
   );
   gpc615_5 gpc2314 (
      {stage2_8[26], stage2_8[27], stage2_8[28], stage2_8[29], stage2_8[30]},
      {stage2_9[28]},
      {stage2_10[24], stage2_10[25], stage2_10[26], stage2_10[27], stage2_10[28], stage2_10[29]},
      {stage3_12[4],stage3_11[8],stage3_10[9],stage3_9[11],stage3_8[14]}
   );
   gpc606_5 gpc2315 (
      {stage2_9[29], stage2_9[30], stage2_9[31], stage2_9[32], stage2_9[33], stage2_9[34]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[5],stage3_11[9],stage3_10[10],stage3_9[12]}
   );
   gpc2116_5 gpc2316 (
      {stage2_11[6], stage2_11[7], stage2_11[8], stage2_11[9], stage2_11[10], stage2_11[11]},
      {stage2_12[0]},
      {stage2_13[0]},
      {stage2_14[0], stage2_14[1]},
      {stage3_15[0],stage3_14[0],stage3_13[1],stage3_12[6],stage3_11[10]}
   );
   gpc615_5 gpc2317 (
      {stage2_11[12], stage2_11[13], stage2_11[14], stage2_11[15], stage2_11[16]},
      {stage2_12[1]},
      {stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5], stage2_13[6]},
      {stage3_15[1],stage3_14[1],stage3_13[2],stage3_12[7],stage3_11[11]}
   );
   gpc615_5 gpc2318 (
      {stage2_11[17], stage2_11[18], stage2_11[19], stage2_11[20], stage2_11[21]},
      {stage2_12[2]},
      {stage2_13[7], stage2_13[8], stage2_13[9], stage2_13[10], stage2_13[11], stage2_13[12]},
      {stage3_15[2],stage3_14[2],stage3_13[3],stage3_12[8],stage3_11[12]}
   );
   gpc606_5 gpc2319 (
      {stage2_12[3], stage2_12[4], stage2_12[5], stage2_12[6], stage2_12[7], stage2_12[8]},
      {stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5], stage2_14[6], stage2_14[7]},
      {stage3_16[0],stage3_15[3],stage3_14[3],stage3_13[4],stage3_12[9]}
   );
   gpc606_5 gpc2320 (
      {stage2_12[9], stage2_12[10], stage2_12[11], stage2_12[12], stage2_12[13], stage2_12[14]},
      {stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11], stage2_14[12], stage2_14[13]},
      {stage3_16[1],stage3_15[4],stage3_14[4],stage3_13[5],stage3_12[10]}
   );
   gpc606_5 gpc2321 (
      {stage2_12[15], stage2_12[16], stage2_12[17], stage2_12[18], stage2_12[19], stage2_12[20]},
      {stage2_14[14], stage2_14[15], stage2_14[16], stage2_14[17], stage2_14[18], stage2_14[19]},
      {stage3_16[2],stage3_15[5],stage3_14[5],stage3_13[6],stage3_12[11]}
   );
   gpc606_5 gpc2322 (
      {stage2_12[21], stage2_12[22], stage2_12[23], stage2_12[24], stage2_12[25], stage2_12[26]},
      {stage2_14[20], stage2_14[21], stage2_14[22], stage2_14[23], stage2_14[24], stage2_14[25]},
      {stage3_16[3],stage3_15[6],stage3_14[6],stage3_13[7],stage3_12[12]}
   );
   gpc606_5 gpc2323 (
      {stage2_14[26], stage2_14[27], stage2_14[28], stage2_14[29], stage2_14[30], stage2_14[31]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[4],stage3_15[7],stage3_14[7]}
   );
   gpc615_5 gpc2324 (
      {stage2_14[32], stage2_14[33], stage2_14[34], stage2_14[35], stage2_14[36]},
      {stage2_15[0]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[1],stage3_16[5],stage3_15[8],stage3_14[8]}
   );
   gpc615_5 gpc2325 (
      {stage2_14[37], stage2_14[38], 1'b0, 1'b0, 1'b0},
      {stage2_15[1]},
      {stage2_16[12], stage2_16[13], stage2_16[14], stage2_16[15], stage2_16[16], stage2_16[17]},
      {stage3_18[2],stage3_17[2],stage3_16[6],stage3_15[9],stage3_14[9]}
   );
   gpc2135_5 gpc2326 (
      {stage2_15[2], stage2_15[3], stage2_15[4], stage2_15[5], stage2_15[6]},
      {stage2_16[18], stage2_16[19], stage2_16[20]},
      {stage2_17[0]},
      {stage2_18[0], stage2_18[1]},
      {stage3_19[0],stage3_18[3],stage3_17[3],stage3_16[7],stage3_15[10]}
   );
   gpc606_5 gpc2327 (
      {stage2_15[7], stage2_15[8], stage2_15[9], stage2_15[10], stage2_15[11], stage2_15[12]},
      {stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5], stage2_17[6]},
      {stage3_19[1],stage3_18[4],stage3_17[4],stage3_16[8],stage3_15[11]}
   );
   gpc615_5 gpc2328 (
      {stage2_15[13], stage2_15[14], stage2_15[15], stage2_15[16], stage2_15[17]},
      {stage2_16[21]},
      {stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11], stage2_17[12]},
      {stage3_19[2],stage3_18[5],stage3_17[5],stage3_16[9],stage3_15[12]}
   );
   gpc1163_5 gpc2329 (
      {stage2_17[13], stage2_17[14], stage2_17[15]},
      {stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5], stage2_18[6], stage2_18[7]},
      {stage2_19[0]},
      {stage2_20[0]},
      {stage3_21[0],stage3_20[0],stage3_19[3],stage3_18[6],stage3_17[6]}
   );
   gpc1163_5 gpc2330 (
      {stage2_17[16], stage2_17[17], stage2_17[18]},
      {stage2_18[8], stage2_18[9], stage2_18[10], stage2_18[11], stage2_18[12], stage2_18[13]},
      {stage2_19[1]},
      {stage2_20[1]},
      {stage3_21[1],stage3_20[1],stage3_19[4],stage3_18[7],stage3_17[7]}
   );
   gpc1163_5 gpc2331 (
      {stage2_17[19], stage2_17[20], stage2_17[21]},
      {stage2_18[14], stage2_18[15], stage2_18[16], stage2_18[17], stage2_18[18], stage2_18[19]},
      {stage2_19[2]},
      {stage2_20[2]},
      {stage3_21[2],stage3_20[2],stage3_19[5],stage3_18[8],stage3_17[8]}
   );
   gpc606_5 gpc2332 (
      {stage2_17[22], stage2_17[23], stage2_17[24], stage2_17[25], stage2_17[26], stage2_17[27]},
      {stage2_19[3], stage2_19[4], stage2_19[5], stage2_19[6], stage2_19[7], stage2_19[8]},
      {stage3_21[3],stage3_20[3],stage3_19[6],stage3_18[9],stage3_17[9]}
   );
   gpc615_5 gpc2333 (
      {stage2_17[28], stage2_17[29], stage2_17[30], stage2_17[31], stage2_17[32]},
      {stage2_18[20]},
      {stage2_19[9], stage2_19[10], stage2_19[11], stage2_19[12], stage2_19[13], stage2_19[14]},
      {stage3_21[4],stage3_20[4],stage3_19[7],stage3_18[10],stage3_17[10]}
   );
   gpc2135_5 gpc2334 (
      {stage2_18[21], stage2_18[22], stage2_18[23], stage2_18[24], stage2_18[25]},
      {stage2_19[15], stage2_19[16], stage2_19[17]},
      {stage2_20[3]},
      {stage2_21[0], stage2_21[1]},
      {stage3_22[0],stage3_21[5],stage3_20[5],stage3_19[8],stage3_18[11]}
   );
   gpc2135_5 gpc2335 (
      {stage2_18[26], stage2_18[27], stage2_18[28], stage2_18[29], stage2_18[30]},
      {stage2_19[18], stage2_19[19], stage2_19[20]},
      {stage2_20[4]},
      {stage2_21[2], stage2_21[3]},
      {stage3_22[1],stage3_21[6],stage3_20[6],stage3_19[9],stage3_18[12]}
   );
   gpc1343_5 gpc2336 (
      {stage2_20[5], stage2_20[6], stage2_20[7]},
      {stage2_21[4], stage2_21[5], stage2_21[6], stage2_21[7]},
      {stage2_22[0], stage2_22[1], stage2_22[2]},
      {stage2_23[0]},
      {stage3_24[0],stage3_23[0],stage3_22[2],stage3_21[7],stage3_20[7]}
   );
   gpc1343_5 gpc2337 (
      {stage2_20[8], stage2_20[9], stage2_20[10]},
      {stage2_21[8], stage2_21[9], stage2_21[10], stage2_21[11]},
      {stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage2_23[1]},
      {stage3_24[1],stage3_23[1],stage3_22[3],stage3_21[8],stage3_20[8]}
   );
   gpc615_5 gpc2338 (
      {stage2_20[11], stage2_20[12], stage2_20[13], stage2_20[14], stage2_20[15]},
      {stage2_21[12]},
      {stage2_22[6], stage2_22[7], stage2_22[8], stage2_22[9], stage2_22[10], stage2_22[11]},
      {stage3_24[2],stage3_23[2],stage3_22[4],stage3_21[9],stage3_20[9]}
   );
   gpc615_5 gpc2339 (
      {stage2_20[16], stage2_20[17], stage2_20[18], stage2_20[19], stage2_20[20]},
      {stage2_21[13]},
      {stage2_22[12], stage2_22[13], stage2_22[14], stage2_22[15], stage2_22[16], stage2_22[17]},
      {stage3_24[3],stage3_23[3],stage3_22[5],stage3_21[10],stage3_20[10]}
   );
   gpc615_5 gpc2340 (
      {stage2_20[21], stage2_20[22], stage2_20[23], stage2_20[24], stage2_20[25]},
      {stage2_21[14]},
      {stage2_22[18], stage2_22[19], stage2_22[20], stage2_22[21], stage2_22[22], stage2_22[23]},
      {stage3_24[4],stage3_23[4],stage3_22[6],stage3_21[11],stage3_20[11]}
   );
   gpc615_5 gpc2341 (
      {stage2_20[26], stage2_20[27], stage2_20[28], stage2_20[29], stage2_20[30]},
      {stage2_21[15]},
      {stage2_22[24], stage2_22[25], stage2_22[26], stage2_22[27], stage2_22[28], stage2_22[29]},
      {stage3_24[5],stage3_23[5],stage3_22[7],stage3_21[12],stage3_20[12]}
   );
   gpc623_5 gpc2342 (
      {stage2_20[31], stage2_20[32], stage2_20[33]},
      {stage2_21[16], stage2_21[17]},
      {stage2_22[30], stage2_22[31], stage2_22[32], stage2_22[33], stage2_22[34], 1'b0},
      {stage3_24[6],stage3_23[6],stage3_22[8],stage3_21[13],stage3_20[13]}
   );
   gpc2135_5 gpc2343 (
      {stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5], stage2_23[6]},
      {stage2_24[0], stage2_24[1], stage2_24[2]},
      {stage2_25[0]},
      {stage2_26[0], stage2_26[1]},
      {stage3_27[0],stage3_26[0],stage3_25[0],stage3_24[7],stage3_23[7]}
   );
   gpc2135_5 gpc2344 (
      {stage2_23[7], stage2_23[8], stage2_23[9], stage2_23[10], stage2_23[11]},
      {stage2_24[3], stage2_24[4], stage2_24[5]},
      {stage2_25[1]},
      {stage2_26[2], stage2_26[3]},
      {stage3_27[1],stage3_26[1],stage3_25[1],stage3_24[8],stage3_23[8]}
   );
   gpc615_5 gpc2345 (
      {stage2_23[12], stage2_23[13], stage2_23[14], stage2_23[15], stage2_23[16]},
      {stage2_24[6]},
      {stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5], stage2_25[6], stage2_25[7]},
      {stage3_27[2],stage3_26[2],stage3_25[2],stage3_24[9],stage3_23[9]}
   );
   gpc615_5 gpc2346 (
      {stage2_23[17], stage2_23[18], stage2_23[19], stage2_23[20], stage2_23[21]},
      {stage2_24[7]},
      {stage2_25[8], stage2_25[9], stage2_25[10], stage2_25[11], stage2_25[12], stage2_25[13]},
      {stage3_27[3],stage3_26[3],stage3_25[3],stage3_24[10],stage3_23[10]}
   );
   gpc615_5 gpc2347 (
      {stage2_23[22], stage2_23[23], stage2_23[24], stage2_23[25], stage2_23[26]},
      {stage2_24[8]},
      {stage2_25[14], stage2_25[15], stage2_25[16], stage2_25[17], stage2_25[18], stage2_25[19]},
      {stage3_27[4],stage3_26[4],stage3_25[4],stage3_24[11],stage3_23[11]}
   );
   gpc606_5 gpc2348 (
      {stage2_24[9], stage2_24[10], stage2_24[11], stage2_24[12], stage2_24[13], stage2_24[14]},
      {stage2_26[4], stage2_26[5], stage2_26[6], stage2_26[7], stage2_26[8], stage2_26[9]},
      {stage3_28[0],stage3_27[5],stage3_26[5],stage3_25[5],stage3_24[12]}
   );
   gpc606_5 gpc2349 (
      {stage2_24[15], stage2_24[16], stage2_24[17], stage2_24[18], stage2_24[19], stage2_24[20]},
      {stage2_26[10], stage2_26[11], stage2_26[12], stage2_26[13], stage2_26[14], stage2_26[15]},
      {stage3_28[1],stage3_27[6],stage3_26[6],stage3_25[6],stage3_24[13]}
   );
   gpc606_5 gpc2350 (
      {stage2_24[21], stage2_24[22], stage2_24[23], stage2_24[24], stage2_24[25], stage2_24[26]},
      {stage2_26[16], stage2_26[17], stage2_26[18], stage2_26[19], stage2_26[20], stage2_26[21]},
      {stage3_28[2],stage3_27[7],stage3_26[7],stage3_25[7],stage3_24[14]}
   );
   gpc2135_5 gpc2351 (
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4]},
      {stage2_28[0], stage2_28[1], stage2_28[2]},
      {stage2_29[0]},
      {stage2_30[0], stage2_30[1]},
      {stage3_31[0],stage3_30[0],stage3_29[0],stage3_28[3],stage3_27[8]}
   );
   gpc2135_5 gpc2352 (
      {stage2_27[5], stage2_27[6], stage2_27[7], stage2_27[8], stage2_27[9]},
      {stage2_28[3], stage2_28[4], stage2_28[5]},
      {stage2_29[1]},
      {stage2_30[2], stage2_30[3]},
      {stage3_31[1],stage3_30[1],stage3_29[1],stage3_28[4],stage3_27[9]}
   );
   gpc2135_5 gpc2353 (
      {stage2_27[10], stage2_27[11], stage2_27[12], stage2_27[13], stage2_27[14]},
      {stage2_28[6], stage2_28[7], stage2_28[8]},
      {stage2_29[2]},
      {stage2_30[4], stage2_30[5]},
      {stage3_31[2],stage3_30[2],stage3_29[2],stage3_28[5],stage3_27[10]}
   );
   gpc606_5 gpc2354 (
      {stage2_27[15], stage2_27[16], stage2_27[17], stage2_27[18], stage2_27[19], stage2_27[20]},
      {stage2_29[3], stage2_29[4], stage2_29[5], stage2_29[6], stage2_29[7], stage2_29[8]},
      {stage3_31[3],stage3_30[3],stage3_29[3],stage3_28[6],stage3_27[11]}
   );
   gpc606_5 gpc2355 (
      {stage2_27[21], stage2_27[22], stage2_27[23], stage2_27[24], stage2_27[25], stage2_27[26]},
      {stage2_29[9], stage2_29[10], stage2_29[11], stage2_29[12], stage2_29[13], stage2_29[14]},
      {stage3_31[4],stage3_30[4],stage3_29[4],stage3_28[7],stage3_27[12]}
   );
   gpc606_5 gpc2356 (
      {stage2_27[27], stage2_27[28], stage2_27[29], stage2_27[30], stage2_27[31], stage2_27[32]},
      {stage2_29[15], stage2_29[16], stage2_29[17], stage2_29[18], stage2_29[19], stage2_29[20]},
      {stage3_31[5],stage3_30[5],stage3_29[5],stage3_28[8],stage3_27[13]}
   );
   gpc606_5 gpc2357 (
      {stage2_28[9], stage2_28[10], stage2_28[11], stage2_28[12], stage2_28[13], stage2_28[14]},
      {stage2_30[6], stage2_30[7], stage2_30[8], stage2_30[9], stage2_30[10], stage2_30[11]},
      {stage3_32[0],stage3_31[6],stage3_30[6],stage3_29[6],stage3_28[9]}
   );
   gpc606_5 gpc2358 (
      {stage2_28[15], stage2_28[16], stage2_28[17], stage2_28[18], stage2_28[19], stage2_28[20]},
      {stage2_30[12], stage2_30[13], stage2_30[14], stage2_30[15], stage2_30[16], stage2_30[17]},
      {stage3_32[1],stage3_31[7],stage3_30[7],stage3_29[7],stage3_28[10]}
   );
   gpc2135_5 gpc2359 (
      {stage2_30[18], stage2_30[19], stage2_30[20], stage2_30[21], stage2_30[22]},
      {stage2_31[0], stage2_31[1], stage2_31[2]},
      {stage2_32[0]},
      {stage2_33[0], stage2_33[1]},
      {stage3_34[0],stage3_33[0],stage3_32[2],stage3_31[8],stage3_30[8]}
   );
   gpc2135_5 gpc2360 (
      {stage2_30[23], stage2_30[24], stage2_30[25], stage2_30[26], stage2_30[27]},
      {stage2_31[3], stage2_31[4], stage2_31[5]},
      {stage2_32[1]},
      {stage2_33[2], stage2_33[3]},
      {stage3_34[1],stage3_33[1],stage3_32[3],stage3_31[9],stage3_30[9]}
   );
   gpc2135_5 gpc2361 (
      {stage2_30[28], stage2_30[29], stage2_30[30], stage2_30[31], stage2_30[32]},
      {stage2_31[6], stage2_31[7], stage2_31[8]},
      {stage2_32[2]},
      {stage2_33[4], stage2_33[5]},
      {stage3_34[2],stage3_33[2],stage3_32[4],stage3_31[10],stage3_30[10]}
   );
   gpc2135_5 gpc2362 (
      {stage2_30[33], stage2_30[34], stage2_30[35], stage2_30[36], stage2_30[37]},
      {stage2_31[9], stage2_31[10], stage2_31[11]},
      {stage2_32[3]},
      {stage2_33[6], stage2_33[7]},
      {stage3_34[3],stage3_33[3],stage3_32[5],stage3_31[11],stage3_30[11]}
   );
   gpc2135_5 gpc2363 (
      {stage2_30[38], stage2_30[39], stage2_30[40], stage2_30[41], stage2_30[42]},
      {stage2_31[12], stage2_31[13], stage2_31[14]},
      {stage2_32[4]},
      {stage2_33[8], stage2_33[9]},
      {stage3_34[4],stage3_33[4],stage3_32[6],stage3_31[12],stage3_30[12]}
   );
   gpc615_5 gpc2364 (
      {stage2_30[43], stage2_30[44], stage2_30[45], stage2_30[46], stage2_30[47]},
      {stage2_31[15]},
      {stage2_32[5], stage2_32[6], stage2_32[7], stage2_32[8], stage2_32[9], stage2_32[10]},
      {stage3_34[5],stage3_33[5],stage3_32[7],stage3_31[13],stage3_30[13]}
   );
   gpc615_5 gpc2365 (
      {stage2_30[48], stage2_30[49], stage2_30[50], stage2_30[51], 1'b0},
      {stage2_31[16]},
      {stage2_32[11], stage2_32[12], stage2_32[13], stage2_32[14], stage2_32[15], stage2_32[16]},
      {stage3_34[6],stage3_33[6],stage3_32[8],stage3_31[14],stage3_30[14]}
   );
   gpc117_4 gpc2366 (
      {stage2_31[17], stage2_31[18], stage2_31[19], stage2_31[20], stage2_31[21], stage2_31[22], stage2_31[23]},
      {stage2_32[17]},
      {stage2_33[10]},
      {stage3_34[7],stage3_33[7],stage3_32[9],stage3_31[15]}
   );
   gpc606_5 gpc2367 (
      {stage2_32[18], stage2_32[19], stage2_32[20], stage2_32[21], stage2_32[22], stage2_32[23]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[0],stage3_34[8],stage3_33[8],stage3_32[10]}
   );
   gpc606_5 gpc2368 (
      {stage2_33[11], stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[1],stage3_35[1],stage3_34[9],stage3_33[9]}
   );
   gpc606_5 gpc2369 (
      {stage2_33[17], stage2_33[18], stage2_33[19], stage2_33[20], stage2_33[21], stage2_33[22]},
      {stage2_35[6], stage2_35[7], stage2_35[8], stage2_35[9], stage2_35[10], stage2_35[11]},
      {stage3_37[1],stage3_36[2],stage3_35[2],stage3_34[10],stage3_33[10]}
   );
   gpc606_5 gpc2370 (
      {stage2_33[23], stage2_33[24], stage2_33[25], stage2_33[26], stage2_33[27], stage2_33[28]},
      {stage2_35[12], stage2_35[13], stage2_35[14], stage2_35[15], stage2_35[16], stage2_35[17]},
      {stage3_37[2],stage3_36[3],stage3_35[3],stage3_34[11],stage3_33[11]}
   );
   gpc135_4 gpc2371 (
      {stage2_34[6], stage2_34[7], stage2_34[8], stage2_34[9], stage2_34[10]},
      {stage2_35[18], stage2_35[19], stage2_35[20]},
      {stage2_36[0]},
      {stage3_37[3],stage3_36[4],stage3_35[4],stage3_34[12]}
   );
   gpc135_4 gpc2372 (
      {stage2_34[11], stage2_34[12], stage2_34[13], stage2_34[14], stage2_34[15]},
      {stage2_35[21], stage2_35[22], stage2_35[23]},
      {stage2_36[1]},
      {stage3_37[4],stage3_36[5],stage3_35[5],stage3_34[13]}
   );
   gpc135_4 gpc2373 (
      {stage2_34[16], stage2_34[17], stage2_34[18], stage2_34[19], stage2_34[20]},
      {stage2_35[24], stage2_35[25], stage2_35[26]},
      {stage2_36[2]},
      {stage3_37[5],stage3_36[6],stage3_35[6],stage3_34[14]}
   );
   gpc615_5 gpc2374 (
      {stage2_34[21], stage2_34[22], stage2_34[23], stage2_34[24], stage2_34[25]},
      {stage2_35[27]},
      {stage2_36[3], stage2_36[4], stage2_36[5], stage2_36[6], stage2_36[7], stage2_36[8]},
      {stage3_38[0],stage3_37[6],stage3_36[7],stage3_35[7],stage3_34[15]}
   );
   gpc615_5 gpc2375 (
      {stage2_34[26], stage2_34[27], stage2_34[28], stage2_34[29], stage2_34[30]},
      {stage2_35[28]},
      {stage2_36[9], stage2_36[10], stage2_36[11], stage2_36[12], stage2_36[13], stage2_36[14]},
      {stage3_38[1],stage3_37[7],stage3_36[8],stage3_35[8],stage3_34[16]}
   );
   gpc1163_5 gpc2376 (
      {stage2_36[15], stage2_36[16], stage2_36[17]},
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5]},
      {stage2_38[0]},
      {stage2_39[0]},
      {stage3_40[0],stage3_39[0],stage3_38[2],stage3_37[8],stage3_36[9]}
   );
   gpc1163_5 gpc2377 (
      {stage2_36[18], stage2_36[19], stage2_36[20]},
      {stage2_37[6], stage2_37[7], stage2_37[8], stage2_37[9], stage2_37[10], stage2_37[11]},
      {stage2_38[1]},
      {stage2_39[1]},
      {stage3_40[1],stage3_39[1],stage3_38[3],stage3_37[9],stage3_36[10]}
   );
   gpc1163_5 gpc2378 (
      {stage2_36[21], stage2_36[22], stage2_36[23]},
      {stage2_37[12], stage2_37[13], stage2_37[14], stage2_37[15], stage2_37[16], stage2_37[17]},
      {stage2_38[2]},
      {stage2_39[2]},
      {stage3_40[2],stage3_39[2],stage3_38[4],stage3_37[10],stage3_36[11]}
   );
   gpc1163_5 gpc2379 (
      {stage2_36[24], stage2_36[25], stage2_36[26]},
      {stage2_37[18], stage2_37[19], stage2_37[20], stage2_37[21], stage2_37[22], stage2_37[23]},
      {stage2_38[3]},
      {stage2_39[3]},
      {stage3_40[3],stage3_39[3],stage3_38[5],stage3_37[11],stage3_36[12]}
   );
   gpc1163_5 gpc2380 (
      {stage2_36[27], stage2_36[28], stage2_36[29]},
      {stage2_37[24], stage2_37[25], stage2_37[26], stage2_37[27], stage2_37[28], stage2_37[29]},
      {stage2_38[4]},
      {stage2_39[4]},
      {stage3_40[4],stage3_39[4],stage3_38[6],stage3_37[12],stage3_36[13]}
   );
   gpc1163_5 gpc2381 (
      {stage2_36[30], stage2_36[31], stage2_36[32]},
      {stage2_37[30], stage2_37[31], stage2_37[32], stage2_37[33], stage2_37[34], stage2_37[35]},
      {stage2_38[5]},
      {stage2_39[5]},
      {stage3_40[5],stage3_39[5],stage3_38[7],stage3_37[13],stage3_36[14]}
   );
   gpc606_5 gpc2382 (
      {stage2_38[6], stage2_38[7], stage2_38[8], stage2_38[9], stage2_38[10], stage2_38[11]},
      {stage2_40[0], stage2_40[1], stage2_40[2], stage2_40[3], stage2_40[4], stage2_40[5]},
      {stage3_42[0],stage3_41[0],stage3_40[6],stage3_39[6],stage3_38[8]}
   );
   gpc606_5 gpc2383 (
      {stage2_38[12], stage2_38[13], stage2_38[14], stage2_38[15], stage2_38[16], stage2_38[17]},
      {stage2_40[6], stage2_40[7], stage2_40[8], stage2_40[9], stage2_40[10], stage2_40[11]},
      {stage3_42[1],stage3_41[1],stage3_40[7],stage3_39[7],stage3_38[9]}
   );
   gpc606_5 gpc2384 (
      {stage2_38[18], stage2_38[19], stage2_38[20], stage2_38[21], stage2_38[22], stage2_38[23]},
      {stage2_40[12], stage2_40[13], stage2_40[14], stage2_40[15], stage2_40[16], stage2_40[17]},
      {stage3_42[2],stage3_41[2],stage3_40[8],stage3_39[8],stage3_38[10]}
   );
   gpc606_5 gpc2385 (
      {stage2_38[24], stage2_38[25], stage2_38[26], stage2_38[27], stage2_38[28], stage2_38[29]},
      {stage2_40[18], stage2_40[19], stage2_40[20], stage2_40[21], stage2_40[22], stage2_40[23]},
      {stage3_42[3],stage3_41[3],stage3_40[9],stage3_39[9],stage3_38[11]}
   );
   gpc606_5 gpc2386 (
      {stage2_38[30], stage2_38[31], stage2_38[32], stage2_38[33], stage2_38[34], stage2_38[35]},
      {stage2_40[24], stage2_40[25], stage2_40[26], stage2_40[27], stage2_40[28], stage2_40[29]},
      {stage3_42[4],stage3_41[4],stage3_40[10],stage3_39[10],stage3_38[12]}
   );
   gpc606_5 gpc2387 (
      {stage2_39[6], stage2_39[7], stage2_39[8], stage2_39[9], stage2_39[10], stage2_39[11]},
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4], stage2_41[5]},
      {stage3_43[0],stage3_42[5],stage3_41[5],stage3_40[11],stage3_39[11]}
   );
   gpc606_5 gpc2388 (
      {stage2_39[12], stage2_39[13], stage2_39[14], stage2_39[15], stage2_39[16], stage2_39[17]},
      {stage2_41[6], stage2_41[7], stage2_41[8], stage2_41[9], stage2_41[10], stage2_41[11]},
      {stage3_43[1],stage3_42[6],stage3_41[6],stage3_40[12],stage3_39[12]}
   );
   gpc615_5 gpc2389 (
      {stage2_39[18], stage2_39[19], stage2_39[20], stage2_39[21], 1'b0},
      {stage2_40[30]},
      {stage2_41[12], stage2_41[13], stage2_41[14], stage2_41[15], stage2_41[16], stage2_41[17]},
      {stage3_43[2],stage3_42[7],stage3_41[7],stage3_40[13],stage3_39[13]}
   );
   gpc606_5 gpc2390 (
      {stage2_41[18], stage2_41[19], stage2_41[20], stage2_41[21], stage2_41[22], stage2_41[23]},
      {stage2_43[0], stage2_43[1], stage2_43[2], stage2_43[3], stage2_43[4], stage2_43[5]},
      {stage3_45[0],stage3_44[0],stage3_43[3],stage3_42[8],stage3_41[8]}
   );
   gpc606_5 gpc2391 (
      {stage2_41[24], stage2_41[25], stage2_41[26], stage2_41[27], stage2_41[28], stage2_41[29]},
      {stage2_43[6], stage2_43[7], stage2_43[8], stage2_43[9], stage2_43[10], stage2_43[11]},
      {stage3_45[1],stage3_44[1],stage3_43[4],stage3_42[9],stage3_41[9]}
   );
   gpc615_5 gpc2392 (
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4]},
      {stage2_43[12]},
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5]},
      {stage3_46[0],stage3_45[2],stage3_44[2],stage3_43[5],stage3_42[10]}
   );
   gpc615_5 gpc2393 (
      {stage2_42[5], stage2_42[6], stage2_42[7], stage2_42[8], stage2_42[9]},
      {stage2_43[13]},
      {stage2_44[6], stage2_44[7], stage2_44[8], stage2_44[9], stage2_44[10], stage2_44[11]},
      {stage3_46[1],stage3_45[3],stage3_44[3],stage3_43[6],stage3_42[11]}
   );
   gpc615_5 gpc2394 (
      {stage2_43[14], stage2_43[15], stage2_43[16], stage2_43[17], stage2_43[18]},
      {stage2_44[12]},
      {stage2_45[0], stage2_45[1], stage2_45[2], stage2_45[3], stage2_45[4], stage2_45[5]},
      {stage3_47[0],stage3_46[2],stage3_45[4],stage3_44[4],stage3_43[7]}
   );
   gpc606_5 gpc2395 (
      {stage2_44[13], stage2_44[14], stage2_44[15], stage2_44[16], stage2_44[17], stage2_44[18]},
      {stage2_46[0], stage2_46[1], stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5]},
      {stage3_48[0],stage3_47[1],stage3_46[3],stage3_45[5],stage3_44[5]}
   );
   gpc606_5 gpc2396 (
      {stage2_44[19], stage2_44[20], stage2_44[21], stage2_44[22], stage2_44[23], stage2_44[24]},
      {stage2_46[6], stage2_46[7], stage2_46[8], stage2_46[9], stage2_46[10], stage2_46[11]},
      {stage3_48[1],stage3_47[2],stage3_46[4],stage3_45[6],stage3_44[6]}
   );
   gpc615_5 gpc2397 (
      {stage2_44[25], stage2_44[26], stage2_44[27], stage2_44[28], stage2_44[29]},
      {stage2_45[6]},
      {stage2_46[12], stage2_46[13], stage2_46[14], stage2_46[15], stage2_46[16], stage2_46[17]},
      {stage3_48[2],stage3_47[3],stage3_46[5],stage3_45[7],stage3_44[7]}
   );
   gpc606_5 gpc2398 (
      {stage2_45[7], stage2_45[8], stage2_45[9], stage2_45[10], stage2_45[11], stage2_45[12]},
      {stage2_47[0], stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage3_49[0],stage3_48[3],stage3_47[4],stage3_46[6],stage3_45[8]}
   );
   gpc615_5 gpc2399 (
      {stage2_45[13], stage2_45[14], stage2_45[15], stage2_45[16], stage2_45[17]},
      {stage2_46[18]},
      {stage2_47[6], stage2_47[7], stage2_47[8], stage2_47[9], stage2_47[10], stage2_47[11]},
      {stage3_49[1],stage3_48[4],stage3_47[5],stage3_46[7],stage3_45[9]}
   );
   gpc615_5 gpc2400 (
      {stage2_45[18], stage2_45[19], stage2_45[20], stage2_45[21], stage2_45[22]},
      {stage2_46[19]},
      {stage2_47[12], stage2_47[13], stage2_47[14], stage2_47[15], stage2_47[16], stage2_47[17]},
      {stage3_49[2],stage3_48[5],stage3_47[6],stage3_46[8],stage3_45[10]}
   );
   gpc615_5 gpc2401 (
      {stage2_45[23], stage2_45[24], stage2_45[25], stage2_45[26], stage2_45[27]},
      {stage2_46[20]},
      {stage2_47[18], stage2_47[19], stage2_47[20], stage2_47[21], stage2_47[22], stage2_47[23]},
      {stage3_49[3],stage3_48[6],stage3_47[7],stage3_46[9],stage3_45[11]}
   );
   gpc615_5 gpc2402 (
      {stage2_45[28], stage2_45[29], stage2_45[30], stage2_45[31], stage2_45[32]},
      {stage2_46[21]},
      {stage2_47[24], stage2_47[25], stage2_47[26], stage2_47[27], stage2_47[28], stage2_47[29]},
      {stage3_49[4],stage3_48[7],stage3_47[8],stage3_46[10],stage3_45[12]}
   );
   gpc615_5 gpc2403 (
      {stage2_47[30], stage2_47[31], stage2_47[32], stage2_47[33], stage2_47[34]},
      {stage2_48[0]},
      {stage2_49[0], stage2_49[1], stage2_49[2], stage2_49[3], stage2_49[4], stage2_49[5]},
      {stage3_51[0],stage3_50[0],stage3_49[5],stage3_48[8],stage3_47[9]}
   );
   gpc615_5 gpc2404 (
      {stage2_48[1], stage2_48[2], stage2_48[3], stage2_48[4], stage2_48[5]},
      {stage2_49[6]},
      {stage2_50[0], stage2_50[1], stage2_50[2], stage2_50[3], stage2_50[4], stage2_50[5]},
      {stage3_52[0],stage3_51[1],stage3_50[1],stage3_49[6],stage3_48[9]}
   );
   gpc615_5 gpc2405 (
      {stage2_48[6], stage2_48[7], stage2_48[8], stage2_48[9], stage2_48[10]},
      {stage2_49[7]},
      {stage2_50[6], stage2_50[7], stage2_50[8], stage2_50[9], stage2_50[10], stage2_50[11]},
      {stage3_52[1],stage3_51[2],stage3_50[2],stage3_49[7],stage3_48[10]}
   );
   gpc615_5 gpc2406 (
      {stage2_48[11], stage2_48[12], stage2_48[13], stage2_48[14], stage2_48[15]},
      {stage2_49[8]},
      {stage2_50[12], stage2_50[13], stage2_50[14], stage2_50[15], stage2_50[16], stage2_50[17]},
      {stage3_52[2],stage3_51[3],stage3_50[3],stage3_49[8],stage3_48[11]}
   );
   gpc615_5 gpc2407 (
      {stage2_48[16], stage2_48[17], stage2_48[18], stage2_48[19], stage2_48[20]},
      {stage2_49[9]},
      {stage2_50[18], stage2_50[19], stage2_50[20], stage2_50[21], stage2_50[22], stage2_50[23]},
      {stage3_52[3],stage3_51[4],stage3_50[4],stage3_49[9],stage3_48[12]}
   );
   gpc615_5 gpc2408 (
      {stage2_48[21], stage2_48[22], stage2_48[23], stage2_48[24], stage2_48[25]},
      {stage2_49[10]},
      {stage2_50[24], stage2_50[25], stage2_50[26], stage2_50[27], stage2_50[28], stage2_50[29]},
      {stage3_52[4],stage3_51[5],stage3_50[5],stage3_49[10],stage3_48[13]}
   );
   gpc135_4 gpc2409 (
      {stage2_49[11], stage2_49[12], stage2_49[13], stage2_49[14], stage2_49[15]},
      {stage2_50[30], stage2_50[31], stage2_50[32]},
      {stage2_51[0]},
      {stage3_52[5],stage3_51[6],stage3_50[6],stage3_49[11]}
   );
   gpc615_5 gpc2410 (
      {stage2_51[1], stage2_51[2], stage2_51[3], stage2_51[4], stage2_51[5]},
      {stage2_52[0]},
      {stage2_53[0], stage2_53[1], stage2_53[2], stage2_53[3], stage2_53[4], stage2_53[5]},
      {stage3_55[0],stage3_54[0],stage3_53[0],stage3_52[6],stage3_51[7]}
   );
   gpc615_5 gpc2411 (
      {stage2_51[6], stage2_51[7], stage2_51[8], stage2_51[9], stage2_51[10]},
      {stage2_52[1]},
      {stage2_53[6], stage2_53[7], stage2_53[8], stage2_53[9], stage2_53[10], stage2_53[11]},
      {stage3_55[1],stage3_54[1],stage3_53[1],stage3_52[7],stage3_51[8]}
   );
   gpc615_5 gpc2412 (
      {stage2_51[11], stage2_51[12], stage2_51[13], stage2_51[14], stage2_51[15]},
      {stage2_52[2]},
      {stage2_53[12], stage2_53[13], stage2_53[14], stage2_53[15], stage2_53[16], stage2_53[17]},
      {stage3_55[2],stage3_54[2],stage3_53[2],stage3_52[8],stage3_51[9]}
   );
   gpc615_5 gpc2413 (
      {stage2_51[16], stage2_51[17], stage2_51[18], stage2_51[19], stage2_51[20]},
      {stage2_52[3]},
      {stage2_53[18], stage2_53[19], stage2_53[20], stage2_53[21], stage2_53[22], stage2_53[23]},
      {stage3_55[3],stage3_54[3],stage3_53[3],stage3_52[9],stage3_51[10]}
   );
   gpc615_5 gpc2414 (
      {stage2_51[21], stage2_51[22], stage2_51[23], stage2_51[24], stage2_51[25]},
      {stage2_52[4]},
      {stage2_53[24], stage2_53[25], stage2_53[26], stage2_53[27], stage2_53[28], stage2_53[29]},
      {stage3_55[4],stage3_54[4],stage3_53[4],stage3_52[10],stage3_51[11]}
   );
   gpc615_5 gpc2415 (
      {stage2_51[26], stage2_51[27], stage2_51[28], stage2_51[29], stage2_51[30]},
      {stage2_52[5]},
      {stage2_53[30], stage2_53[31], stage2_53[32], stage2_53[33], stage2_53[34], stage2_53[35]},
      {stage3_55[5],stage3_54[5],stage3_53[5],stage3_52[11],stage3_51[12]}
   );
   gpc615_5 gpc2416 (
      {stage2_52[6], stage2_52[7], stage2_52[8], stage2_52[9], stage2_52[10]},
      {stage2_53[36]},
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3], stage2_54[4], stage2_54[5]},
      {stage3_56[0],stage3_55[6],stage3_54[6],stage3_53[6],stage3_52[12]}
   );
   gpc1163_5 gpc2417 (
      {stage2_54[6], stage2_54[7], stage2_54[8]},
      {stage2_55[0], stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5]},
      {stage2_56[0]},
      {stage2_57[0]},
      {stage3_58[0],stage3_57[0],stage3_56[1],stage3_55[7],stage3_54[7]}
   );
   gpc1163_5 gpc2418 (
      {stage2_54[9], stage2_54[10], stage2_54[11]},
      {stage2_55[6], stage2_55[7], stage2_55[8], stage2_55[9], stage2_55[10], stage2_55[11]},
      {stage2_56[1]},
      {stage2_57[1]},
      {stage3_58[1],stage3_57[1],stage3_56[2],stage3_55[8],stage3_54[8]}
   );
   gpc1163_5 gpc2419 (
      {stage2_54[12], stage2_54[13], stage2_54[14]},
      {stage2_55[12], stage2_55[13], stage2_55[14], stage2_55[15], stage2_55[16], stage2_55[17]},
      {stage2_56[2]},
      {stage2_57[2]},
      {stage3_58[2],stage3_57[2],stage3_56[3],stage3_55[9],stage3_54[9]}
   );
   gpc606_5 gpc2420 (
      {stage2_56[3], stage2_56[4], stage2_56[5], stage2_56[6], stage2_56[7], stage2_56[8]},
      {stage2_58[0], stage2_58[1], stage2_58[2], stage2_58[3], stage2_58[4], stage2_58[5]},
      {stage3_60[0],stage3_59[0],stage3_58[3],stage3_57[3],stage3_56[4]}
   );
   gpc606_5 gpc2421 (
      {stage2_56[9], stage2_56[10], stage2_56[11], stage2_56[12], stage2_56[13], stage2_56[14]},
      {stage2_58[6], stage2_58[7], stage2_58[8], stage2_58[9], stage2_58[10], stage2_58[11]},
      {stage3_60[1],stage3_59[1],stage3_58[4],stage3_57[4],stage3_56[5]}
   );
   gpc606_5 gpc2422 (
      {stage2_56[15], stage2_56[16], stage2_56[17], stage2_56[18], stage2_56[19], stage2_56[20]},
      {stage2_58[12], stage2_58[13], stage2_58[14], stage2_58[15], stage2_58[16], stage2_58[17]},
      {stage3_60[2],stage3_59[2],stage3_58[5],stage3_57[5],stage3_56[6]}
   );
   gpc606_5 gpc2423 (
      {stage2_56[21], stage2_56[22], stage2_56[23], stage2_56[24], stage2_56[25], stage2_56[26]},
      {stage2_58[18], stage2_58[19], stage2_58[20], stage2_58[21], stage2_58[22], stage2_58[23]},
      {stage3_60[3],stage3_59[3],stage3_58[6],stage3_57[6],stage3_56[7]}
   );
   gpc606_5 gpc2424 (
      {stage2_57[3], stage2_57[4], stage2_57[5], stage2_57[6], stage2_57[7], stage2_57[8]},
      {stage2_59[0], stage2_59[1], stage2_59[2], stage2_59[3], stage2_59[4], stage2_59[5]},
      {stage3_61[0],stage3_60[4],stage3_59[4],stage3_58[7],stage3_57[7]}
   );
   gpc606_5 gpc2425 (
      {stage2_57[9], stage2_57[10], stage2_57[11], stage2_57[12], stage2_57[13], stage2_57[14]},
      {stage2_59[6], stage2_59[7], stage2_59[8], stage2_59[9], stage2_59[10], stage2_59[11]},
      {stage3_61[1],stage3_60[5],stage3_59[5],stage3_58[8],stage3_57[8]}
   );
   gpc606_5 gpc2426 (
      {stage2_57[15], stage2_57[16], stage2_57[17], stage2_57[18], stage2_57[19], stage2_57[20]},
      {stage2_59[12], stage2_59[13], stage2_59[14], stage2_59[15], stage2_59[16], stage2_59[17]},
      {stage3_61[2],stage3_60[6],stage3_59[6],stage3_58[9],stage3_57[9]}
   );
   gpc606_5 gpc2427 (
      {stage2_57[21], stage2_57[22], stage2_57[23], stage2_57[24], stage2_57[25], stage2_57[26]},
      {stage2_59[18], stage2_59[19], stage2_59[20], stage2_59[21], stage2_59[22], stage2_59[23]},
      {stage3_61[3],stage3_60[7],stage3_59[7],stage3_58[10],stage3_57[10]}
   );
   gpc606_5 gpc2428 (
      {stage2_57[27], stage2_57[28], stage2_57[29], stage2_57[30], stage2_57[31], stage2_57[32]},
      {stage2_59[24], stage2_59[25], stage2_59[26], stage2_59[27], stage2_59[28], stage2_59[29]},
      {stage3_61[4],stage3_60[8],stage3_59[8],stage3_58[11],stage3_57[11]}
   );
   gpc606_5 gpc2429 (
      {stage2_60[0], stage2_60[1], stage2_60[2], stage2_60[3], stage2_60[4], stage2_60[5]},
      {stage2_62[0], stage2_62[1], stage2_62[2], stage2_62[3], stage2_62[4], stage2_62[5]},
      {stage3_64[0],stage3_63[0],stage3_62[0],stage3_61[5],stage3_60[9]}
   );
   gpc606_5 gpc2430 (
      {stage2_60[6], stage2_60[7], stage2_60[8], stage2_60[9], stage2_60[10], stage2_60[11]},
      {stage2_62[6], stage2_62[7], stage2_62[8], stage2_62[9], stage2_62[10], stage2_62[11]},
      {stage3_64[1],stage3_63[1],stage3_62[1],stage3_61[6],stage3_60[10]}
   );
   gpc606_5 gpc2431 (
      {stage2_60[12], stage2_60[13], stage2_60[14], stage2_60[15], stage2_60[16], stage2_60[17]},
      {stage2_62[12], stage2_62[13], stage2_62[14], stage2_62[15], stage2_62[16], stage2_62[17]},
      {stage3_64[2],stage3_63[2],stage3_62[2],stage3_61[7],stage3_60[11]}
   );
   gpc623_5 gpc2432 (
      {stage2_60[18], stage2_60[19], stage2_60[20]},
      {stage2_61[0], stage2_61[1]},
      {stage2_62[18], stage2_62[19], stage2_62[20], stage2_62[21], stage2_62[22], stage2_62[23]},
      {stage3_64[3],stage3_63[3],stage3_62[3],stage3_61[8],stage3_60[12]}
   );
   gpc606_5 gpc2433 (
      {stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5], stage2_61[6], stage2_61[7]},
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5]},
      {stage3_65[0],stage3_64[4],stage3_63[4],stage3_62[4],stage3_61[9]}
   );
   gpc606_5 gpc2434 (
      {stage2_61[8], stage2_61[9], stage2_61[10], stage2_61[11], stage2_61[12], stage2_61[13]},
      {stage2_63[6], stage2_63[7], stage2_63[8], stage2_63[9], stage2_63[10], stage2_63[11]},
      {stage3_65[1],stage3_64[5],stage3_63[5],stage3_62[5],stage3_61[10]}
   );
   gpc606_5 gpc2435 (
      {stage2_61[14], stage2_61[15], stage2_61[16], stage2_61[17], stage2_61[18], stage2_61[19]},
      {stage2_63[12], stage2_63[13], stage2_63[14], stage2_63[15], stage2_63[16], stage2_63[17]},
      {stage3_65[2],stage3_64[6],stage3_63[6],stage3_62[6],stage3_61[11]}
   );
   gpc606_5 gpc2436 (
      {stage2_62[24], stage2_62[25], stage2_62[26], stage2_62[27], stage2_62[28], stage2_62[29]},
      {stage2_64[0], stage2_64[1], stage2_64[2], stage2_64[3], stage2_64[4], stage2_64[5]},
      {stage3_66[0],stage3_65[3],stage3_64[7],stage3_63[7],stage3_62[7]}
   );
   gpc1343_5 gpc2437 (
      {stage2_63[18], stage2_63[19], stage2_63[20]},
      {stage2_64[6], stage2_64[7], stage2_64[8], stage2_64[9]},
      {stage2_65[0], stage2_65[1], stage2_65[2]},
      {stage2_66[0]},
      {stage3_67[0],stage3_66[1],stage3_65[4],stage3_64[8],stage3_63[8]}
   );
   gpc1343_5 gpc2438 (
      {stage2_63[21], stage2_63[22], stage2_63[23]},
      {stage2_64[10], stage2_64[11], stage2_64[12], stage2_64[13]},
      {stage2_65[3], stage2_65[4], stage2_65[5]},
      {stage2_66[1]},
      {stage3_67[1],stage3_66[2],stage3_65[5],stage3_64[9],stage3_63[9]}
   );
   gpc1343_5 gpc2439 (
      {stage2_63[24], stage2_63[25], stage2_63[26]},
      {stage2_64[14], stage2_64[15], stage2_64[16], stage2_64[17]},
      {stage2_65[6], stage2_65[7], stage2_65[8]},
      {stage2_66[2]},
      {stage3_67[2],stage3_66[3],stage3_65[6],stage3_64[10],stage3_63[10]}
   );
   gpc1343_5 gpc2440 (
      {stage2_63[27], stage2_63[28], stage2_63[29]},
      {stage2_64[18], stage2_64[19], stage2_64[20], stage2_64[21]},
      {stage2_65[9], stage2_65[10], stage2_65[11]},
      {stage2_66[3]},
      {stage3_67[3],stage3_66[4],stage3_65[7],stage3_64[11],stage3_63[11]}
   );
   gpc1343_5 gpc2441 (
      {stage2_63[30], stage2_63[31], stage2_63[32]},
      {stage2_64[22], stage2_64[23], stage2_64[24], stage2_64[25]},
      {stage2_65[12], stage2_65[13], stage2_65[14]},
      {stage2_66[4]},
      {stage3_67[4],stage3_66[5],stage3_65[8],stage3_64[12],stage3_63[12]}
   );
   gpc1_1 gpc2442 (
      {stage2_0[18]},
      {stage3_0[3]}
   );
   gpc1_1 gpc2443 (
      {stage2_0[19]},
      {stage3_0[4]}
   );
   gpc1_1 gpc2444 (
      {stage2_1[10]},
      {stage3_1[5]}
   );
   gpc1_1 gpc2445 (
      {stage2_1[11]},
      {stage3_1[6]}
   );
   gpc1_1 gpc2446 (
      {stage2_1[12]},
      {stage3_1[7]}
   );
   gpc1_1 gpc2447 (
      {stage2_3[12]},
      {stage3_3[6]}
   );
   gpc1_1 gpc2448 (
      {stage2_3[13]},
      {stage3_3[7]}
   );
   gpc1_1 gpc2449 (
      {stage2_3[14]},
      {stage3_3[8]}
   );
   gpc1_1 gpc2450 (
      {stage2_3[15]},
      {stage3_3[9]}
   );
   gpc1_1 gpc2451 (
      {stage2_3[16]},
      {stage3_3[10]}
   );
   gpc1_1 gpc2452 (
      {stage2_3[17]},
      {stage3_3[11]}
   );
   gpc1_1 gpc2453 (
      {stage2_3[18]},
      {stage3_3[12]}
   );
   gpc1_1 gpc2454 (
      {stage2_3[19]},
      {stage3_3[13]}
   );
   gpc1_1 gpc2455 (
      {stage2_3[20]},
      {stage3_3[14]}
   );
   gpc1_1 gpc2456 (
      {stage2_3[21]},
      {stage3_3[15]}
   );
   gpc1_1 gpc2457 (
      {stage2_3[22]},
      {stage3_3[16]}
   );
   gpc1_1 gpc2458 (
      {stage2_3[23]},
      {stage3_3[17]}
   );
   gpc1_1 gpc2459 (
      {stage2_3[24]},
      {stage3_3[18]}
   );
   gpc1_1 gpc2460 (
      {stage2_3[25]},
      {stage3_3[19]}
   );
   gpc1_1 gpc2461 (
      {stage2_3[26]},
      {stage3_3[20]}
   );
   gpc1_1 gpc2462 (
      {stage2_3[27]},
      {stage3_3[21]}
   );
   gpc1_1 gpc2463 (
      {stage2_4[23]},
      {stage3_4[9]}
   );
   gpc1_1 gpc2464 (
      {stage2_4[24]},
      {stage3_4[10]}
   );
   gpc1_1 gpc2465 (
      {stage2_4[25]},
      {stage3_4[11]}
   );
   gpc1_1 gpc2466 (
      {stage2_5[13]},
      {stage3_5[8]}
   );
   gpc1_1 gpc2467 (
      {stage2_5[14]},
      {stage3_5[9]}
   );
   gpc1_1 gpc2468 (
      {stage2_5[15]},
      {stage3_5[10]}
   );
   gpc1_1 gpc2469 (
      {stage2_5[16]},
      {stage3_5[11]}
   );
   gpc1_1 gpc2470 (
      {stage2_5[17]},
      {stage3_5[12]}
   );
   gpc1_1 gpc2471 (
      {stage2_5[18]},
      {stage3_5[13]}
   );
   gpc1_1 gpc2472 (
      {stage2_5[19]},
      {stage3_5[14]}
   );
   gpc1_1 gpc2473 (
      {stage2_5[20]},
      {stage3_5[15]}
   );
   gpc1_1 gpc2474 (
      {stage2_5[21]},
      {stage3_5[16]}
   );
   gpc1_1 gpc2475 (
      {stage2_5[22]},
      {stage3_5[17]}
   );
   gpc1_1 gpc2476 (
      {stage2_5[23]},
      {stage3_5[18]}
   );
   gpc1_1 gpc2477 (
      {stage2_5[24]},
      {stage3_5[19]}
   );
   gpc1_1 gpc2478 (
      {stage2_5[25]},
      {stage3_5[20]}
   );
   gpc1_1 gpc2479 (
      {stage2_5[26]},
      {stage3_5[21]}
   );
   gpc1_1 gpc2480 (
      {stage2_5[27]},
      {stage3_5[22]}
   );
   gpc1_1 gpc2481 (
      {stage2_5[28]},
      {stage3_5[23]}
   );
   gpc1_1 gpc2482 (
      {stage2_6[23]},
      {stage3_6[7]}
   );
   gpc1_1 gpc2483 (
      {stage2_6[24]},
      {stage3_6[8]}
   );
   gpc1_1 gpc2484 (
      {stage2_6[25]},
      {stage3_6[9]}
   );
   gpc1_1 gpc2485 (
      {stage2_7[37]},
      {stage3_7[10]}
   );
   gpc1_1 gpc2486 (
      {stage2_7[38]},
      {stage3_7[11]}
   );
   gpc1_1 gpc2487 (
      {stage2_8[31]},
      {stage3_8[15]}
   );
   gpc1_1 gpc2488 (
      {stage2_9[35]},
      {stage3_9[13]}
   );
   gpc1_1 gpc2489 (
      {stage2_9[36]},
      {stage3_9[14]}
   );
   gpc1_1 gpc2490 (
      {stage2_9[37]},
      {stage3_9[15]}
   );
   gpc1_1 gpc2491 (
      {stage2_9[38]},
      {stage3_9[16]}
   );
   gpc1_1 gpc2492 (
      {stage2_9[39]},
      {stage3_9[17]}
   );
   gpc1_1 gpc2493 (
      {stage2_9[40]},
      {stage3_9[18]}
   );
   gpc1_1 gpc2494 (
      {stage2_9[41]},
      {stage3_9[19]}
   );
   gpc1_1 gpc2495 (
      {stage2_10[30]},
      {stage3_10[11]}
   );
   gpc1_1 gpc2496 (
      {stage2_12[27]},
      {stage3_12[13]}
   );
   gpc1_1 gpc2497 (
      {stage2_13[13]},
      {stage3_13[8]}
   );
   gpc1_1 gpc2498 (
      {stage2_13[14]},
      {stage3_13[9]}
   );
   gpc1_1 gpc2499 (
      {stage2_13[15]},
      {stage3_13[10]}
   );
   gpc1_1 gpc2500 (
      {stage2_13[16]},
      {stage3_13[11]}
   );
   gpc1_1 gpc2501 (
      {stage2_15[18]},
      {stage3_15[13]}
   );
   gpc1_1 gpc2502 (
      {stage2_15[19]},
      {stage3_15[14]}
   );
   gpc1_1 gpc2503 (
      {stage2_15[20]},
      {stage3_15[15]}
   );
   gpc1_1 gpc2504 (
      {stage2_15[21]},
      {stage3_15[16]}
   );
   gpc1_1 gpc2505 (
      {stage2_15[22]},
      {stage3_15[17]}
   );
   gpc1_1 gpc2506 (
      {stage2_15[23]},
      {stage3_15[18]}
   );
   gpc1_1 gpc2507 (
      {stage2_15[24]},
      {stage3_15[19]}
   );
   gpc1_1 gpc2508 (
      {stage2_15[25]},
      {stage3_15[20]}
   );
   gpc1_1 gpc2509 (
      {stage2_15[26]},
      {stage3_15[21]}
   );
   gpc1_1 gpc2510 (
      {stage2_15[27]},
      {stage3_15[22]}
   );
   gpc1_1 gpc2511 (
      {stage2_15[28]},
      {stage3_15[23]}
   );
   gpc1_1 gpc2512 (
      {stage2_15[29]},
      {stage3_15[24]}
   );
   gpc1_1 gpc2513 (
      {stage2_15[30]},
      {stage3_15[25]}
   );
   gpc1_1 gpc2514 (
      {stage2_16[22]},
      {stage3_16[10]}
   );
   gpc1_1 gpc2515 (
      {stage2_16[23]},
      {stage3_16[11]}
   );
   gpc1_1 gpc2516 (
      {stage2_17[33]},
      {stage3_17[11]}
   );
   gpc1_1 gpc2517 (
      {stage2_19[21]},
      {stage3_19[10]}
   );
   gpc1_1 gpc2518 (
      {stage2_19[22]},
      {stage3_19[11]}
   );
   gpc1_1 gpc2519 (
      {stage2_19[23]},
      {stage3_19[12]}
   );
   gpc1_1 gpc2520 (
      {stage2_19[24]},
      {stage3_19[13]}
   );
   gpc1_1 gpc2521 (
      {stage2_19[25]},
      {stage3_19[14]}
   );
   gpc1_1 gpc2522 (
      {stage2_19[26]},
      {stage3_19[15]}
   );
   gpc1_1 gpc2523 (
      {stage2_21[18]},
      {stage3_21[14]}
   );
   gpc1_1 gpc2524 (
      {stage2_21[19]},
      {stage3_21[15]}
   );
   gpc1_1 gpc2525 (
      {stage2_21[20]},
      {stage3_21[16]}
   );
   gpc1_1 gpc2526 (
      {stage2_21[21]},
      {stage3_21[17]}
   );
   gpc1_1 gpc2527 (
      {stage2_23[27]},
      {stage3_23[12]}
   );
   gpc1_1 gpc2528 (
      {stage2_24[27]},
      {stage3_24[15]}
   );
   gpc1_1 gpc2529 (
      {stage2_25[20]},
      {stage3_25[8]}
   );
   gpc1_1 gpc2530 (
      {stage2_25[21]},
      {stage3_25[9]}
   );
   gpc1_1 gpc2531 (
      {stage2_25[22]},
      {stage3_25[10]}
   );
   gpc1_1 gpc2532 (
      {stage2_25[23]},
      {stage3_25[11]}
   );
   gpc1_1 gpc2533 (
      {stage2_25[24]},
      {stage3_25[12]}
   );
   gpc1_1 gpc2534 (
      {stage2_25[25]},
      {stage3_25[13]}
   );
   gpc1_1 gpc2535 (
      {stage2_25[26]},
      {stage3_25[14]}
   );
   gpc1_1 gpc2536 (
      {stage2_25[27]},
      {stage3_25[15]}
   );
   gpc1_1 gpc2537 (
      {stage2_25[28]},
      {stage3_25[16]}
   );
   gpc1_1 gpc2538 (
      {stage2_25[29]},
      {stage3_25[17]}
   );
   gpc1_1 gpc2539 (
      {stage2_25[30]},
      {stage3_25[18]}
   );
   gpc1_1 gpc2540 (
      {stage2_25[31]},
      {stage3_25[19]}
   );
   gpc1_1 gpc2541 (
      {stage2_26[22]},
      {stage3_26[8]}
   );
   gpc1_1 gpc2542 (
      {stage2_26[23]},
      {stage3_26[9]}
   );
   gpc1_1 gpc2543 (
      {stage2_26[24]},
      {stage3_26[10]}
   );
   gpc1_1 gpc2544 (
      {stage2_26[25]},
      {stage3_26[11]}
   );
   gpc1_1 gpc2545 (
      {stage2_26[26]},
      {stage3_26[12]}
   );
   gpc1_1 gpc2546 (
      {stage2_28[21]},
      {stage3_28[11]}
   );
   gpc1_1 gpc2547 (
      {stage2_28[22]},
      {stage3_28[12]}
   );
   gpc1_1 gpc2548 (
      {stage2_28[23]},
      {stage3_28[13]}
   );
   gpc1_1 gpc2549 (
      {stage2_28[24]},
      {stage3_28[14]}
   );
   gpc1_1 gpc2550 (
      {stage2_28[25]},
      {stage3_28[15]}
   );
   gpc1_1 gpc2551 (
      {stage2_28[26]},
      {stage3_28[16]}
   );
   gpc1_1 gpc2552 (
      {stage2_31[24]},
      {stage3_31[16]}
   );
   gpc1_1 gpc2553 (
      {stage2_31[25]},
      {stage3_31[17]}
   );
   gpc1_1 gpc2554 (
      {stage2_31[26]},
      {stage3_31[18]}
   );
   gpc1_1 gpc2555 (
      {stage2_31[27]},
      {stage3_31[19]}
   );
   gpc1_1 gpc2556 (
      {stage2_32[24]},
      {stage3_32[11]}
   );
   gpc1_1 gpc2557 (
      {stage2_34[31]},
      {stage3_34[17]}
   );
   gpc1_1 gpc2558 (
      {stage2_35[29]},
      {stage3_35[9]}
   );
   gpc1_1 gpc2559 (
      {stage2_37[36]},
      {stage3_37[14]}
   );
   gpc1_1 gpc2560 (
      {stage2_40[31]},
      {stage3_40[14]}
   );
   gpc1_1 gpc2561 (
      {stage2_40[32]},
      {stage3_40[15]}
   );
   gpc1_1 gpc2562 (
      {stage2_40[33]},
      {stage3_40[16]}
   );
   gpc1_1 gpc2563 (
      {stage2_40[34]},
      {stage3_40[17]}
   );
   gpc1_1 gpc2564 (
      {stage2_41[30]},
      {stage3_41[10]}
   );
   gpc1_1 gpc2565 (
      {stage2_41[31]},
      {stage3_41[11]}
   );
   gpc1_1 gpc2566 (
      {stage2_42[10]},
      {stage3_42[12]}
   );
   gpc1_1 gpc2567 (
      {stage2_42[11]},
      {stage3_42[13]}
   );
   gpc1_1 gpc2568 (
      {stage2_42[12]},
      {stage3_42[14]}
   );
   gpc1_1 gpc2569 (
      {stage2_42[13]},
      {stage3_42[15]}
   );
   gpc1_1 gpc2570 (
      {stage2_42[14]},
      {stage3_42[16]}
   );
   gpc1_1 gpc2571 (
      {stage2_42[15]},
      {stage3_42[17]}
   );
   gpc1_1 gpc2572 (
      {stage2_42[16]},
      {stage3_42[18]}
   );
   gpc1_1 gpc2573 (
      {stage2_42[17]},
      {stage3_42[19]}
   );
   gpc1_1 gpc2574 (
      {stage2_43[19]},
      {stage3_43[8]}
   );
   gpc1_1 gpc2575 (
      {stage2_43[20]},
      {stage3_43[9]}
   );
   gpc1_1 gpc2576 (
      {stage2_45[33]},
      {stage3_45[13]}
   );
   gpc1_1 gpc2577 (
      {stage2_45[34]},
      {stage3_45[14]}
   );
   gpc1_1 gpc2578 (
      {stage2_46[22]},
      {stage3_46[11]}
   );
   gpc1_1 gpc2579 (
      {stage2_47[35]},
      {stage3_47[10]}
   );
   gpc1_1 gpc2580 (
      {stage2_48[26]},
      {stage3_48[14]}
   );
   gpc1_1 gpc2581 (
      {stage2_48[27]},
      {stage3_48[15]}
   );
   gpc1_1 gpc2582 (
      {stage2_48[28]},
      {stage3_48[16]}
   );
   gpc1_1 gpc2583 (
      {stage2_48[29]},
      {stage3_48[17]}
   );
   gpc1_1 gpc2584 (
      {stage2_48[30]},
      {stage3_48[18]}
   );
   gpc1_1 gpc2585 (
      {stage2_52[11]},
      {stage3_52[13]}
   );
   gpc1_1 gpc2586 (
      {stage2_52[12]},
      {stage3_52[14]}
   );
   gpc1_1 gpc2587 (
      {stage2_52[13]},
      {stage3_52[15]}
   );
   gpc1_1 gpc2588 (
      {stage2_52[14]},
      {stage3_52[16]}
   );
   gpc1_1 gpc2589 (
      {stage2_52[15]},
      {stage3_52[17]}
   );
   gpc1_1 gpc2590 (
      {stage2_52[16]},
      {stage3_52[18]}
   );
   gpc1_1 gpc2591 (
      {stage2_52[17]},
      {stage3_52[19]}
   );
   gpc1_1 gpc2592 (
      {stage2_53[37]},
      {stage3_53[7]}
   );
   gpc1_1 gpc2593 (
      {stage2_53[38]},
      {stage3_53[8]}
   );
   gpc1_1 gpc2594 (
      {stage2_54[15]},
      {stage3_54[10]}
   );
   gpc1_1 gpc2595 (
      {stage2_54[16]},
      {stage3_54[11]}
   );
   gpc1_1 gpc2596 (
      {stage2_54[17]},
      {stage3_54[12]}
   );
   gpc1_1 gpc2597 (
      {stage2_54[18]},
      {stage3_54[13]}
   );
   gpc1_1 gpc2598 (
      {stage2_54[19]},
      {stage3_54[14]}
   );
   gpc1_1 gpc2599 (
      {stage2_54[20]},
      {stage3_54[15]}
   );
   gpc1_1 gpc2600 (
      {stage2_54[21]},
      {stage3_54[16]}
   );
   gpc1_1 gpc2601 (
      {stage2_54[22]},
      {stage3_54[17]}
   );
   gpc1_1 gpc2602 (
      {stage2_54[23]},
      {stage3_54[18]}
   );
   gpc1_1 gpc2603 (
      {stage2_54[24]},
      {stage3_54[19]}
   );
   gpc1_1 gpc2604 (
      {stage2_54[25]},
      {stage3_54[20]}
   );
   gpc1_1 gpc2605 (
      {stage2_54[26]},
      {stage3_54[21]}
   );
   gpc1_1 gpc2606 (
      {stage2_54[27]},
      {stage3_54[22]}
   );
   gpc1_1 gpc2607 (
      {stage2_54[28]},
      {stage3_54[23]}
   );
   gpc1_1 gpc2608 (
      {stage2_55[18]},
      {stage3_55[10]}
   );
   gpc1_1 gpc2609 (
      {stage2_55[19]},
      {stage3_55[11]}
   );
   gpc1_1 gpc2610 (
      {stage2_59[30]},
      {stage3_59[9]}
   );
   gpc1_1 gpc2611 (
      {stage2_59[31]},
      {stage3_59[10]}
   );
   gpc1_1 gpc2612 (
      {stage2_59[32]},
      {stage3_59[11]}
   );
   gpc1_1 gpc2613 (
      {stage2_59[33]},
      {stage3_59[12]}
   );
   gpc1_1 gpc2614 (
      {stage2_59[34]},
      {stage3_59[13]}
   );
   gpc1_1 gpc2615 (
      {stage2_60[21]},
      {stage3_60[13]}
   );
   gpc1_1 gpc2616 (
      {stage2_61[20]},
      {stage3_61[12]}
   );
   gpc1_1 gpc2617 (
      {stage2_61[21]},
      {stage3_61[13]}
   );
   gpc1_1 gpc2618 (
      {stage2_61[22]},
      {stage3_61[14]}
   );
   gpc1_1 gpc2619 (
      {stage2_61[23]},
      {stage3_61[15]}
   );
   gpc1_1 gpc2620 (
      {stage2_61[24]},
      {stage3_61[16]}
   );
   gpc1_1 gpc2621 (
      {stage2_61[25]},
      {stage3_61[17]}
   );
   gpc1_1 gpc2622 (
      {stage2_61[26]},
      {stage3_61[18]}
   );
   gpc1_1 gpc2623 (
      {stage2_61[27]},
      {stage3_61[19]}
   );
   gpc1_1 gpc2624 (
      {stage2_61[28]},
      {stage3_61[20]}
   );
   gpc1_1 gpc2625 (
      {stage2_62[30]},
      {stage3_62[8]}
   );
   gpc1_1 gpc2626 (
      {stage2_62[31]},
      {stage3_62[9]}
   );
   gpc1_1 gpc2627 (
      {stage2_62[32]},
      {stage3_62[10]}
   );
   gpc1_1 gpc2628 (
      {stage2_62[33]},
      {stage3_62[11]}
   );
   gpc1_1 gpc2629 (
      {stage2_62[34]},
      {stage3_62[12]}
   );
   gpc1_1 gpc2630 (
      {stage2_62[35]},
      {stage3_62[13]}
   );
   gpc1_1 gpc2631 (
      {stage2_62[36]},
      {stage3_62[14]}
   );
   gpc1_1 gpc2632 (
      {stage2_62[37]},
      {stage3_62[15]}
   );
   gpc1_1 gpc2633 (
      {stage2_63[33]},
      {stage3_63[13]}
   );
   gpc1_1 gpc2634 (
      {stage2_63[34]},
      {stage3_63[14]}
   );
   gpc1_1 gpc2635 (
      {stage2_63[35]},
      {stage3_63[15]}
   );
   gpc1_1 gpc2636 (
      {stage2_63[36]},
      {stage3_63[16]}
   );
   gpc1_1 gpc2637 (
      {stage2_63[37]},
      {stage3_63[17]}
   );
   gpc1_1 gpc2638 (
      {stage2_65[15]},
      {stage3_65[9]}
   );
   gpc1_1 gpc2639 (
      {stage2_65[16]},
      {stage3_65[10]}
   );
   gpc1_1 gpc2640 (
      {stage2_65[17]},
      {stage3_65[11]}
   );
   gpc1_1 gpc2641 (
      {stage2_66[5]},
      {stage3_66[6]}
   );
   gpc1_1 gpc2642 (
      {stage2_67[0]},
      {stage3_67[5]}
   );
   gpc1_1 gpc2643 (
      {stage2_67[1]},
      {stage3_67[6]}
   );
   gpc615_5 gpc2644 (
      {stage3_0[0], stage3_0[1], stage3_0[2], stage3_0[3], stage3_0[4]},
      {stage3_1[0]},
      {stage3_2[0], stage3_2[1], stage3_2[2], stage3_2[3], stage3_2[4], stage3_2[5]},
      {stage4_4[0],stage4_3[0],stage4_2[0],stage4_1[0],stage4_0[0]}
   );
   gpc207_4 gpc2645 (
      {stage3_1[1], stage3_1[2], stage3_1[3], stage3_1[4], stage3_1[5], stage3_1[6], stage3_1[7]},
      {stage3_3[0], stage3_3[1]},
      {stage4_4[1],stage4_3[1],stage4_2[1],stage4_1[1]}
   );
   gpc615_5 gpc2646 (
      {stage3_3[2], stage3_3[3], stage3_3[4], stage3_3[5], stage3_3[6]},
      {stage3_4[0]},
      {stage3_5[0], stage3_5[1], stage3_5[2], stage3_5[3], stage3_5[4], stage3_5[5]},
      {stage4_7[0],stage4_6[0],stage4_5[0],stage4_4[2],stage4_3[2]}
   );
   gpc615_5 gpc2647 (
      {stage3_3[7], stage3_3[8], stage3_3[9], stage3_3[10], stage3_3[11]},
      {stage3_4[1]},
      {stage3_5[6], stage3_5[7], stage3_5[8], stage3_5[9], stage3_5[10], stage3_5[11]},
      {stage4_7[1],stage4_6[1],stage4_5[1],stage4_4[3],stage4_3[3]}
   );
   gpc615_5 gpc2648 (
      {stage3_3[12], stage3_3[13], stage3_3[14], stage3_3[15], stage3_3[16]},
      {stage3_4[2]},
      {stage3_5[12], stage3_5[13], stage3_5[14], stage3_5[15], stage3_5[16], stage3_5[17]},
      {stage4_7[2],stage4_6[2],stage4_5[2],stage4_4[4],stage4_3[4]}
   );
   gpc615_5 gpc2649 (
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4]},
      {stage3_7[0]},
      {stage3_8[0], stage3_8[1], stage3_8[2], stage3_8[3], stage3_8[4], stage3_8[5]},
      {stage4_10[0],stage4_9[0],stage4_8[0],stage4_7[3],stage4_6[3]}
   );
   gpc615_5 gpc2650 (
      {stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4], stage3_7[5]},
      {stage3_8[6]},
      {stage3_9[0], stage3_9[1], stage3_9[2], stage3_9[3], stage3_9[4], stage3_9[5]},
      {stage4_11[0],stage4_10[1],stage4_9[1],stage4_8[1],stage4_7[4]}
   );
   gpc615_5 gpc2651 (
      {stage3_7[6], stage3_7[7], stage3_7[8], stage3_7[9], stage3_7[10]},
      {stage3_8[7]},
      {stage3_9[6], stage3_9[7], stage3_9[8], stage3_9[9], stage3_9[10], stage3_9[11]},
      {stage4_11[1],stage4_10[2],stage4_9[2],stage4_8[2],stage4_7[5]}
   );
   gpc606_5 gpc2652 (
      {stage3_8[8], stage3_8[9], stage3_8[10], stage3_8[11], stage3_8[12], stage3_8[13]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage4_12[0],stage4_11[2],stage4_10[3],stage4_9[3],stage4_8[3]}
   );
   gpc606_5 gpc2653 (
      {stage3_9[12], stage3_9[13], stage3_9[14], stage3_9[15], stage3_9[16], stage3_9[17]},
      {stage3_11[0], stage3_11[1], stage3_11[2], stage3_11[3], stage3_11[4], stage3_11[5]},
      {stage4_13[0],stage4_12[1],stage4_11[3],stage4_10[4],stage4_9[4]}
   );
   gpc606_5 gpc2654 (
      {stage3_11[6], stage3_11[7], stage3_11[8], stage3_11[9], stage3_11[10], stage3_11[11]},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], stage3_13[5]},
      {stage4_15[0],stage4_14[0],stage4_13[1],stage4_12[2],stage4_11[4]}
   );
   gpc207_4 gpc2655 (
      {stage3_12[0], stage3_12[1], stage3_12[2], stage3_12[3], stage3_12[4], stage3_12[5], stage3_12[6]},
      {stage3_14[0], stage3_14[1]},
      {stage4_15[1],stage4_14[1],stage4_13[2],stage4_12[3]}
   );
   gpc606_5 gpc2656 (
      {stage3_12[7], stage3_12[8], stage3_12[9], stage3_12[10], stage3_12[11], stage3_12[12]},
      {stage3_14[2], stage3_14[3], stage3_14[4], stage3_14[5], stage3_14[6], stage3_14[7]},
      {stage4_16[0],stage4_15[2],stage4_14[2],stage4_13[3],stage4_12[4]}
   );
   gpc606_5 gpc2657 (
      {stage3_13[6], stage3_13[7], stage3_13[8], stage3_13[9], stage3_13[10], stage3_13[11]},
      {stage3_15[0], stage3_15[1], stage3_15[2], stage3_15[3], stage3_15[4], stage3_15[5]},
      {stage4_17[0],stage4_16[1],stage4_15[3],stage4_14[3],stage4_13[4]}
   );
   gpc207_4 gpc2658 (
      {stage3_15[6], stage3_15[7], stage3_15[8], stage3_15[9], stage3_15[10], stage3_15[11], stage3_15[12]},
      {stage3_17[0], stage3_17[1]},
      {stage4_18[0],stage4_17[1],stage4_16[2],stage4_15[4]}
   );
   gpc207_4 gpc2659 (
      {stage3_15[13], stage3_15[14], stage3_15[15], stage3_15[16], stage3_15[17], stage3_15[18], stage3_15[19]},
      {stage3_17[2], stage3_17[3]},
      {stage4_18[1],stage4_17[2],stage4_16[3],stage4_15[5]}
   );
   gpc615_5 gpc2660 (
      {stage3_15[20], stage3_15[21], stage3_15[22], stage3_15[23], stage3_15[24]},
      {stage3_16[0]},
      {stage3_17[4], stage3_17[5], stage3_17[6], stage3_17[7], stage3_17[8], stage3_17[9]},
      {stage4_19[0],stage4_18[2],stage4_17[3],stage4_16[4],stage4_15[6]}
   );
   gpc606_5 gpc2661 (
      {stage3_16[1], stage3_16[2], stage3_16[3], stage3_16[4], stage3_16[5], stage3_16[6]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage4_20[0],stage4_19[1],stage4_18[3],stage4_17[4],stage4_16[5]}
   );
   gpc606_5 gpc2662 (
      {stage3_16[7], stage3_16[8], stage3_16[9], stage3_16[10], stage3_16[11], 1'b0},
      {stage3_18[6], stage3_18[7], stage3_18[8], stage3_18[9], stage3_18[10], stage3_18[11]},
      {stage4_20[1],stage4_19[2],stage4_18[4],stage4_17[5],stage4_16[6]}
   );
   gpc615_5 gpc2663 (
      {stage3_19[0], stage3_19[1], stage3_19[2], stage3_19[3], stage3_19[4]},
      {stage3_20[0]},
      {stage3_21[0], stage3_21[1], stage3_21[2], stage3_21[3], stage3_21[4], stage3_21[5]},
      {stage4_23[0],stage4_22[0],stage4_21[0],stage4_20[2],stage4_19[3]}
   );
   gpc615_5 gpc2664 (
      {stage3_19[5], stage3_19[6], stage3_19[7], stage3_19[8], stage3_19[9]},
      {stage3_20[1]},
      {stage3_21[6], stage3_21[7], stage3_21[8], stage3_21[9], stage3_21[10], stage3_21[11]},
      {stage4_23[1],stage4_22[1],stage4_21[1],stage4_20[3],stage4_19[4]}
   );
   gpc615_5 gpc2665 (
      {stage3_19[10], stage3_19[11], stage3_19[12], stage3_19[13], stage3_19[14]},
      {stage3_20[2]},
      {stage3_21[12], stage3_21[13], stage3_21[14], stage3_21[15], stage3_21[16], stage3_21[17]},
      {stage4_23[2],stage4_22[2],stage4_21[2],stage4_20[4],stage4_19[5]}
   );
   gpc606_5 gpc2666 (
      {stage3_20[3], stage3_20[4], stage3_20[5], stage3_20[6], stage3_20[7], stage3_20[8]},
      {stage3_22[0], stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], stage3_22[5]},
      {stage4_24[0],stage4_23[3],stage4_22[3],stage4_21[3],stage4_20[5]}
   );
   gpc1163_5 gpc2667 (
      {stage3_22[6], stage3_22[7], stage3_22[8]},
      {stage3_23[0], stage3_23[1], stage3_23[2], stage3_23[3], stage3_23[4], stage3_23[5]},
      {stage3_24[0]},
      {stage3_25[0]},
      {stage4_26[0],stage4_25[0],stage4_24[1],stage4_23[4],stage4_22[4]}
   );
   gpc117_4 gpc2668 (
      {stage3_23[6], stage3_23[7], stage3_23[8], stage3_23[9], stage3_23[10], stage3_23[11], stage3_23[12]},
      {stage3_24[1]},
      {stage3_25[1]},
      {stage4_26[1],stage4_25[1],stage4_24[2],stage4_23[5]}
   );
   gpc207_4 gpc2669 (
      {stage3_24[2], stage3_24[3], stage3_24[4], stage3_24[5], stage3_24[6], stage3_24[7], stage3_24[8]},
      {stage3_26[0], stage3_26[1]},
      {stage4_27[0],stage4_26[2],stage4_25[2],stage4_24[3]}
   );
   gpc135_4 gpc2670 (
      {stage3_25[2], stage3_25[3], stage3_25[4], stage3_25[5], stage3_25[6]},
      {stage3_26[2], stage3_26[3], stage3_26[4]},
      {stage3_27[0]},
      {stage4_28[0],stage4_27[1],stage4_26[3],stage4_25[3]}
   );
   gpc135_4 gpc2671 (
      {stage3_25[7], stage3_25[8], stage3_25[9], stage3_25[10], stage3_25[11]},
      {stage3_26[5], stage3_26[6], stage3_26[7]},
      {stage3_27[1]},
      {stage4_28[1],stage4_27[2],stage4_26[4],stage4_25[4]}
   );
   gpc606_5 gpc2672 (
      {stage3_25[12], stage3_25[13], stage3_25[14], stage3_25[15], stage3_25[16], stage3_25[17]},
      {stage3_27[2], stage3_27[3], stage3_27[4], stage3_27[5], stage3_27[6], stage3_27[7]},
      {stage4_29[0],stage4_28[2],stage4_27[3],stage4_26[5],stage4_25[5]}
   );
   gpc1163_5 gpc2673 (
      {stage3_27[8], stage3_27[9], stage3_27[10]},
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4], stage3_28[5]},
      {stage3_29[0]},
      {stage3_30[0]},
      {stage4_31[0],stage4_30[0],stage4_29[1],stage4_28[3],stage4_27[4]}
   );
   gpc1163_5 gpc2674 (
      {stage3_27[11], stage3_27[12], stage3_27[13]},
      {stage3_28[6], stage3_28[7], stage3_28[8], stage3_28[9], stage3_28[10], stage3_28[11]},
      {stage3_29[1]},
      {stage3_30[1]},
      {stage4_31[1],stage4_30[1],stage4_29[2],stage4_28[4],stage4_27[5]}
   );
   gpc606_5 gpc2675 (
      {stage3_28[12], stage3_28[13], stage3_28[14], stage3_28[15], stage3_28[16], 1'b0},
      {stage3_30[2], stage3_30[3], stage3_30[4], stage3_30[5], stage3_30[6], stage3_30[7]},
      {stage4_32[0],stage4_31[2],stage4_30[2],stage4_29[3],stage4_28[5]}
   );
   gpc207_4 gpc2676 (
      {stage3_30[8], stage3_30[9], stage3_30[10], stage3_30[11], stage3_30[12], stage3_30[13], stage3_30[14]},
      {stage3_32[0], stage3_32[1]},
      {stage4_33[0],stage4_32[1],stage4_31[3],stage4_30[3]}
   );
   gpc207_4 gpc2677 (
      {stage3_31[0], stage3_31[1], stage3_31[2], stage3_31[3], stage3_31[4], stage3_31[5], stage3_31[6]},
      {stage3_33[0], stage3_33[1]},
      {stage4_34[0],stage4_33[1],stage4_32[2],stage4_31[4]}
   );
   gpc207_4 gpc2678 (
      {stage3_31[7], stage3_31[8], stage3_31[9], stage3_31[10], stage3_31[11], stage3_31[12], stage3_31[13]},
      {stage3_33[2], stage3_33[3]},
      {stage4_34[1],stage4_33[2],stage4_32[3],stage4_31[5]}
   );
   gpc606_5 gpc2679 (
      {stage3_31[14], stage3_31[15], stage3_31[16], stage3_31[17], stage3_31[18], stage3_31[19]},
      {stage3_33[4], stage3_33[5], stage3_33[6], stage3_33[7], stage3_33[8], stage3_33[9]},
      {stage4_35[0],stage4_34[2],stage4_33[3],stage4_32[4],stage4_31[6]}
   );
   gpc615_5 gpc2680 (
      {stage3_32[2], stage3_32[3], stage3_32[4], stage3_32[5], stage3_32[6]},
      {stage3_33[10]},
      {stage3_34[0], stage3_34[1], stage3_34[2], stage3_34[3], stage3_34[4], stage3_34[5]},
      {stage4_36[0],stage4_35[1],stage4_34[3],stage4_33[4],stage4_32[5]}
   );
   gpc615_5 gpc2681 (
      {stage3_32[7], stage3_32[8], stage3_32[9], stage3_32[10], stage3_32[11]},
      {stage3_33[11]},
      {stage3_34[6], stage3_34[7], stage3_34[8], stage3_34[9], stage3_34[10], stage3_34[11]},
      {stage4_36[1],stage4_35[2],stage4_34[4],stage4_33[5],stage4_32[6]}
   );
   gpc606_5 gpc2682 (
      {stage3_34[12], stage3_34[13], stage3_34[14], stage3_34[15], stage3_34[16], stage3_34[17]},
      {stage3_36[0], stage3_36[1], stage3_36[2], stage3_36[3], stage3_36[4], stage3_36[5]},
      {stage4_38[0],stage4_37[0],stage4_36[2],stage4_35[3],stage4_34[5]}
   );
   gpc117_4 gpc2683 (
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3], stage3_35[4], stage3_35[5], stage3_35[6]},
      {stage3_36[6]},
      {stage3_37[0]},
      {stage4_38[1],stage4_37[1],stage4_36[3],stage4_35[4]}
   );
   gpc1163_5 gpc2684 (
      {stage3_35[7], stage3_35[8], stage3_35[9]},
      {stage3_36[7], stage3_36[8], stage3_36[9], stage3_36[10], stage3_36[11], stage3_36[12]},
      {stage3_37[1]},
      {stage3_38[0]},
      {stage4_39[0],stage4_38[2],stage4_37[2],stage4_36[4],stage4_35[5]}
   );
   gpc1163_5 gpc2685 (
      {stage3_37[2], stage3_37[3], stage3_37[4]},
      {stage3_38[1], stage3_38[2], stage3_38[3], stage3_38[4], stage3_38[5], stage3_38[6]},
      {stage3_39[0]},
      {stage3_40[0]},
      {stage4_41[0],stage4_40[0],stage4_39[1],stage4_38[3],stage4_37[3]}
   );
   gpc1163_5 gpc2686 (
      {stage3_37[5], stage3_37[6], stage3_37[7]},
      {stage3_38[7], stage3_38[8], stage3_38[9], stage3_38[10], stage3_38[11], stage3_38[12]},
      {stage3_39[1]},
      {stage3_40[1]},
      {stage4_41[1],stage4_40[1],stage4_39[2],stage4_38[4],stage4_37[4]}
   );
   gpc606_5 gpc2687 (
      {stage3_37[8], stage3_37[9], stage3_37[10], stage3_37[11], stage3_37[12], stage3_37[13]},
      {stage3_39[2], stage3_39[3], stage3_39[4], stage3_39[5], stage3_39[6], stage3_39[7]},
      {stage4_41[2],stage4_40[2],stage4_39[3],stage4_38[5],stage4_37[5]}
   );
   gpc223_4 gpc2688 (
      {stage3_39[8], stage3_39[9], stage3_39[10]},
      {stage3_40[2], stage3_40[3]},
      {stage3_41[0], stage3_41[1]},
      {stage4_42[0],stage4_41[3],stage4_40[3],stage4_39[4]}
   );
   gpc623_5 gpc2689 (
      {stage3_40[4], stage3_40[5], stage3_40[6]},
      {stage3_41[2], stage3_41[3]},
      {stage3_42[0], stage3_42[1], stage3_42[2], stage3_42[3], stage3_42[4], stage3_42[5]},
      {stage4_44[0],stage4_43[0],stage4_42[1],stage4_41[4],stage4_40[4]}
   );
   gpc623_5 gpc2690 (
      {stage3_40[7], stage3_40[8], stage3_40[9]},
      {stage3_41[4], stage3_41[5]},
      {stage3_42[6], stage3_42[7], stage3_42[8], stage3_42[9], stage3_42[10], stage3_42[11]},
      {stage4_44[1],stage4_43[1],stage4_42[2],stage4_41[5],stage4_40[5]}
   );
   gpc623_5 gpc2691 (
      {stage3_40[10], stage3_40[11], stage3_40[12]},
      {stage3_41[6], stage3_41[7]},
      {stage3_42[12], stage3_42[13], stage3_42[14], stage3_42[15], stage3_42[16], stage3_42[17]},
      {stage4_44[2],stage4_43[2],stage4_42[3],stage4_41[6],stage4_40[6]}
   );
   gpc615_5 gpc2692 (
      {stage3_43[0], stage3_43[1], stage3_43[2], stage3_43[3], stage3_43[4]},
      {stage3_44[0]},
      {stage3_45[0], stage3_45[1], stage3_45[2], stage3_45[3], stage3_45[4], stage3_45[5]},
      {stage4_47[0],stage4_46[0],stage4_45[0],stage4_44[3],stage4_43[3]}
   );
   gpc615_5 gpc2693 (
      {stage3_43[5], stage3_43[6], stage3_43[7], stage3_43[8], stage3_43[9]},
      {stage3_44[1]},
      {stage3_45[6], stage3_45[7], stage3_45[8], stage3_45[9], stage3_45[10], stage3_45[11]},
      {stage4_47[1],stage4_46[1],stage4_45[1],stage4_44[4],stage4_43[4]}
   );
   gpc207_4 gpc2694 (
      {stage3_44[2], stage3_44[3], stage3_44[4], stage3_44[5], stage3_44[6], stage3_44[7], 1'b0},
      {stage3_46[0], stage3_46[1]},
      {stage4_47[2],stage4_46[2],stage4_45[2],stage4_44[5]}
   );
   gpc606_5 gpc2695 (
      {stage3_46[2], stage3_46[3], stage3_46[4], stage3_46[5], stage3_46[6], stage3_46[7]},
      {stage3_48[0], stage3_48[1], stage3_48[2], stage3_48[3], stage3_48[4], stage3_48[5]},
      {stage4_50[0],stage4_49[0],stage4_48[0],stage4_47[3],stage4_46[3]}
   );
   gpc623_5 gpc2696 (
      {stage3_46[8], stage3_46[9], stage3_46[10]},
      {stage3_47[0], stage3_47[1]},
      {stage3_48[6], stage3_48[7], stage3_48[8], stage3_48[9], stage3_48[10], stage3_48[11]},
      {stage4_50[1],stage4_49[1],stage4_48[1],stage4_47[4],stage4_46[4]}
   );
   gpc135_4 gpc2697 (
      {stage3_47[2], stage3_47[3], stage3_47[4], stage3_47[5], stage3_47[6]},
      {stage3_48[12], stage3_48[13], stage3_48[14]},
      {stage3_49[0]},
      {stage4_50[2],stage4_49[2],stage4_48[2],stage4_47[5]}
   );
   gpc135_4 gpc2698 (
      {stage3_47[7], stage3_47[8], stage3_47[9], stage3_47[10], 1'b0},
      {stage3_48[15], stage3_48[16], stage3_48[17]},
      {stage3_49[1]},
      {stage4_50[3],stage4_49[3],stage4_48[3],stage4_47[6]}
   );
   gpc615_5 gpc2699 (
      {stage3_49[2], stage3_49[3], stage3_49[4], stage3_49[5], stage3_49[6]},
      {stage3_50[0]},
      {stage3_51[0], stage3_51[1], stage3_51[2], stage3_51[3], stage3_51[4], stage3_51[5]},
      {stage4_53[0],stage4_52[0],stage4_51[0],stage4_50[4],stage4_49[4]}
   );
   gpc615_5 gpc2700 (
      {stage3_49[7], stage3_49[8], stage3_49[9], stage3_49[10], stage3_49[11]},
      {stage3_50[1]},
      {stage3_51[6], stage3_51[7], stage3_51[8], stage3_51[9], stage3_51[10], stage3_51[11]},
      {stage4_53[1],stage4_52[1],stage4_51[1],stage4_50[5],stage4_49[5]}
   );
   gpc615_5 gpc2701 (
      {stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5], stage3_50[6]},
      {stage3_51[12]},
      {stage3_52[0], stage3_52[1], stage3_52[2], stage3_52[3], stage3_52[4], stage3_52[5]},
      {stage4_54[0],stage4_53[2],stage4_52[2],stage4_51[2],stage4_50[6]}
   );
   gpc1343_5 gpc2702 (
      {stage3_53[0], stage3_53[1], stage3_53[2]},
      {stage3_54[0], stage3_54[1], stage3_54[2], stage3_54[3]},
      {stage3_55[0], stage3_55[1], stage3_55[2]},
      {stage3_56[0]},
      {stage4_57[0],stage4_56[0],stage4_55[0],stage4_54[1],stage4_53[3]}
   );
   gpc1343_5 gpc2703 (
      {stage3_53[3], stage3_53[4], stage3_53[5]},
      {stage3_54[4], stage3_54[5], stage3_54[6], stage3_54[7]},
      {stage3_55[3], stage3_55[4], stage3_55[5]},
      {stage3_56[1]},
      {stage4_57[1],stage4_56[1],stage4_55[1],stage4_54[2],stage4_53[4]}
   );
   gpc1343_5 gpc2704 (
      {stage3_53[6], stage3_53[7], stage3_53[8]},
      {stage3_54[8], stage3_54[9], stage3_54[10], stage3_54[11]},
      {stage3_55[6], stage3_55[7], stage3_55[8]},
      {stage3_56[2]},
      {stage4_57[2],stage4_56[2],stage4_55[2],stage4_54[3],stage4_53[5]}
   );
   gpc135_4 gpc2705 (
      {stage3_54[12], stage3_54[13], stage3_54[14], stage3_54[15], stage3_54[16]},
      {stage3_55[9], stage3_55[10], stage3_55[11]},
      {stage3_56[3]},
      {stage4_57[3],stage4_56[3],stage4_55[3],stage4_54[4]}
   );
   gpc606_5 gpc2706 (
      {stage3_57[0], stage3_57[1], stage3_57[2], stage3_57[3], stage3_57[4], stage3_57[5]},
      {stage3_59[0], stage3_59[1], stage3_59[2], stage3_59[3], stage3_59[4], stage3_59[5]},
      {stage4_61[0],stage4_60[0],stage4_59[0],stage4_58[0],stage4_57[4]}
   );
   gpc606_5 gpc2707 (
      {stage3_57[6], stage3_57[7], stage3_57[8], stage3_57[9], stage3_57[10], stage3_57[11]},
      {stage3_59[6], stage3_59[7], stage3_59[8], stage3_59[9], stage3_59[10], stage3_59[11]},
      {stage4_61[1],stage4_60[1],stage4_59[1],stage4_58[1],stage4_57[5]}
   );
   gpc207_4 gpc2708 (
      {stage3_58[0], stage3_58[1], stage3_58[2], stage3_58[3], stage3_58[4], stage3_58[5], stage3_58[6]},
      {stage3_60[0], stage3_60[1]},
      {stage4_61[2],stage4_60[2],stage4_59[2],stage4_58[2]}
   );
   gpc207_4 gpc2709 (
      {stage3_58[7], stage3_58[8], stage3_58[9], stage3_58[10], stage3_58[11], 1'b0, 1'b0},
      {stage3_60[2], stage3_60[3]},
      {stage4_61[3],stage4_60[3],stage4_59[3],stage4_58[3]}
   );
   gpc606_5 gpc2710 (
      {stage3_60[4], stage3_60[5], stage3_60[6], stage3_60[7], stage3_60[8], stage3_60[9]},
      {stage3_62[0], stage3_62[1], stage3_62[2], stage3_62[3], stage3_62[4], stage3_62[5]},
      {stage4_64[0],stage4_63[0],stage4_62[0],stage4_61[4],stage4_60[4]}
   );
   gpc606_5 gpc2711 (
      {stage3_60[10], stage3_60[11], stage3_60[12], stage3_60[13], 1'b0, 1'b0},
      {stage3_62[6], stage3_62[7], stage3_62[8], stage3_62[9], stage3_62[10], stage3_62[11]},
      {stage4_64[1],stage4_63[1],stage4_62[1],stage4_61[5],stage4_60[5]}
   );
   gpc117_4 gpc2712 (
      {stage3_61[0], stage3_61[1], stage3_61[2], stage3_61[3], stage3_61[4], stage3_61[5], stage3_61[6]},
      {stage3_62[12]},
      {stage3_63[0]},
      {stage4_64[2],stage4_63[2],stage4_62[2],stage4_61[6]}
   );
   gpc207_4 gpc2713 (
      {stage3_61[7], stage3_61[8], stage3_61[9], stage3_61[10], stage3_61[11], stage3_61[12], stage3_61[13]},
      {stage3_63[1], stage3_63[2]},
      {stage4_64[3],stage4_63[3],stage4_62[3],stage4_61[7]}
   );
   gpc606_5 gpc2714 (
      {stage3_61[14], stage3_61[15], stage3_61[16], stage3_61[17], stage3_61[18], stage3_61[19]},
      {stage3_63[3], stage3_63[4], stage3_63[5], stage3_63[6], stage3_63[7], stage3_63[8]},
      {stage4_65[0],stage4_64[4],stage4_63[4],stage4_62[4],stage4_61[8]}
   );
   gpc615_5 gpc2715 (
      {stage3_62[13], stage3_62[14], stage3_62[15], 1'b0, 1'b0},
      {stage3_63[9]},
      {stage3_64[0], stage3_64[1], stage3_64[2], stage3_64[3], stage3_64[4], stage3_64[5]},
      {stage4_66[0],stage4_65[1],stage4_64[5],stage4_63[5],stage4_62[5]}
   );
   gpc606_5 gpc2716 (
      {stage3_63[10], stage3_63[11], stage3_63[12], stage3_63[13], stage3_63[14], stage3_63[15]},
      {stage3_65[0], stage3_65[1], stage3_65[2], stage3_65[3], stage3_65[4], stage3_65[5]},
      {stage4_67[0],stage4_66[1],stage4_65[2],stage4_64[6],stage4_63[6]}
   );
   gpc606_5 gpc2717 (
      {stage3_64[6], stage3_64[7], stage3_64[8], stage3_64[9], stage3_64[10], stage3_64[11]},
      {stage3_66[0], stage3_66[1], stage3_66[2], stage3_66[3], stage3_66[4], stage3_66[5]},
      {stage4_68[0],stage4_67[1],stage4_66[2],stage4_65[3],stage4_64[7]}
   );
   gpc606_5 gpc2718 (
      {stage3_65[6], stage3_65[7], stage3_65[8], stage3_65[9], stage3_65[10], stage3_65[11]},
      {stage3_67[0], stage3_67[1], stage3_67[2], stage3_67[3], stage3_67[4], stage3_67[5]},
      {stage4_69[0],stage4_68[1],stage4_67[2],stage4_66[3],stage4_65[4]}
   );
   gpc1_1 gpc2719 (
      {stage3_3[17]},
      {stage4_3[5]}
   );
   gpc1_1 gpc2720 (
      {stage3_3[18]},
      {stage4_3[6]}
   );
   gpc1_1 gpc2721 (
      {stage3_3[19]},
      {stage4_3[7]}
   );
   gpc1_1 gpc2722 (
      {stage3_3[20]},
      {stage4_3[8]}
   );
   gpc1_1 gpc2723 (
      {stage3_3[21]},
      {stage4_3[9]}
   );
   gpc1_1 gpc2724 (
      {stage3_4[3]},
      {stage4_4[5]}
   );
   gpc1_1 gpc2725 (
      {stage3_4[4]},
      {stage4_4[6]}
   );
   gpc1_1 gpc2726 (
      {stage3_4[5]},
      {stage4_4[7]}
   );
   gpc1_1 gpc2727 (
      {stage3_4[6]},
      {stage4_4[8]}
   );
   gpc1_1 gpc2728 (
      {stage3_4[7]},
      {stage4_4[9]}
   );
   gpc1_1 gpc2729 (
      {stage3_4[8]},
      {stage4_4[10]}
   );
   gpc1_1 gpc2730 (
      {stage3_4[9]},
      {stage4_4[11]}
   );
   gpc1_1 gpc2731 (
      {stage3_4[10]},
      {stage4_4[12]}
   );
   gpc1_1 gpc2732 (
      {stage3_4[11]},
      {stage4_4[13]}
   );
   gpc1_1 gpc2733 (
      {stage3_5[18]},
      {stage4_5[3]}
   );
   gpc1_1 gpc2734 (
      {stage3_5[19]},
      {stage4_5[4]}
   );
   gpc1_1 gpc2735 (
      {stage3_5[20]},
      {stage4_5[5]}
   );
   gpc1_1 gpc2736 (
      {stage3_5[21]},
      {stage4_5[6]}
   );
   gpc1_1 gpc2737 (
      {stage3_5[22]},
      {stage4_5[7]}
   );
   gpc1_1 gpc2738 (
      {stage3_5[23]},
      {stage4_5[8]}
   );
   gpc1_1 gpc2739 (
      {stage3_6[5]},
      {stage4_6[4]}
   );
   gpc1_1 gpc2740 (
      {stage3_6[6]},
      {stage4_6[5]}
   );
   gpc1_1 gpc2741 (
      {stage3_6[7]},
      {stage4_6[6]}
   );
   gpc1_1 gpc2742 (
      {stage3_6[8]},
      {stage4_6[7]}
   );
   gpc1_1 gpc2743 (
      {stage3_6[9]},
      {stage4_6[8]}
   );
   gpc1_1 gpc2744 (
      {stage3_7[11]},
      {stage4_7[6]}
   );
   gpc1_1 gpc2745 (
      {stage3_8[14]},
      {stage4_8[4]}
   );
   gpc1_1 gpc2746 (
      {stage3_8[15]},
      {stage4_8[5]}
   );
   gpc1_1 gpc2747 (
      {stage3_9[18]},
      {stage4_9[5]}
   );
   gpc1_1 gpc2748 (
      {stage3_9[19]},
      {stage4_9[6]}
   );
   gpc1_1 gpc2749 (
      {stage3_10[6]},
      {stage4_10[5]}
   );
   gpc1_1 gpc2750 (
      {stage3_10[7]},
      {stage4_10[6]}
   );
   gpc1_1 gpc2751 (
      {stage3_10[8]},
      {stage4_10[7]}
   );
   gpc1_1 gpc2752 (
      {stage3_10[9]},
      {stage4_10[8]}
   );
   gpc1_1 gpc2753 (
      {stage3_10[10]},
      {stage4_10[9]}
   );
   gpc1_1 gpc2754 (
      {stage3_10[11]},
      {stage4_10[10]}
   );
   gpc1_1 gpc2755 (
      {stage3_11[12]},
      {stage4_11[5]}
   );
   gpc1_1 gpc2756 (
      {stage3_12[13]},
      {stage4_12[5]}
   );
   gpc1_1 gpc2757 (
      {stage3_14[8]},
      {stage4_14[4]}
   );
   gpc1_1 gpc2758 (
      {stage3_14[9]},
      {stage4_14[5]}
   );
   gpc1_1 gpc2759 (
      {stage3_15[25]},
      {stage4_15[7]}
   );
   gpc1_1 gpc2760 (
      {stage3_17[10]},
      {stage4_17[6]}
   );
   gpc1_1 gpc2761 (
      {stage3_17[11]},
      {stage4_17[7]}
   );
   gpc1_1 gpc2762 (
      {stage3_18[12]},
      {stage4_18[5]}
   );
   gpc1_1 gpc2763 (
      {stage3_19[15]},
      {stage4_19[6]}
   );
   gpc1_1 gpc2764 (
      {stage3_20[9]},
      {stage4_20[6]}
   );
   gpc1_1 gpc2765 (
      {stage3_20[10]},
      {stage4_20[7]}
   );
   gpc1_1 gpc2766 (
      {stage3_20[11]},
      {stage4_20[8]}
   );
   gpc1_1 gpc2767 (
      {stage3_20[12]},
      {stage4_20[9]}
   );
   gpc1_1 gpc2768 (
      {stage3_20[13]},
      {stage4_20[10]}
   );
   gpc1_1 gpc2769 (
      {stage3_24[9]},
      {stage4_24[4]}
   );
   gpc1_1 gpc2770 (
      {stage3_24[10]},
      {stage4_24[5]}
   );
   gpc1_1 gpc2771 (
      {stage3_24[11]},
      {stage4_24[6]}
   );
   gpc1_1 gpc2772 (
      {stage3_24[12]},
      {stage4_24[7]}
   );
   gpc1_1 gpc2773 (
      {stage3_24[13]},
      {stage4_24[8]}
   );
   gpc1_1 gpc2774 (
      {stage3_24[14]},
      {stage4_24[9]}
   );
   gpc1_1 gpc2775 (
      {stage3_24[15]},
      {stage4_24[10]}
   );
   gpc1_1 gpc2776 (
      {stage3_25[18]},
      {stage4_25[6]}
   );
   gpc1_1 gpc2777 (
      {stage3_25[19]},
      {stage4_25[7]}
   );
   gpc1_1 gpc2778 (
      {stage3_26[8]},
      {stage4_26[6]}
   );
   gpc1_1 gpc2779 (
      {stage3_26[9]},
      {stage4_26[7]}
   );
   gpc1_1 gpc2780 (
      {stage3_26[10]},
      {stage4_26[8]}
   );
   gpc1_1 gpc2781 (
      {stage3_26[11]},
      {stage4_26[9]}
   );
   gpc1_1 gpc2782 (
      {stage3_26[12]},
      {stage4_26[10]}
   );
   gpc1_1 gpc2783 (
      {stage3_29[2]},
      {stage4_29[4]}
   );
   gpc1_1 gpc2784 (
      {stage3_29[3]},
      {stage4_29[5]}
   );
   gpc1_1 gpc2785 (
      {stage3_29[4]},
      {stage4_29[6]}
   );
   gpc1_1 gpc2786 (
      {stage3_29[5]},
      {stage4_29[7]}
   );
   gpc1_1 gpc2787 (
      {stage3_29[6]},
      {stage4_29[8]}
   );
   gpc1_1 gpc2788 (
      {stage3_29[7]},
      {stage4_29[9]}
   );
   gpc1_1 gpc2789 (
      {stage3_36[13]},
      {stage4_36[5]}
   );
   gpc1_1 gpc2790 (
      {stage3_36[14]},
      {stage4_36[6]}
   );
   gpc1_1 gpc2791 (
      {stage3_37[14]},
      {stage4_37[6]}
   );
   gpc1_1 gpc2792 (
      {stage3_39[11]},
      {stage4_39[5]}
   );
   gpc1_1 gpc2793 (
      {stage3_39[12]},
      {stage4_39[6]}
   );
   gpc1_1 gpc2794 (
      {stage3_39[13]},
      {stage4_39[7]}
   );
   gpc1_1 gpc2795 (
      {stage3_40[13]},
      {stage4_40[7]}
   );
   gpc1_1 gpc2796 (
      {stage3_40[14]},
      {stage4_40[8]}
   );
   gpc1_1 gpc2797 (
      {stage3_40[15]},
      {stage4_40[9]}
   );
   gpc1_1 gpc2798 (
      {stage3_40[16]},
      {stage4_40[10]}
   );
   gpc1_1 gpc2799 (
      {stage3_40[17]},
      {stage4_40[11]}
   );
   gpc1_1 gpc2800 (
      {stage3_41[8]},
      {stage4_41[7]}
   );
   gpc1_1 gpc2801 (
      {stage3_41[9]},
      {stage4_41[8]}
   );
   gpc1_1 gpc2802 (
      {stage3_41[10]},
      {stage4_41[9]}
   );
   gpc1_1 gpc2803 (
      {stage3_41[11]},
      {stage4_41[10]}
   );
   gpc1_1 gpc2804 (
      {stage3_42[18]},
      {stage4_42[4]}
   );
   gpc1_1 gpc2805 (
      {stage3_42[19]},
      {stage4_42[5]}
   );
   gpc1_1 gpc2806 (
      {stage3_45[12]},
      {stage4_45[3]}
   );
   gpc1_1 gpc2807 (
      {stage3_45[13]},
      {stage4_45[4]}
   );
   gpc1_1 gpc2808 (
      {stage3_45[14]},
      {stage4_45[5]}
   );
   gpc1_1 gpc2809 (
      {stage3_46[11]},
      {stage4_46[5]}
   );
   gpc1_1 gpc2810 (
      {stage3_48[18]},
      {stage4_48[4]}
   );
   gpc1_1 gpc2811 (
      {stage3_52[6]},
      {stage4_52[3]}
   );
   gpc1_1 gpc2812 (
      {stage3_52[7]},
      {stage4_52[4]}
   );
   gpc1_1 gpc2813 (
      {stage3_52[8]},
      {stage4_52[5]}
   );
   gpc1_1 gpc2814 (
      {stage3_52[9]},
      {stage4_52[6]}
   );
   gpc1_1 gpc2815 (
      {stage3_52[10]},
      {stage4_52[7]}
   );
   gpc1_1 gpc2816 (
      {stage3_52[11]},
      {stage4_52[8]}
   );
   gpc1_1 gpc2817 (
      {stage3_52[12]},
      {stage4_52[9]}
   );
   gpc1_1 gpc2818 (
      {stage3_52[13]},
      {stage4_52[10]}
   );
   gpc1_1 gpc2819 (
      {stage3_52[14]},
      {stage4_52[11]}
   );
   gpc1_1 gpc2820 (
      {stage3_52[15]},
      {stage4_52[12]}
   );
   gpc1_1 gpc2821 (
      {stage3_52[16]},
      {stage4_52[13]}
   );
   gpc1_1 gpc2822 (
      {stage3_52[17]},
      {stage4_52[14]}
   );
   gpc1_1 gpc2823 (
      {stage3_52[18]},
      {stage4_52[15]}
   );
   gpc1_1 gpc2824 (
      {stage3_52[19]},
      {stage4_52[16]}
   );
   gpc1_1 gpc2825 (
      {stage3_54[17]},
      {stage4_54[5]}
   );
   gpc1_1 gpc2826 (
      {stage3_54[18]},
      {stage4_54[6]}
   );
   gpc1_1 gpc2827 (
      {stage3_54[19]},
      {stage4_54[7]}
   );
   gpc1_1 gpc2828 (
      {stage3_54[20]},
      {stage4_54[8]}
   );
   gpc1_1 gpc2829 (
      {stage3_54[21]},
      {stage4_54[9]}
   );
   gpc1_1 gpc2830 (
      {stage3_54[22]},
      {stage4_54[10]}
   );
   gpc1_1 gpc2831 (
      {stage3_54[23]},
      {stage4_54[11]}
   );
   gpc1_1 gpc2832 (
      {stage3_56[4]},
      {stage4_56[4]}
   );
   gpc1_1 gpc2833 (
      {stage3_56[5]},
      {stage4_56[5]}
   );
   gpc1_1 gpc2834 (
      {stage3_56[6]},
      {stage4_56[6]}
   );
   gpc1_1 gpc2835 (
      {stage3_56[7]},
      {stage4_56[7]}
   );
   gpc1_1 gpc2836 (
      {stage3_59[12]},
      {stage4_59[4]}
   );
   gpc1_1 gpc2837 (
      {stage3_59[13]},
      {stage4_59[5]}
   );
   gpc1_1 gpc2838 (
      {stage3_61[20]},
      {stage4_61[9]}
   );
   gpc1_1 gpc2839 (
      {stage3_63[16]},
      {stage4_63[7]}
   );
   gpc1_1 gpc2840 (
      {stage3_63[17]},
      {stage4_63[8]}
   );
   gpc1_1 gpc2841 (
      {stage3_64[12]},
      {stage4_64[8]}
   );
   gpc1_1 gpc2842 (
      {stage3_66[6]},
      {stage4_66[4]}
   );
   gpc1_1 gpc2843 (
      {stage3_67[6]},
      {stage4_67[3]}
   );
   gpc117_4 gpc2844 (
      {stage4_3[0], stage4_3[1], stage4_3[2], stage4_3[3], stage4_3[4], stage4_3[5], stage4_3[6]},
      {stage4_4[0]},
      {stage4_5[0]},
      {stage5_6[0],stage5_5[0],stage5_4[0],stage5_3[0]}
   );
   gpc606_5 gpc2845 (
      {stage4_4[1], stage4_4[2], stage4_4[3], stage4_4[4], stage4_4[5], stage4_4[6]},
      {stage4_6[0], stage4_6[1], stage4_6[2], stage4_6[3], stage4_6[4], stage4_6[5]},
      {stage5_8[0],stage5_7[0],stage5_6[1],stage5_5[1],stage5_4[1]}
   );
   gpc1325_5 gpc2846 (
      {stage4_4[7], stage4_4[8], stage4_4[9], stage4_4[10], stage4_4[11]},
      {stage4_5[1], stage4_5[2]},
      {stage4_6[6], stage4_6[7], stage4_6[8]},
      {stage4_7[0]},
      {stage5_8[1],stage5_7[1],stage5_6[2],stage5_5[2],stage5_4[2]}
   );
   gpc606_5 gpc2847 (
      {stage4_5[3], stage4_5[4], stage4_5[5], stage4_5[6], stage4_5[7], stage4_5[8]},
      {stage4_7[1], stage4_7[2], stage4_7[3], stage4_7[4], stage4_7[5], stage4_7[6]},
      {stage5_9[0],stage5_8[2],stage5_7[2],stage5_6[3],stage5_5[3]}
   );
   gpc606_5 gpc2848 (
      {stage4_8[0], stage4_8[1], stage4_8[2], stage4_8[3], stage4_8[4], stage4_8[5]},
      {stage4_10[0], stage4_10[1], stage4_10[2], stage4_10[3], stage4_10[4], stage4_10[5]},
      {stage5_12[0],stage5_11[0],stage5_10[0],stage5_9[1],stage5_8[3]}
   );
   gpc606_5 gpc2849 (
      {stage4_9[0], stage4_9[1], stage4_9[2], stage4_9[3], stage4_9[4], stage4_9[5]},
      {stage4_11[0], stage4_11[1], stage4_11[2], stage4_11[3], stage4_11[4], stage4_11[5]},
      {stage5_13[0],stage5_12[1],stage5_11[1],stage5_10[1],stage5_9[2]}
   );
   gpc623_5 gpc2850 (
      {stage4_12[0], stage4_12[1], stage4_12[2]},
      {stage4_13[0], stage4_13[1]},
      {stage4_14[0], stage4_14[1], stage4_14[2], stage4_14[3], stage4_14[4], stage4_14[5]},
      {stage5_16[0],stage5_15[0],stage5_14[0],stage5_13[1],stage5_12[2]}
   );
   gpc615_5 gpc2851 (
      {stage4_16[0], stage4_16[1], stage4_16[2], stage4_16[3], stage4_16[4]},
      {stage4_17[0]},
      {stage4_18[0], stage4_18[1], stage4_18[2], stage4_18[3], stage4_18[4], stage4_18[5]},
      {stage5_20[0],stage5_19[0],stage5_18[0],stage5_17[0],stage5_16[1]}
   );
   gpc606_5 gpc2852 (
      {stage4_17[1], stage4_17[2], stage4_17[3], stage4_17[4], stage4_17[5], stage4_17[6]},
      {stage4_19[0], stage4_19[1], stage4_19[2], stage4_19[3], stage4_19[4], stage4_19[5]},
      {stage5_21[0],stage5_20[1],stage5_19[1],stage5_18[1],stage5_17[1]}
   );
   gpc15_3 gpc2853 (
      {stage4_20[0], stage4_20[1], stage4_20[2], stage4_20[3], stage4_20[4]},
      {stage4_21[0]},
      {stage5_22[0],stage5_21[1],stage5_20[2]}
   );
   gpc1163_5 gpc2854 (
      {stage4_22[0], stage4_22[1], stage4_22[2]},
      {stage4_23[0], stage4_23[1], stage4_23[2], stage4_23[3], stage4_23[4], stage4_23[5]},
      {stage4_24[0]},
      {stage4_25[0]},
      {stage5_26[0],stage5_25[0],stage5_24[0],stage5_23[0],stage5_22[1]}
   );
   gpc606_5 gpc2855 (
      {stage4_24[1], stage4_24[2], stage4_24[3], stage4_24[4], stage4_24[5], stage4_24[6]},
      {stage4_26[0], stage4_26[1], stage4_26[2], stage4_26[3], stage4_26[4], stage4_26[5]},
      {stage5_28[0],stage5_27[0],stage5_26[1],stage5_25[1],stage5_24[1]}
   );
   gpc7_3 gpc2856 (
      {stage4_25[1], stage4_25[2], stage4_25[3], stage4_25[4], stage4_25[5], stage4_25[6], stage4_25[7]},
      {stage5_27[1],stage5_26[2],stage5_25[2]}
   );
   gpc615_5 gpc2857 (
      {stage4_26[6], stage4_26[7], stage4_26[8], stage4_26[9], stage4_26[10]},
      {stage4_27[0]},
      {stage4_28[0], stage4_28[1], stage4_28[2], stage4_28[3], stage4_28[4], stage4_28[5]},
      {stage5_30[0],stage5_29[0],stage5_28[1],stage5_27[2],stage5_26[3]}
   );
   gpc606_5 gpc2858 (
      {stage4_29[0], stage4_29[1], stage4_29[2], stage4_29[3], stage4_29[4], stage4_29[5]},
      {stage4_31[0], stage4_31[1], stage4_31[2], stage4_31[3], stage4_31[4], stage4_31[5]},
      {stage5_33[0],stage5_32[0],stage5_31[0],stage5_30[1],stage5_29[1]}
   );
   gpc623_5 gpc2859 (
      {stage4_30[0], stage4_30[1], stage4_30[2]},
      {stage4_31[6], 1'b0},
      {stage4_32[0], stage4_32[1], stage4_32[2], stage4_32[3], stage4_32[4], stage4_32[5]},
      {stage5_34[0],stage5_33[1],stage5_32[1],stage5_31[1],stage5_30[2]}
   );
   gpc606_5 gpc2860 (
      {stage4_33[0], stage4_33[1], stage4_33[2], stage4_33[3], stage4_33[4], stage4_33[5]},
      {stage4_35[0], stage4_35[1], stage4_35[2], stage4_35[3], stage4_35[4], stage4_35[5]},
      {stage5_37[0],stage5_36[0],stage5_35[0],stage5_34[1],stage5_33[2]}
   );
   gpc7_3 gpc2861 (
      {stage4_36[0], stage4_36[1], stage4_36[2], stage4_36[3], stage4_36[4], stage4_36[5], stage4_36[6]},
      {stage5_38[0],stage5_37[1],stage5_36[1]}
   );
   gpc7_3 gpc2862 (
      {stage4_37[0], stage4_37[1], stage4_37[2], stage4_37[3], stage4_37[4], stage4_37[5], stage4_37[6]},
      {stage5_39[0],stage5_38[1],stage5_37[2]}
   );
   gpc615_5 gpc2863 (
      {stage4_38[0], stage4_38[1], stage4_38[2], stage4_38[3], stage4_38[4]},
      {stage4_39[0]},
      {stage4_40[0], stage4_40[1], stage4_40[2], stage4_40[3], stage4_40[4], stage4_40[5]},
      {stage5_42[0],stage5_41[0],stage5_40[0],stage5_39[1],stage5_38[2]}
   );
   gpc615_5 gpc2864 (
      {stage4_39[1], stage4_39[2], stage4_39[3], stage4_39[4], stage4_39[5]},
      {stage4_40[6]},
      {stage4_41[0], stage4_41[1], stage4_41[2], stage4_41[3], stage4_41[4], stage4_41[5]},
      {stage5_43[0],stage5_42[1],stage5_41[1],stage5_40[1],stage5_39[2]}
   );
   gpc606_5 gpc2865 (
      {stage4_40[7], stage4_40[8], stage4_40[9], stage4_40[10], stage4_40[11], 1'b0},
      {stage4_42[0], stage4_42[1], stage4_42[2], stage4_42[3], stage4_42[4], stage4_42[5]},
      {stage5_44[0],stage5_43[1],stage5_42[2],stage5_41[2],stage5_40[2]}
   );
   gpc15_3 gpc2866 (
      {stage4_41[6], stage4_41[7], stage4_41[8], stage4_41[9], stage4_41[10]},
      {1'b0},
      {stage5_43[2],stage5_42[3],stage5_41[3]}
   );
   gpc606_5 gpc2867 (
      {stage4_43[0], stage4_43[1], stage4_43[2], stage4_43[3], stage4_43[4], 1'b0},
      {stage4_45[0], stage4_45[1], stage4_45[2], stage4_45[3], stage4_45[4], stage4_45[5]},
      {stage5_47[0],stage5_46[0],stage5_45[0],stage5_44[1],stage5_43[3]}
   );
   gpc615_5 gpc2868 (
      {stage4_44[0], stage4_44[1], stage4_44[2], stage4_44[3], stage4_44[4]},
      {1'b0},
      {stage4_46[0], stage4_46[1], stage4_46[2], stage4_46[3], stage4_46[4], stage4_46[5]},
      {stage5_48[0],stage5_47[1],stage5_46[1],stage5_45[1],stage5_44[2]}
   );
   gpc615_5 gpc2869 (
      {stage4_47[0], stage4_47[1], stage4_47[2], stage4_47[3], stage4_47[4]},
      {stage4_48[0]},
      {stage4_49[0], stage4_49[1], stage4_49[2], stage4_49[3], stage4_49[4], stage4_49[5]},
      {stage5_51[0],stage5_50[0],stage5_49[0],stage5_48[1],stage5_47[2]}
   );
   gpc117_4 gpc2870 (
      {stage4_50[0], stage4_50[1], stage4_50[2], stage4_50[3], stage4_50[4], stage4_50[5], stage4_50[6]},
      {stage4_51[0]},
      {stage4_52[0]},
      {stage5_53[0],stage5_52[0],stage5_51[1],stage5_50[1]}
   );
   gpc615_5 gpc2871 (
      {stage4_51[1], stage4_51[2], 1'b0, 1'b0, 1'b0},
      {stage4_52[1]},
      {stage4_53[0], stage4_53[1], stage4_53[2], stage4_53[3], stage4_53[4], stage4_53[5]},
      {stage5_55[0],stage5_54[0],stage5_53[1],stage5_52[1],stage5_51[2]}
   );
   gpc606_5 gpc2872 (
      {stage4_52[2], stage4_52[3], stage4_52[4], stage4_52[5], stage4_52[6], stage4_52[7]},
      {stage4_54[0], stage4_54[1], stage4_54[2], stage4_54[3], stage4_54[4], stage4_54[5]},
      {stage5_56[0],stage5_55[1],stage5_54[1],stage5_53[2],stage5_52[2]}
   );
   gpc606_5 gpc2873 (
      {stage4_52[8], stage4_52[9], stage4_52[10], stage4_52[11], stage4_52[12], stage4_52[13]},
      {stage4_54[6], stage4_54[7], stage4_54[8], stage4_54[9], stage4_54[10], stage4_54[11]},
      {stage5_56[1],stage5_55[2],stage5_54[2],stage5_53[3],stage5_52[3]}
   );
   gpc1415_5 gpc2874 (
      {stage4_55[0], stage4_55[1], stage4_55[2], stage4_55[3], 1'b0},
      {stage4_56[0]},
      {stage4_57[0], stage4_57[1], stage4_57[2], stage4_57[3]},
      {stage4_58[0]},
      {stage5_59[0],stage5_58[0],stage5_57[0],stage5_56[2],stage5_55[3]}
   );
   gpc135_4 gpc2875 (
      {stage4_56[1], stage4_56[2], stage4_56[3], stage4_56[4], stage4_56[5]},
      {stage4_57[4], stage4_57[5], 1'b0},
      {stage4_58[1]},
      {stage5_59[1],stage5_58[1],stage5_57[1],stage5_56[3]}
   );
   gpc606_5 gpc2876 (
      {stage4_59[0], stage4_59[1], stage4_59[2], stage4_59[3], stage4_59[4], stage4_59[5]},
      {stage4_61[0], stage4_61[1], stage4_61[2], stage4_61[3], stage4_61[4], stage4_61[5]},
      {stage5_63[0],stage5_62[0],stage5_61[0],stage5_60[0],stage5_59[2]}
   );
   gpc606_5 gpc2877 (
      {stage4_60[0], stage4_60[1], stage4_60[2], stage4_60[3], stage4_60[4], stage4_60[5]},
      {stage4_62[0], stage4_62[1], stage4_62[2], stage4_62[3], stage4_62[4], stage4_62[5]},
      {stage5_64[0],stage5_63[1],stage5_62[1],stage5_61[1],stage5_60[1]}
   );
   gpc1325_5 gpc2878 (
      {stage4_61[6], stage4_61[7], stage4_61[8], stage4_61[9], 1'b0},
      {1'b0, 1'b0},
      {stage4_63[0], stage4_63[1], stage4_63[2]},
      {stage4_64[0]},
      {stage5_65[0],stage5_64[1],stage5_63[2],stage5_62[2],stage5_61[2]}
   );
   gpc606_5 gpc2879 (
      {stage4_63[3], stage4_63[4], stage4_63[5], stage4_63[6], stage4_63[7], stage4_63[8]},
      {stage4_65[0], stage4_65[1], stage4_65[2], stage4_65[3], stage4_65[4], 1'b0},
      {stage5_67[0],stage5_66[0],stage5_65[1],stage5_64[2],stage5_63[3]}
   );
   gpc606_5 gpc2880 (
      {stage4_64[1], stage4_64[2], stage4_64[3], stage4_64[4], stage4_64[5], stage4_64[6]},
      {stage4_66[0], stage4_66[1], stage4_66[2], stage4_66[3], stage4_66[4], 1'b0},
      {stage5_68[0],stage5_67[1],stage5_66[1],stage5_65[2],stage5_64[3]}
   );
   gpc2135_5 gpc2881 (
      {stage4_67[0], stage4_67[1], stage4_67[2], stage4_67[3], 1'b0},
      {stage4_68[0], stage4_68[1], 1'b0},
      {stage4_69[0]},
      {1'b0, 1'b0},
      {stage5_70[0],stage5_69[0],stage5_68[1],stage5_67[2]}
   );
   gpc1_1 gpc2882 (
      {stage4_0[0]},
      {stage5_0[0]}
   );
   gpc1_1 gpc2883 (
      {stage4_1[0]},
      {stage5_1[0]}
   );
   gpc1_1 gpc2884 (
      {stage4_1[1]},
      {stage5_1[1]}
   );
   gpc1_1 gpc2885 (
      {stage4_2[0]},
      {stage5_2[0]}
   );
   gpc1_1 gpc2886 (
      {stage4_2[1]},
      {stage5_2[1]}
   );
   gpc1_1 gpc2887 (
      {stage4_3[7]},
      {stage5_3[1]}
   );
   gpc1_1 gpc2888 (
      {stage4_3[8]},
      {stage5_3[2]}
   );
   gpc1_1 gpc2889 (
      {stage4_3[9]},
      {stage5_3[3]}
   );
   gpc1_1 gpc2890 (
      {stage4_4[12]},
      {stage5_4[3]}
   );
   gpc1_1 gpc2891 (
      {stage4_4[13]},
      {stage5_4[4]}
   );
   gpc1_1 gpc2892 (
      {stage4_9[6]},
      {stage5_9[3]}
   );
   gpc1_1 gpc2893 (
      {stage4_10[6]},
      {stage5_10[2]}
   );
   gpc1_1 gpc2894 (
      {stage4_10[7]},
      {stage5_10[3]}
   );
   gpc1_1 gpc2895 (
      {stage4_10[8]},
      {stage5_10[4]}
   );
   gpc1_1 gpc2896 (
      {stage4_10[9]},
      {stage5_10[5]}
   );
   gpc1_1 gpc2897 (
      {stage4_10[10]},
      {stage5_10[6]}
   );
   gpc1_1 gpc2898 (
      {stage4_12[3]},
      {stage5_12[3]}
   );
   gpc1_1 gpc2899 (
      {stage4_12[4]},
      {stage5_12[4]}
   );
   gpc1_1 gpc2900 (
      {stage4_12[5]},
      {stage5_12[5]}
   );
   gpc1_1 gpc2901 (
      {stage4_13[2]},
      {stage5_13[2]}
   );
   gpc1_1 gpc2902 (
      {stage4_13[3]},
      {stage5_13[3]}
   );
   gpc1_1 gpc2903 (
      {stage4_13[4]},
      {stage5_13[4]}
   );
   gpc1_1 gpc2904 (
      {stage4_15[0]},
      {stage5_15[1]}
   );
   gpc1_1 gpc2905 (
      {stage4_15[1]},
      {stage5_15[2]}
   );
   gpc1_1 gpc2906 (
      {stage4_15[2]},
      {stage5_15[3]}
   );
   gpc1_1 gpc2907 (
      {stage4_15[3]},
      {stage5_15[4]}
   );
   gpc1_1 gpc2908 (
      {stage4_15[4]},
      {stage5_15[5]}
   );
   gpc1_1 gpc2909 (
      {stage4_15[5]},
      {stage5_15[6]}
   );
   gpc1_1 gpc2910 (
      {stage4_15[6]},
      {stage5_15[7]}
   );
   gpc1_1 gpc2911 (
      {stage4_15[7]},
      {stage5_15[8]}
   );
   gpc1_1 gpc2912 (
      {stage4_16[5]},
      {stage5_16[2]}
   );
   gpc1_1 gpc2913 (
      {stage4_16[6]},
      {stage5_16[3]}
   );
   gpc1_1 gpc2914 (
      {stage4_17[7]},
      {stage5_17[2]}
   );
   gpc1_1 gpc2915 (
      {stage4_19[6]},
      {stage5_19[2]}
   );
   gpc1_1 gpc2916 (
      {stage4_20[5]},
      {stage5_20[3]}
   );
   gpc1_1 gpc2917 (
      {stage4_20[6]},
      {stage5_20[4]}
   );
   gpc1_1 gpc2918 (
      {stage4_20[7]},
      {stage5_20[5]}
   );
   gpc1_1 gpc2919 (
      {stage4_20[8]},
      {stage5_20[6]}
   );
   gpc1_1 gpc2920 (
      {stage4_20[9]},
      {stage5_20[7]}
   );
   gpc1_1 gpc2921 (
      {stage4_20[10]},
      {stage5_20[8]}
   );
   gpc1_1 gpc2922 (
      {stage4_21[1]},
      {stage5_21[2]}
   );
   gpc1_1 gpc2923 (
      {stage4_21[2]},
      {stage5_21[3]}
   );
   gpc1_1 gpc2924 (
      {stage4_21[3]},
      {stage5_21[4]}
   );
   gpc1_1 gpc2925 (
      {stage4_22[3]},
      {stage5_22[2]}
   );
   gpc1_1 gpc2926 (
      {stage4_22[4]},
      {stage5_22[3]}
   );
   gpc1_1 gpc2927 (
      {stage4_24[7]},
      {stage5_24[2]}
   );
   gpc1_1 gpc2928 (
      {stage4_24[8]},
      {stage5_24[3]}
   );
   gpc1_1 gpc2929 (
      {stage4_24[9]},
      {stage5_24[4]}
   );
   gpc1_1 gpc2930 (
      {stage4_24[10]},
      {stage5_24[5]}
   );
   gpc1_1 gpc2931 (
      {stage4_27[1]},
      {stage5_27[3]}
   );
   gpc1_1 gpc2932 (
      {stage4_27[2]},
      {stage5_27[4]}
   );
   gpc1_1 gpc2933 (
      {stage4_27[3]},
      {stage5_27[5]}
   );
   gpc1_1 gpc2934 (
      {stage4_27[4]},
      {stage5_27[6]}
   );
   gpc1_1 gpc2935 (
      {stage4_27[5]},
      {stage5_27[7]}
   );
   gpc1_1 gpc2936 (
      {stage4_29[6]},
      {stage5_29[2]}
   );
   gpc1_1 gpc2937 (
      {stage4_29[7]},
      {stage5_29[3]}
   );
   gpc1_1 gpc2938 (
      {stage4_29[8]},
      {stage5_29[4]}
   );
   gpc1_1 gpc2939 (
      {stage4_29[9]},
      {stage5_29[5]}
   );
   gpc1_1 gpc2940 (
      {stage4_30[3]},
      {stage5_30[3]}
   );
   gpc1_1 gpc2941 (
      {stage4_32[6]},
      {stage5_32[2]}
   );
   gpc1_1 gpc2942 (
      {stage4_34[0]},
      {stage5_34[2]}
   );
   gpc1_1 gpc2943 (
      {stage4_34[1]},
      {stage5_34[3]}
   );
   gpc1_1 gpc2944 (
      {stage4_34[2]},
      {stage5_34[4]}
   );
   gpc1_1 gpc2945 (
      {stage4_34[3]},
      {stage5_34[5]}
   );
   gpc1_1 gpc2946 (
      {stage4_34[4]},
      {stage5_34[6]}
   );
   gpc1_1 gpc2947 (
      {stage4_34[5]},
      {stage5_34[7]}
   );
   gpc1_1 gpc2948 (
      {stage4_38[5]},
      {stage5_38[3]}
   );
   gpc1_1 gpc2949 (
      {stage4_39[6]},
      {stage5_39[3]}
   );
   gpc1_1 gpc2950 (
      {stage4_39[7]},
      {stage5_39[4]}
   );
   gpc1_1 gpc2951 (
      {stage4_44[5]},
      {stage5_44[3]}
   );
   gpc1_1 gpc2952 (
      {stage4_47[5]},
      {stage5_47[3]}
   );
   gpc1_1 gpc2953 (
      {stage4_47[6]},
      {stage5_47[4]}
   );
   gpc1_1 gpc2954 (
      {stage4_48[1]},
      {stage5_48[2]}
   );
   gpc1_1 gpc2955 (
      {stage4_48[2]},
      {stage5_48[3]}
   );
   gpc1_1 gpc2956 (
      {stage4_48[3]},
      {stage5_48[4]}
   );
   gpc1_1 gpc2957 (
      {stage4_48[4]},
      {stage5_48[5]}
   );
   gpc1_1 gpc2958 (
      {stage4_52[14]},
      {stage5_52[4]}
   );
   gpc1_1 gpc2959 (
      {stage4_52[15]},
      {stage5_52[5]}
   );
   gpc1_1 gpc2960 (
      {stage4_52[16]},
      {stage5_52[6]}
   );
   gpc1_1 gpc2961 (
      {stage4_56[6]},
      {stage5_56[4]}
   );
   gpc1_1 gpc2962 (
      {stage4_56[7]},
      {stage5_56[5]}
   );
   gpc1_1 gpc2963 (
      {stage4_58[2]},
      {stage5_58[2]}
   );
   gpc1_1 gpc2964 (
      {stage4_58[3]},
      {stage5_58[3]}
   );
   gpc1_1 gpc2965 (
      {stage4_64[7]},
      {stage5_64[4]}
   );
   gpc1_1 gpc2966 (
      {stage4_64[8]},
      {stage5_64[5]}
   );
   gpc1343_5 gpc2967 (
      {stage5_3[0], stage5_3[1], stage5_3[2]},
      {stage5_4[0], stage5_4[1], stage5_4[2], stage5_4[3]},
      {stage5_5[0], stage5_5[1], stage5_5[2]},
      {stage5_6[0]},
      {stage6_7[0],stage6_6[0],stage6_5[0],stage6_4[0],stage6_3[0]}
   );
   gpc135_4 gpc2968 (
      {stage5_6[1], stage5_6[2], stage5_6[3], 1'b0, 1'b0},
      {stage5_7[0], stage5_7[1], stage5_7[2]},
      {stage5_8[0]},
      {stage6_9[0],stage6_8[0],stage6_7[1],stage6_6[1]}
   );
   gpc1343_5 gpc2969 (
      {stage5_8[1], stage5_8[2], stage5_8[3]},
      {stage5_9[0], stage5_9[1], stage5_9[2], stage5_9[3]},
      {stage5_10[0], stage5_10[1], stage5_10[2]},
      {stage5_11[0]},
      {stage6_12[0],stage6_11[0],stage6_10[0],stage6_9[1],stage6_8[1]}
   );
   gpc615_5 gpc2970 (
      {stage5_10[3], stage5_10[4], stage5_10[5], stage5_10[6], 1'b0},
      {stage5_11[1]},
      {stage5_12[0], stage5_12[1], stage5_12[2], stage5_12[3], stage5_12[4], stage5_12[5]},
      {stage6_14[0],stage6_13[0],stage6_12[1],stage6_11[1],stage6_10[1]}
   );
   gpc615_5 gpc2971 (
      {stage5_13[0], stage5_13[1], stage5_13[2], stage5_13[3], stage5_13[4]},
      {stage5_14[0]},
      {stage5_15[0], stage5_15[1], stage5_15[2], stage5_15[3], stage5_15[4], stage5_15[5]},
      {stage6_17[0],stage6_16[0],stage6_15[0],stage6_14[1],stage6_13[1]}
   );
   gpc1343_5 gpc2972 (
      {stage5_15[6], stage5_15[7], stage5_15[8]},
      {stage5_16[0], stage5_16[1], stage5_16[2], stage5_16[3]},
      {stage5_17[0], stage5_17[1], stage5_17[2]},
      {stage5_18[0]},
      {stage6_19[0],stage6_18[0],stage6_17[1],stage6_16[1],stage6_15[1]}
   );
   gpc1163_5 gpc2973 (
      {stage5_19[0], stage5_19[1], stage5_19[2]},
      {stage5_20[0], stage5_20[1], stage5_20[2], stage5_20[3], stage5_20[4], stage5_20[5]},
      {stage5_21[0]},
      {stage5_22[0]},
      {stage6_23[0],stage6_22[0],stage6_21[0],stage6_20[0],stage6_19[1]}
   );
   gpc1343_5 gpc2974 (
      {stage5_20[6], stage5_20[7], stage5_20[8]},
      {stage5_21[1], stage5_21[2], stage5_21[3], stage5_21[4]},
      {stage5_22[1], stage5_22[2], stage5_22[3]},
      {stage5_23[0]},
      {stage6_24[0],stage6_23[1],stage6_22[1],stage6_21[1],stage6_20[1]}
   );
   gpc7_3 gpc2975 (
      {stage5_24[0], stage5_24[1], stage5_24[2], stage5_24[3], stage5_24[4], stage5_24[5], 1'b0},
      {stage6_26[0],stage6_25[0],stage6_24[1]}
   );
   gpc1343_5 gpc2976 (
      {stage5_25[0], stage5_25[1], stage5_25[2]},
      {stage5_26[0], stage5_26[1], stage5_26[2], stage5_26[3]},
      {stage5_27[0], stage5_27[1], stage5_27[2]},
      {stage5_28[0]},
      {stage6_29[0],stage6_28[0],stage6_27[0],stage6_26[1],stage6_25[1]}
   );
   gpc615_5 gpc2977 (
      {stage5_27[3], stage5_27[4], stage5_27[5], stage5_27[6], stage5_27[7]},
      {stage5_28[1]},
      {stage5_29[0], stage5_29[1], stage5_29[2], stage5_29[3], stage5_29[4], stage5_29[5]},
      {stage6_31[0],stage6_30[0],stage6_29[1],stage6_28[1],stage6_27[1]}
   );
   gpc135_4 gpc2978 (
      {stage5_30[0], stage5_30[1], stage5_30[2], stage5_30[3], 1'b0},
      {stage5_31[0], stage5_31[1], 1'b0},
      {stage5_32[0]},
      {stage6_33[0],stage6_32[0],stage6_31[1],stage6_30[1]}
   );
   gpc135_4 gpc2979 (
      {stage5_32[1], stage5_32[2], 1'b0, 1'b0, 1'b0},
      {stage5_33[0], stage5_33[1], stage5_33[2]},
      {stage5_34[0]},
      {stage6_35[0],stage6_34[0],stage6_33[1],stage6_32[1]}
   );
   gpc117_4 gpc2980 (
      {stage5_34[1], stage5_34[2], stage5_34[3], stage5_34[4], stage5_34[5], stage5_34[6], stage5_34[7]},
      {stage5_35[0]},
      {stage5_36[0]},
      {stage6_37[0],stage6_36[0],stage6_35[1],stage6_34[1]}
   );
   gpc1343_5 gpc2981 (
      {stage5_37[0], stage5_37[1], stage5_37[2]},
      {stage5_38[0], stage5_38[1], stage5_38[2], stage5_38[3]},
      {stage5_39[0], stage5_39[1], stage5_39[2]},
      {stage5_40[0]},
      {stage6_41[0],stage6_40[0],stage6_39[0],stage6_38[0],stage6_37[1]}
   );
   gpc1423_5 gpc2982 (
      {stage5_39[3], stage5_39[4], 1'b0},
      {stage5_40[1], stage5_40[2]},
      {stage5_41[0], stage5_41[1], stage5_41[2], stage5_41[3]},
      {stage5_42[0]},
      {stage6_43[0],stage6_42[0],stage6_41[1],stage6_40[1],stage6_39[1]}
   );
   gpc1343_5 gpc2983 (
      {stage5_42[1], stage5_42[2], stage5_42[3]},
      {stage5_43[0], stage5_43[1], stage5_43[2], stage5_43[3]},
      {stage5_44[0], stage5_44[1], stage5_44[2]},
      {stage5_45[0]},
      {stage6_46[0],stage6_45[0],stage6_44[0],stage6_43[1],stage6_42[1]}
   );
   gpc1343_5 gpc2984 (
      {stage5_46[0], stage5_46[1], 1'b0},
      {stage5_47[0], stage5_47[1], stage5_47[2], stage5_47[3]},
      {stage5_48[0], stage5_48[1], stage5_48[2]},
      {stage5_49[0]},
      {stage6_50[0],stage6_49[0],stage6_48[0],stage6_47[0],stage6_46[1]}
   );
   gpc223_4 gpc2985 (
      {stage5_48[3], stage5_48[4], stage5_48[5]},
      {1'b0, 1'b0},
      {stage5_50[0], stage5_50[1]},
      {stage6_51[0],stage6_50[1],stage6_49[1],stage6_48[1]}
   );
   gpc223_4 gpc2986 (
      {stage5_51[0], stage5_51[1], stage5_51[2]},
      {stage5_52[0], stage5_52[1]},
      {stage5_53[0], stage5_53[1]},
      {stage6_54[0],stage6_53[0],stage6_52[0],stage6_51[1]}
   );
   gpc1325_5 gpc2987 (
      {stage5_52[2], stage5_52[3], stage5_52[4], stage5_52[5], stage5_52[6]},
      {stage5_53[2], stage5_53[3]},
      {stage5_54[0], stage5_54[1], stage5_54[2]},
      {stage5_55[0]},
      {stage6_56[0],stage6_55[0],stage6_54[1],stage6_53[1],stage6_52[1]}
   );
   gpc1163_5 gpc2988 (
      {stage5_55[1], stage5_55[2], stage5_55[3]},
      {stage5_56[0], stage5_56[1], stage5_56[2], stage5_56[3], stage5_56[4], stage5_56[5]},
      {stage5_57[0]},
      {stage5_58[0]},
      {stage6_59[0],stage6_58[0],stage6_57[0],stage6_56[1],stage6_55[1]}
   );
   gpc1343_5 gpc2989 (
      {stage5_57[1], 1'b0, 1'b0},
      {stage5_58[1], stage5_58[2], stage5_58[3], 1'b0},
      {stage5_59[0], stage5_59[1], stage5_59[2]},
      {stage5_60[0]},
      {stage6_61[0],stage6_60[0],stage6_59[1],stage6_58[1],stage6_57[1]}
   );
   gpc1423_5 gpc2990 (
      {stage5_61[0], stage5_61[1], stage5_61[2]},
      {stage5_62[0], stage5_62[1]},
      {stage5_63[0], stage5_63[1], stage5_63[2], stage5_63[3]},
      {stage5_64[0]},
      {stage6_65[0],stage6_64[0],stage6_63[0],stage6_62[0],stage6_61[1]}
   );
   gpc135_4 gpc2991 (
      {stage5_64[1], stage5_64[2], stage5_64[3], stage5_64[4], stage5_64[5]},
      {stage5_65[0], stage5_65[1], stage5_65[2]},
      {stage5_66[0]},
      {stage6_67[0],stage6_66[0],stage6_65[1],stage6_64[1]}
   );
   gpc1163_5 gpc2992 (
      {stage5_66[1], 1'b0, 1'b0},
      {stage5_67[0], stage5_67[1], stage5_67[2], 1'b0, 1'b0, 1'b0},
      {stage5_68[0]},
      {stage5_69[0]},
      {stage6_70[0],stage6_69[0],stage6_68[0],stage6_67[1],stage6_66[1]}
   );
   gpc1_1 gpc2993 (
      {stage5_0[0]},
      {stage6_0[0]}
   );
   gpc1_1 gpc2994 (
      {stage5_1[0]},
      {stage6_1[0]}
   );
   gpc1_1 gpc2995 (
      {stage5_1[1]},
      {stage6_1[1]}
   );
   gpc1_1 gpc2996 (
      {stage5_2[0]},
      {stage6_2[0]}
   );
   gpc1_1 gpc2997 (
      {stage5_2[1]},
      {stage6_2[1]}
   );
   gpc1_1 gpc2998 (
      {stage5_3[3]},
      {stage6_3[1]}
   );
   gpc1_1 gpc2999 (
      {stage5_4[4]},
      {stage6_4[1]}
   );
   gpc1_1 gpc3000 (
      {stage5_5[3]},
      {stage6_5[1]}
   );
   gpc1_1 gpc3001 (
      {stage5_18[1]},
      {stage6_18[1]}
   );
   gpc1_1 gpc3002 (
      {stage5_36[1]},
      {stage6_36[1]}
   );
   gpc1_1 gpc3003 (
      {stage5_44[3]},
      {stage6_44[1]}
   );
   gpc1_1 gpc3004 (
      {stage5_45[1]},
      {stage6_45[1]}
   );
   gpc1_1 gpc3005 (
      {stage5_47[4]},
      {stage6_47[1]}
   );
   gpc1_1 gpc3006 (
      {stage5_60[1]},
      {stage6_60[1]}
   );
   gpc1_1 gpc3007 (
      {stage5_62[2]},
      {stage6_62[1]}
   );
   gpc1_1 gpc3008 (
      {stage5_68[1]},
      {stage6_68[1]}
   );
   gpc1_1 gpc3009 (
      {stage5_70[0]},
      {stage6_70[1]}
   );
endmodule

module testbench();
    reg [127:0] src0;
    reg [127:0] src1;
    reg [127:0] src2;
    reg [127:0] src3;
    reg [127:0] src4;
    reg [127:0] src5;
    reg [127:0] src6;
    reg [127:0] src7;
    reg [127:0] src8;
    reg [127:0] src9;
    reg [127:0] src10;
    reg [127:0] src11;
    reg [127:0] src12;
    reg [127:0] src13;
    reg [127:0] src14;
    reg [127:0] src15;
    reg [127:0] src16;
    reg [127:0] src17;
    reg [127:0] src18;
    reg [127:0] src19;
    reg [127:0] src20;
    reg [127:0] src21;
    reg [127:0] src22;
    reg [127:0] src23;
    reg [127:0] src24;
    reg [127:0] src25;
    reg [127:0] src26;
    reg [127:0] src27;
    reg [127:0] src28;
    reg [127:0] src29;
    reg [127:0] src30;
    reg [127:0] src31;
    reg [127:0] src32;
    reg [127:0] src33;
    reg [127:0] src34;
    reg [127:0] src35;
    reg [127:0] src36;
    reg [127:0] src37;
    reg [127:0] src38;
    reg [127:0] src39;
    reg [127:0] src40;
    reg [127:0] src41;
    reg [127:0] src42;
    reg [127:0] src43;
    reg [127:0] src44;
    reg [127:0] src45;
    reg [127:0] src46;
    reg [127:0] src47;
    reg [127:0] src48;
    reg [127:0] src49;
    reg [127:0] src50;
    reg [127:0] src51;
    reg [127:0] src52;
    reg [127:0] src53;
    reg [127:0] src54;
    reg [127:0] src55;
    reg [127:0] src56;
    reg [127:0] src57;
    reg [127:0] src58;
    reg [127:0] src59;
    reg [127:0] src60;
    reg [127:0] src61;
    reg [127:0] src62;
    reg [127:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [0:0] dst69;
    wire [0:0] dst70;
    wire [70:0] srcsum;
    wire [70:0] dstsum;
    wire test;
    compressor_CLA128_64 compressor_CLA128_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68),
        .dst69(dst69),
        .dst70(dst70));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31] + src0[32] + src0[33] + src0[34] + src0[35] + src0[36] + src0[37] + src0[38] + src0[39] + src0[40] + src0[41] + src0[42] + src0[43] + src0[44] + src0[45] + src0[46] + src0[47] + src0[48] + src0[49] + src0[50] + src0[51] + src0[52] + src0[53] + src0[54] + src0[55] + src0[56] + src0[57] + src0[58] + src0[59] + src0[60] + src0[61] + src0[62] + src0[63] + src0[64] + src0[65] + src0[66] + src0[67] + src0[68] + src0[69] + src0[70] + src0[71] + src0[72] + src0[73] + src0[74] + src0[75] + src0[76] + src0[77] + src0[78] + src0[79] + src0[80] + src0[81] + src0[82] + src0[83] + src0[84] + src0[85] + src0[86] + src0[87] + src0[88] + src0[89] + src0[90] + src0[91] + src0[92] + src0[93] + src0[94] + src0[95] + src0[96] + src0[97] + src0[98] + src0[99] + src0[100] + src0[101] + src0[102] + src0[103] + src0[104] + src0[105] + src0[106] + src0[107] + src0[108] + src0[109] + src0[110] + src0[111] + src0[112] + src0[113] + src0[114] + src0[115] + src0[116] + src0[117] + src0[118] + src0[119] + src0[120] + src0[121] + src0[122] + src0[123] + src0[124] + src0[125] + src0[126] + src0[127])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31] + src1[32] + src1[33] + src1[34] + src1[35] + src1[36] + src1[37] + src1[38] + src1[39] + src1[40] + src1[41] + src1[42] + src1[43] + src1[44] + src1[45] + src1[46] + src1[47] + src1[48] + src1[49] + src1[50] + src1[51] + src1[52] + src1[53] + src1[54] + src1[55] + src1[56] + src1[57] + src1[58] + src1[59] + src1[60] + src1[61] + src1[62] + src1[63] + src1[64] + src1[65] + src1[66] + src1[67] + src1[68] + src1[69] + src1[70] + src1[71] + src1[72] + src1[73] + src1[74] + src1[75] + src1[76] + src1[77] + src1[78] + src1[79] + src1[80] + src1[81] + src1[82] + src1[83] + src1[84] + src1[85] + src1[86] + src1[87] + src1[88] + src1[89] + src1[90] + src1[91] + src1[92] + src1[93] + src1[94] + src1[95] + src1[96] + src1[97] + src1[98] + src1[99] + src1[100] + src1[101] + src1[102] + src1[103] + src1[104] + src1[105] + src1[106] + src1[107] + src1[108] + src1[109] + src1[110] + src1[111] + src1[112] + src1[113] + src1[114] + src1[115] + src1[116] + src1[117] + src1[118] + src1[119] + src1[120] + src1[121] + src1[122] + src1[123] + src1[124] + src1[125] + src1[126] + src1[127])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31] + src2[32] + src2[33] + src2[34] + src2[35] + src2[36] + src2[37] + src2[38] + src2[39] + src2[40] + src2[41] + src2[42] + src2[43] + src2[44] + src2[45] + src2[46] + src2[47] + src2[48] + src2[49] + src2[50] + src2[51] + src2[52] + src2[53] + src2[54] + src2[55] + src2[56] + src2[57] + src2[58] + src2[59] + src2[60] + src2[61] + src2[62] + src2[63] + src2[64] + src2[65] + src2[66] + src2[67] + src2[68] + src2[69] + src2[70] + src2[71] + src2[72] + src2[73] + src2[74] + src2[75] + src2[76] + src2[77] + src2[78] + src2[79] + src2[80] + src2[81] + src2[82] + src2[83] + src2[84] + src2[85] + src2[86] + src2[87] + src2[88] + src2[89] + src2[90] + src2[91] + src2[92] + src2[93] + src2[94] + src2[95] + src2[96] + src2[97] + src2[98] + src2[99] + src2[100] + src2[101] + src2[102] + src2[103] + src2[104] + src2[105] + src2[106] + src2[107] + src2[108] + src2[109] + src2[110] + src2[111] + src2[112] + src2[113] + src2[114] + src2[115] + src2[116] + src2[117] + src2[118] + src2[119] + src2[120] + src2[121] + src2[122] + src2[123] + src2[124] + src2[125] + src2[126] + src2[127])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31] + src3[32] + src3[33] + src3[34] + src3[35] + src3[36] + src3[37] + src3[38] + src3[39] + src3[40] + src3[41] + src3[42] + src3[43] + src3[44] + src3[45] + src3[46] + src3[47] + src3[48] + src3[49] + src3[50] + src3[51] + src3[52] + src3[53] + src3[54] + src3[55] + src3[56] + src3[57] + src3[58] + src3[59] + src3[60] + src3[61] + src3[62] + src3[63] + src3[64] + src3[65] + src3[66] + src3[67] + src3[68] + src3[69] + src3[70] + src3[71] + src3[72] + src3[73] + src3[74] + src3[75] + src3[76] + src3[77] + src3[78] + src3[79] + src3[80] + src3[81] + src3[82] + src3[83] + src3[84] + src3[85] + src3[86] + src3[87] + src3[88] + src3[89] + src3[90] + src3[91] + src3[92] + src3[93] + src3[94] + src3[95] + src3[96] + src3[97] + src3[98] + src3[99] + src3[100] + src3[101] + src3[102] + src3[103] + src3[104] + src3[105] + src3[106] + src3[107] + src3[108] + src3[109] + src3[110] + src3[111] + src3[112] + src3[113] + src3[114] + src3[115] + src3[116] + src3[117] + src3[118] + src3[119] + src3[120] + src3[121] + src3[122] + src3[123] + src3[124] + src3[125] + src3[126] + src3[127])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31] + src4[32] + src4[33] + src4[34] + src4[35] + src4[36] + src4[37] + src4[38] + src4[39] + src4[40] + src4[41] + src4[42] + src4[43] + src4[44] + src4[45] + src4[46] + src4[47] + src4[48] + src4[49] + src4[50] + src4[51] + src4[52] + src4[53] + src4[54] + src4[55] + src4[56] + src4[57] + src4[58] + src4[59] + src4[60] + src4[61] + src4[62] + src4[63] + src4[64] + src4[65] + src4[66] + src4[67] + src4[68] + src4[69] + src4[70] + src4[71] + src4[72] + src4[73] + src4[74] + src4[75] + src4[76] + src4[77] + src4[78] + src4[79] + src4[80] + src4[81] + src4[82] + src4[83] + src4[84] + src4[85] + src4[86] + src4[87] + src4[88] + src4[89] + src4[90] + src4[91] + src4[92] + src4[93] + src4[94] + src4[95] + src4[96] + src4[97] + src4[98] + src4[99] + src4[100] + src4[101] + src4[102] + src4[103] + src4[104] + src4[105] + src4[106] + src4[107] + src4[108] + src4[109] + src4[110] + src4[111] + src4[112] + src4[113] + src4[114] + src4[115] + src4[116] + src4[117] + src4[118] + src4[119] + src4[120] + src4[121] + src4[122] + src4[123] + src4[124] + src4[125] + src4[126] + src4[127])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31] + src5[32] + src5[33] + src5[34] + src5[35] + src5[36] + src5[37] + src5[38] + src5[39] + src5[40] + src5[41] + src5[42] + src5[43] + src5[44] + src5[45] + src5[46] + src5[47] + src5[48] + src5[49] + src5[50] + src5[51] + src5[52] + src5[53] + src5[54] + src5[55] + src5[56] + src5[57] + src5[58] + src5[59] + src5[60] + src5[61] + src5[62] + src5[63] + src5[64] + src5[65] + src5[66] + src5[67] + src5[68] + src5[69] + src5[70] + src5[71] + src5[72] + src5[73] + src5[74] + src5[75] + src5[76] + src5[77] + src5[78] + src5[79] + src5[80] + src5[81] + src5[82] + src5[83] + src5[84] + src5[85] + src5[86] + src5[87] + src5[88] + src5[89] + src5[90] + src5[91] + src5[92] + src5[93] + src5[94] + src5[95] + src5[96] + src5[97] + src5[98] + src5[99] + src5[100] + src5[101] + src5[102] + src5[103] + src5[104] + src5[105] + src5[106] + src5[107] + src5[108] + src5[109] + src5[110] + src5[111] + src5[112] + src5[113] + src5[114] + src5[115] + src5[116] + src5[117] + src5[118] + src5[119] + src5[120] + src5[121] + src5[122] + src5[123] + src5[124] + src5[125] + src5[126] + src5[127])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31] + src6[32] + src6[33] + src6[34] + src6[35] + src6[36] + src6[37] + src6[38] + src6[39] + src6[40] + src6[41] + src6[42] + src6[43] + src6[44] + src6[45] + src6[46] + src6[47] + src6[48] + src6[49] + src6[50] + src6[51] + src6[52] + src6[53] + src6[54] + src6[55] + src6[56] + src6[57] + src6[58] + src6[59] + src6[60] + src6[61] + src6[62] + src6[63] + src6[64] + src6[65] + src6[66] + src6[67] + src6[68] + src6[69] + src6[70] + src6[71] + src6[72] + src6[73] + src6[74] + src6[75] + src6[76] + src6[77] + src6[78] + src6[79] + src6[80] + src6[81] + src6[82] + src6[83] + src6[84] + src6[85] + src6[86] + src6[87] + src6[88] + src6[89] + src6[90] + src6[91] + src6[92] + src6[93] + src6[94] + src6[95] + src6[96] + src6[97] + src6[98] + src6[99] + src6[100] + src6[101] + src6[102] + src6[103] + src6[104] + src6[105] + src6[106] + src6[107] + src6[108] + src6[109] + src6[110] + src6[111] + src6[112] + src6[113] + src6[114] + src6[115] + src6[116] + src6[117] + src6[118] + src6[119] + src6[120] + src6[121] + src6[122] + src6[123] + src6[124] + src6[125] + src6[126] + src6[127])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31] + src7[32] + src7[33] + src7[34] + src7[35] + src7[36] + src7[37] + src7[38] + src7[39] + src7[40] + src7[41] + src7[42] + src7[43] + src7[44] + src7[45] + src7[46] + src7[47] + src7[48] + src7[49] + src7[50] + src7[51] + src7[52] + src7[53] + src7[54] + src7[55] + src7[56] + src7[57] + src7[58] + src7[59] + src7[60] + src7[61] + src7[62] + src7[63] + src7[64] + src7[65] + src7[66] + src7[67] + src7[68] + src7[69] + src7[70] + src7[71] + src7[72] + src7[73] + src7[74] + src7[75] + src7[76] + src7[77] + src7[78] + src7[79] + src7[80] + src7[81] + src7[82] + src7[83] + src7[84] + src7[85] + src7[86] + src7[87] + src7[88] + src7[89] + src7[90] + src7[91] + src7[92] + src7[93] + src7[94] + src7[95] + src7[96] + src7[97] + src7[98] + src7[99] + src7[100] + src7[101] + src7[102] + src7[103] + src7[104] + src7[105] + src7[106] + src7[107] + src7[108] + src7[109] + src7[110] + src7[111] + src7[112] + src7[113] + src7[114] + src7[115] + src7[116] + src7[117] + src7[118] + src7[119] + src7[120] + src7[121] + src7[122] + src7[123] + src7[124] + src7[125] + src7[126] + src7[127])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31] + src8[32] + src8[33] + src8[34] + src8[35] + src8[36] + src8[37] + src8[38] + src8[39] + src8[40] + src8[41] + src8[42] + src8[43] + src8[44] + src8[45] + src8[46] + src8[47] + src8[48] + src8[49] + src8[50] + src8[51] + src8[52] + src8[53] + src8[54] + src8[55] + src8[56] + src8[57] + src8[58] + src8[59] + src8[60] + src8[61] + src8[62] + src8[63] + src8[64] + src8[65] + src8[66] + src8[67] + src8[68] + src8[69] + src8[70] + src8[71] + src8[72] + src8[73] + src8[74] + src8[75] + src8[76] + src8[77] + src8[78] + src8[79] + src8[80] + src8[81] + src8[82] + src8[83] + src8[84] + src8[85] + src8[86] + src8[87] + src8[88] + src8[89] + src8[90] + src8[91] + src8[92] + src8[93] + src8[94] + src8[95] + src8[96] + src8[97] + src8[98] + src8[99] + src8[100] + src8[101] + src8[102] + src8[103] + src8[104] + src8[105] + src8[106] + src8[107] + src8[108] + src8[109] + src8[110] + src8[111] + src8[112] + src8[113] + src8[114] + src8[115] + src8[116] + src8[117] + src8[118] + src8[119] + src8[120] + src8[121] + src8[122] + src8[123] + src8[124] + src8[125] + src8[126] + src8[127])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31] + src9[32] + src9[33] + src9[34] + src9[35] + src9[36] + src9[37] + src9[38] + src9[39] + src9[40] + src9[41] + src9[42] + src9[43] + src9[44] + src9[45] + src9[46] + src9[47] + src9[48] + src9[49] + src9[50] + src9[51] + src9[52] + src9[53] + src9[54] + src9[55] + src9[56] + src9[57] + src9[58] + src9[59] + src9[60] + src9[61] + src9[62] + src9[63] + src9[64] + src9[65] + src9[66] + src9[67] + src9[68] + src9[69] + src9[70] + src9[71] + src9[72] + src9[73] + src9[74] + src9[75] + src9[76] + src9[77] + src9[78] + src9[79] + src9[80] + src9[81] + src9[82] + src9[83] + src9[84] + src9[85] + src9[86] + src9[87] + src9[88] + src9[89] + src9[90] + src9[91] + src9[92] + src9[93] + src9[94] + src9[95] + src9[96] + src9[97] + src9[98] + src9[99] + src9[100] + src9[101] + src9[102] + src9[103] + src9[104] + src9[105] + src9[106] + src9[107] + src9[108] + src9[109] + src9[110] + src9[111] + src9[112] + src9[113] + src9[114] + src9[115] + src9[116] + src9[117] + src9[118] + src9[119] + src9[120] + src9[121] + src9[122] + src9[123] + src9[124] + src9[125] + src9[126] + src9[127])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31] + src10[32] + src10[33] + src10[34] + src10[35] + src10[36] + src10[37] + src10[38] + src10[39] + src10[40] + src10[41] + src10[42] + src10[43] + src10[44] + src10[45] + src10[46] + src10[47] + src10[48] + src10[49] + src10[50] + src10[51] + src10[52] + src10[53] + src10[54] + src10[55] + src10[56] + src10[57] + src10[58] + src10[59] + src10[60] + src10[61] + src10[62] + src10[63] + src10[64] + src10[65] + src10[66] + src10[67] + src10[68] + src10[69] + src10[70] + src10[71] + src10[72] + src10[73] + src10[74] + src10[75] + src10[76] + src10[77] + src10[78] + src10[79] + src10[80] + src10[81] + src10[82] + src10[83] + src10[84] + src10[85] + src10[86] + src10[87] + src10[88] + src10[89] + src10[90] + src10[91] + src10[92] + src10[93] + src10[94] + src10[95] + src10[96] + src10[97] + src10[98] + src10[99] + src10[100] + src10[101] + src10[102] + src10[103] + src10[104] + src10[105] + src10[106] + src10[107] + src10[108] + src10[109] + src10[110] + src10[111] + src10[112] + src10[113] + src10[114] + src10[115] + src10[116] + src10[117] + src10[118] + src10[119] + src10[120] + src10[121] + src10[122] + src10[123] + src10[124] + src10[125] + src10[126] + src10[127])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31] + src11[32] + src11[33] + src11[34] + src11[35] + src11[36] + src11[37] + src11[38] + src11[39] + src11[40] + src11[41] + src11[42] + src11[43] + src11[44] + src11[45] + src11[46] + src11[47] + src11[48] + src11[49] + src11[50] + src11[51] + src11[52] + src11[53] + src11[54] + src11[55] + src11[56] + src11[57] + src11[58] + src11[59] + src11[60] + src11[61] + src11[62] + src11[63] + src11[64] + src11[65] + src11[66] + src11[67] + src11[68] + src11[69] + src11[70] + src11[71] + src11[72] + src11[73] + src11[74] + src11[75] + src11[76] + src11[77] + src11[78] + src11[79] + src11[80] + src11[81] + src11[82] + src11[83] + src11[84] + src11[85] + src11[86] + src11[87] + src11[88] + src11[89] + src11[90] + src11[91] + src11[92] + src11[93] + src11[94] + src11[95] + src11[96] + src11[97] + src11[98] + src11[99] + src11[100] + src11[101] + src11[102] + src11[103] + src11[104] + src11[105] + src11[106] + src11[107] + src11[108] + src11[109] + src11[110] + src11[111] + src11[112] + src11[113] + src11[114] + src11[115] + src11[116] + src11[117] + src11[118] + src11[119] + src11[120] + src11[121] + src11[122] + src11[123] + src11[124] + src11[125] + src11[126] + src11[127])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31] + src12[32] + src12[33] + src12[34] + src12[35] + src12[36] + src12[37] + src12[38] + src12[39] + src12[40] + src12[41] + src12[42] + src12[43] + src12[44] + src12[45] + src12[46] + src12[47] + src12[48] + src12[49] + src12[50] + src12[51] + src12[52] + src12[53] + src12[54] + src12[55] + src12[56] + src12[57] + src12[58] + src12[59] + src12[60] + src12[61] + src12[62] + src12[63] + src12[64] + src12[65] + src12[66] + src12[67] + src12[68] + src12[69] + src12[70] + src12[71] + src12[72] + src12[73] + src12[74] + src12[75] + src12[76] + src12[77] + src12[78] + src12[79] + src12[80] + src12[81] + src12[82] + src12[83] + src12[84] + src12[85] + src12[86] + src12[87] + src12[88] + src12[89] + src12[90] + src12[91] + src12[92] + src12[93] + src12[94] + src12[95] + src12[96] + src12[97] + src12[98] + src12[99] + src12[100] + src12[101] + src12[102] + src12[103] + src12[104] + src12[105] + src12[106] + src12[107] + src12[108] + src12[109] + src12[110] + src12[111] + src12[112] + src12[113] + src12[114] + src12[115] + src12[116] + src12[117] + src12[118] + src12[119] + src12[120] + src12[121] + src12[122] + src12[123] + src12[124] + src12[125] + src12[126] + src12[127])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31] + src13[32] + src13[33] + src13[34] + src13[35] + src13[36] + src13[37] + src13[38] + src13[39] + src13[40] + src13[41] + src13[42] + src13[43] + src13[44] + src13[45] + src13[46] + src13[47] + src13[48] + src13[49] + src13[50] + src13[51] + src13[52] + src13[53] + src13[54] + src13[55] + src13[56] + src13[57] + src13[58] + src13[59] + src13[60] + src13[61] + src13[62] + src13[63] + src13[64] + src13[65] + src13[66] + src13[67] + src13[68] + src13[69] + src13[70] + src13[71] + src13[72] + src13[73] + src13[74] + src13[75] + src13[76] + src13[77] + src13[78] + src13[79] + src13[80] + src13[81] + src13[82] + src13[83] + src13[84] + src13[85] + src13[86] + src13[87] + src13[88] + src13[89] + src13[90] + src13[91] + src13[92] + src13[93] + src13[94] + src13[95] + src13[96] + src13[97] + src13[98] + src13[99] + src13[100] + src13[101] + src13[102] + src13[103] + src13[104] + src13[105] + src13[106] + src13[107] + src13[108] + src13[109] + src13[110] + src13[111] + src13[112] + src13[113] + src13[114] + src13[115] + src13[116] + src13[117] + src13[118] + src13[119] + src13[120] + src13[121] + src13[122] + src13[123] + src13[124] + src13[125] + src13[126] + src13[127])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31] + src14[32] + src14[33] + src14[34] + src14[35] + src14[36] + src14[37] + src14[38] + src14[39] + src14[40] + src14[41] + src14[42] + src14[43] + src14[44] + src14[45] + src14[46] + src14[47] + src14[48] + src14[49] + src14[50] + src14[51] + src14[52] + src14[53] + src14[54] + src14[55] + src14[56] + src14[57] + src14[58] + src14[59] + src14[60] + src14[61] + src14[62] + src14[63] + src14[64] + src14[65] + src14[66] + src14[67] + src14[68] + src14[69] + src14[70] + src14[71] + src14[72] + src14[73] + src14[74] + src14[75] + src14[76] + src14[77] + src14[78] + src14[79] + src14[80] + src14[81] + src14[82] + src14[83] + src14[84] + src14[85] + src14[86] + src14[87] + src14[88] + src14[89] + src14[90] + src14[91] + src14[92] + src14[93] + src14[94] + src14[95] + src14[96] + src14[97] + src14[98] + src14[99] + src14[100] + src14[101] + src14[102] + src14[103] + src14[104] + src14[105] + src14[106] + src14[107] + src14[108] + src14[109] + src14[110] + src14[111] + src14[112] + src14[113] + src14[114] + src14[115] + src14[116] + src14[117] + src14[118] + src14[119] + src14[120] + src14[121] + src14[122] + src14[123] + src14[124] + src14[125] + src14[126] + src14[127])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31] + src15[32] + src15[33] + src15[34] + src15[35] + src15[36] + src15[37] + src15[38] + src15[39] + src15[40] + src15[41] + src15[42] + src15[43] + src15[44] + src15[45] + src15[46] + src15[47] + src15[48] + src15[49] + src15[50] + src15[51] + src15[52] + src15[53] + src15[54] + src15[55] + src15[56] + src15[57] + src15[58] + src15[59] + src15[60] + src15[61] + src15[62] + src15[63] + src15[64] + src15[65] + src15[66] + src15[67] + src15[68] + src15[69] + src15[70] + src15[71] + src15[72] + src15[73] + src15[74] + src15[75] + src15[76] + src15[77] + src15[78] + src15[79] + src15[80] + src15[81] + src15[82] + src15[83] + src15[84] + src15[85] + src15[86] + src15[87] + src15[88] + src15[89] + src15[90] + src15[91] + src15[92] + src15[93] + src15[94] + src15[95] + src15[96] + src15[97] + src15[98] + src15[99] + src15[100] + src15[101] + src15[102] + src15[103] + src15[104] + src15[105] + src15[106] + src15[107] + src15[108] + src15[109] + src15[110] + src15[111] + src15[112] + src15[113] + src15[114] + src15[115] + src15[116] + src15[117] + src15[118] + src15[119] + src15[120] + src15[121] + src15[122] + src15[123] + src15[124] + src15[125] + src15[126] + src15[127])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31] + src16[32] + src16[33] + src16[34] + src16[35] + src16[36] + src16[37] + src16[38] + src16[39] + src16[40] + src16[41] + src16[42] + src16[43] + src16[44] + src16[45] + src16[46] + src16[47] + src16[48] + src16[49] + src16[50] + src16[51] + src16[52] + src16[53] + src16[54] + src16[55] + src16[56] + src16[57] + src16[58] + src16[59] + src16[60] + src16[61] + src16[62] + src16[63] + src16[64] + src16[65] + src16[66] + src16[67] + src16[68] + src16[69] + src16[70] + src16[71] + src16[72] + src16[73] + src16[74] + src16[75] + src16[76] + src16[77] + src16[78] + src16[79] + src16[80] + src16[81] + src16[82] + src16[83] + src16[84] + src16[85] + src16[86] + src16[87] + src16[88] + src16[89] + src16[90] + src16[91] + src16[92] + src16[93] + src16[94] + src16[95] + src16[96] + src16[97] + src16[98] + src16[99] + src16[100] + src16[101] + src16[102] + src16[103] + src16[104] + src16[105] + src16[106] + src16[107] + src16[108] + src16[109] + src16[110] + src16[111] + src16[112] + src16[113] + src16[114] + src16[115] + src16[116] + src16[117] + src16[118] + src16[119] + src16[120] + src16[121] + src16[122] + src16[123] + src16[124] + src16[125] + src16[126] + src16[127])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31] + src17[32] + src17[33] + src17[34] + src17[35] + src17[36] + src17[37] + src17[38] + src17[39] + src17[40] + src17[41] + src17[42] + src17[43] + src17[44] + src17[45] + src17[46] + src17[47] + src17[48] + src17[49] + src17[50] + src17[51] + src17[52] + src17[53] + src17[54] + src17[55] + src17[56] + src17[57] + src17[58] + src17[59] + src17[60] + src17[61] + src17[62] + src17[63] + src17[64] + src17[65] + src17[66] + src17[67] + src17[68] + src17[69] + src17[70] + src17[71] + src17[72] + src17[73] + src17[74] + src17[75] + src17[76] + src17[77] + src17[78] + src17[79] + src17[80] + src17[81] + src17[82] + src17[83] + src17[84] + src17[85] + src17[86] + src17[87] + src17[88] + src17[89] + src17[90] + src17[91] + src17[92] + src17[93] + src17[94] + src17[95] + src17[96] + src17[97] + src17[98] + src17[99] + src17[100] + src17[101] + src17[102] + src17[103] + src17[104] + src17[105] + src17[106] + src17[107] + src17[108] + src17[109] + src17[110] + src17[111] + src17[112] + src17[113] + src17[114] + src17[115] + src17[116] + src17[117] + src17[118] + src17[119] + src17[120] + src17[121] + src17[122] + src17[123] + src17[124] + src17[125] + src17[126] + src17[127])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31] + src18[32] + src18[33] + src18[34] + src18[35] + src18[36] + src18[37] + src18[38] + src18[39] + src18[40] + src18[41] + src18[42] + src18[43] + src18[44] + src18[45] + src18[46] + src18[47] + src18[48] + src18[49] + src18[50] + src18[51] + src18[52] + src18[53] + src18[54] + src18[55] + src18[56] + src18[57] + src18[58] + src18[59] + src18[60] + src18[61] + src18[62] + src18[63] + src18[64] + src18[65] + src18[66] + src18[67] + src18[68] + src18[69] + src18[70] + src18[71] + src18[72] + src18[73] + src18[74] + src18[75] + src18[76] + src18[77] + src18[78] + src18[79] + src18[80] + src18[81] + src18[82] + src18[83] + src18[84] + src18[85] + src18[86] + src18[87] + src18[88] + src18[89] + src18[90] + src18[91] + src18[92] + src18[93] + src18[94] + src18[95] + src18[96] + src18[97] + src18[98] + src18[99] + src18[100] + src18[101] + src18[102] + src18[103] + src18[104] + src18[105] + src18[106] + src18[107] + src18[108] + src18[109] + src18[110] + src18[111] + src18[112] + src18[113] + src18[114] + src18[115] + src18[116] + src18[117] + src18[118] + src18[119] + src18[120] + src18[121] + src18[122] + src18[123] + src18[124] + src18[125] + src18[126] + src18[127])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31] + src19[32] + src19[33] + src19[34] + src19[35] + src19[36] + src19[37] + src19[38] + src19[39] + src19[40] + src19[41] + src19[42] + src19[43] + src19[44] + src19[45] + src19[46] + src19[47] + src19[48] + src19[49] + src19[50] + src19[51] + src19[52] + src19[53] + src19[54] + src19[55] + src19[56] + src19[57] + src19[58] + src19[59] + src19[60] + src19[61] + src19[62] + src19[63] + src19[64] + src19[65] + src19[66] + src19[67] + src19[68] + src19[69] + src19[70] + src19[71] + src19[72] + src19[73] + src19[74] + src19[75] + src19[76] + src19[77] + src19[78] + src19[79] + src19[80] + src19[81] + src19[82] + src19[83] + src19[84] + src19[85] + src19[86] + src19[87] + src19[88] + src19[89] + src19[90] + src19[91] + src19[92] + src19[93] + src19[94] + src19[95] + src19[96] + src19[97] + src19[98] + src19[99] + src19[100] + src19[101] + src19[102] + src19[103] + src19[104] + src19[105] + src19[106] + src19[107] + src19[108] + src19[109] + src19[110] + src19[111] + src19[112] + src19[113] + src19[114] + src19[115] + src19[116] + src19[117] + src19[118] + src19[119] + src19[120] + src19[121] + src19[122] + src19[123] + src19[124] + src19[125] + src19[126] + src19[127])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31] + src20[32] + src20[33] + src20[34] + src20[35] + src20[36] + src20[37] + src20[38] + src20[39] + src20[40] + src20[41] + src20[42] + src20[43] + src20[44] + src20[45] + src20[46] + src20[47] + src20[48] + src20[49] + src20[50] + src20[51] + src20[52] + src20[53] + src20[54] + src20[55] + src20[56] + src20[57] + src20[58] + src20[59] + src20[60] + src20[61] + src20[62] + src20[63] + src20[64] + src20[65] + src20[66] + src20[67] + src20[68] + src20[69] + src20[70] + src20[71] + src20[72] + src20[73] + src20[74] + src20[75] + src20[76] + src20[77] + src20[78] + src20[79] + src20[80] + src20[81] + src20[82] + src20[83] + src20[84] + src20[85] + src20[86] + src20[87] + src20[88] + src20[89] + src20[90] + src20[91] + src20[92] + src20[93] + src20[94] + src20[95] + src20[96] + src20[97] + src20[98] + src20[99] + src20[100] + src20[101] + src20[102] + src20[103] + src20[104] + src20[105] + src20[106] + src20[107] + src20[108] + src20[109] + src20[110] + src20[111] + src20[112] + src20[113] + src20[114] + src20[115] + src20[116] + src20[117] + src20[118] + src20[119] + src20[120] + src20[121] + src20[122] + src20[123] + src20[124] + src20[125] + src20[126] + src20[127])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31] + src21[32] + src21[33] + src21[34] + src21[35] + src21[36] + src21[37] + src21[38] + src21[39] + src21[40] + src21[41] + src21[42] + src21[43] + src21[44] + src21[45] + src21[46] + src21[47] + src21[48] + src21[49] + src21[50] + src21[51] + src21[52] + src21[53] + src21[54] + src21[55] + src21[56] + src21[57] + src21[58] + src21[59] + src21[60] + src21[61] + src21[62] + src21[63] + src21[64] + src21[65] + src21[66] + src21[67] + src21[68] + src21[69] + src21[70] + src21[71] + src21[72] + src21[73] + src21[74] + src21[75] + src21[76] + src21[77] + src21[78] + src21[79] + src21[80] + src21[81] + src21[82] + src21[83] + src21[84] + src21[85] + src21[86] + src21[87] + src21[88] + src21[89] + src21[90] + src21[91] + src21[92] + src21[93] + src21[94] + src21[95] + src21[96] + src21[97] + src21[98] + src21[99] + src21[100] + src21[101] + src21[102] + src21[103] + src21[104] + src21[105] + src21[106] + src21[107] + src21[108] + src21[109] + src21[110] + src21[111] + src21[112] + src21[113] + src21[114] + src21[115] + src21[116] + src21[117] + src21[118] + src21[119] + src21[120] + src21[121] + src21[122] + src21[123] + src21[124] + src21[125] + src21[126] + src21[127])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31] + src22[32] + src22[33] + src22[34] + src22[35] + src22[36] + src22[37] + src22[38] + src22[39] + src22[40] + src22[41] + src22[42] + src22[43] + src22[44] + src22[45] + src22[46] + src22[47] + src22[48] + src22[49] + src22[50] + src22[51] + src22[52] + src22[53] + src22[54] + src22[55] + src22[56] + src22[57] + src22[58] + src22[59] + src22[60] + src22[61] + src22[62] + src22[63] + src22[64] + src22[65] + src22[66] + src22[67] + src22[68] + src22[69] + src22[70] + src22[71] + src22[72] + src22[73] + src22[74] + src22[75] + src22[76] + src22[77] + src22[78] + src22[79] + src22[80] + src22[81] + src22[82] + src22[83] + src22[84] + src22[85] + src22[86] + src22[87] + src22[88] + src22[89] + src22[90] + src22[91] + src22[92] + src22[93] + src22[94] + src22[95] + src22[96] + src22[97] + src22[98] + src22[99] + src22[100] + src22[101] + src22[102] + src22[103] + src22[104] + src22[105] + src22[106] + src22[107] + src22[108] + src22[109] + src22[110] + src22[111] + src22[112] + src22[113] + src22[114] + src22[115] + src22[116] + src22[117] + src22[118] + src22[119] + src22[120] + src22[121] + src22[122] + src22[123] + src22[124] + src22[125] + src22[126] + src22[127])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31] + src23[32] + src23[33] + src23[34] + src23[35] + src23[36] + src23[37] + src23[38] + src23[39] + src23[40] + src23[41] + src23[42] + src23[43] + src23[44] + src23[45] + src23[46] + src23[47] + src23[48] + src23[49] + src23[50] + src23[51] + src23[52] + src23[53] + src23[54] + src23[55] + src23[56] + src23[57] + src23[58] + src23[59] + src23[60] + src23[61] + src23[62] + src23[63] + src23[64] + src23[65] + src23[66] + src23[67] + src23[68] + src23[69] + src23[70] + src23[71] + src23[72] + src23[73] + src23[74] + src23[75] + src23[76] + src23[77] + src23[78] + src23[79] + src23[80] + src23[81] + src23[82] + src23[83] + src23[84] + src23[85] + src23[86] + src23[87] + src23[88] + src23[89] + src23[90] + src23[91] + src23[92] + src23[93] + src23[94] + src23[95] + src23[96] + src23[97] + src23[98] + src23[99] + src23[100] + src23[101] + src23[102] + src23[103] + src23[104] + src23[105] + src23[106] + src23[107] + src23[108] + src23[109] + src23[110] + src23[111] + src23[112] + src23[113] + src23[114] + src23[115] + src23[116] + src23[117] + src23[118] + src23[119] + src23[120] + src23[121] + src23[122] + src23[123] + src23[124] + src23[125] + src23[126] + src23[127])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31] + src24[32] + src24[33] + src24[34] + src24[35] + src24[36] + src24[37] + src24[38] + src24[39] + src24[40] + src24[41] + src24[42] + src24[43] + src24[44] + src24[45] + src24[46] + src24[47] + src24[48] + src24[49] + src24[50] + src24[51] + src24[52] + src24[53] + src24[54] + src24[55] + src24[56] + src24[57] + src24[58] + src24[59] + src24[60] + src24[61] + src24[62] + src24[63] + src24[64] + src24[65] + src24[66] + src24[67] + src24[68] + src24[69] + src24[70] + src24[71] + src24[72] + src24[73] + src24[74] + src24[75] + src24[76] + src24[77] + src24[78] + src24[79] + src24[80] + src24[81] + src24[82] + src24[83] + src24[84] + src24[85] + src24[86] + src24[87] + src24[88] + src24[89] + src24[90] + src24[91] + src24[92] + src24[93] + src24[94] + src24[95] + src24[96] + src24[97] + src24[98] + src24[99] + src24[100] + src24[101] + src24[102] + src24[103] + src24[104] + src24[105] + src24[106] + src24[107] + src24[108] + src24[109] + src24[110] + src24[111] + src24[112] + src24[113] + src24[114] + src24[115] + src24[116] + src24[117] + src24[118] + src24[119] + src24[120] + src24[121] + src24[122] + src24[123] + src24[124] + src24[125] + src24[126] + src24[127])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31] + src25[32] + src25[33] + src25[34] + src25[35] + src25[36] + src25[37] + src25[38] + src25[39] + src25[40] + src25[41] + src25[42] + src25[43] + src25[44] + src25[45] + src25[46] + src25[47] + src25[48] + src25[49] + src25[50] + src25[51] + src25[52] + src25[53] + src25[54] + src25[55] + src25[56] + src25[57] + src25[58] + src25[59] + src25[60] + src25[61] + src25[62] + src25[63] + src25[64] + src25[65] + src25[66] + src25[67] + src25[68] + src25[69] + src25[70] + src25[71] + src25[72] + src25[73] + src25[74] + src25[75] + src25[76] + src25[77] + src25[78] + src25[79] + src25[80] + src25[81] + src25[82] + src25[83] + src25[84] + src25[85] + src25[86] + src25[87] + src25[88] + src25[89] + src25[90] + src25[91] + src25[92] + src25[93] + src25[94] + src25[95] + src25[96] + src25[97] + src25[98] + src25[99] + src25[100] + src25[101] + src25[102] + src25[103] + src25[104] + src25[105] + src25[106] + src25[107] + src25[108] + src25[109] + src25[110] + src25[111] + src25[112] + src25[113] + src25[114] + src25[115] + src25[116] + src25[117] + src25[118] + src25[119] + src25[120] + src25[121] + src25[122] + src25[123] + src25[124] + src25[125] + src25[126] + src25[127])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31] + src26[32] + src26[33] + src26[34] + src26[35] + src26[36] + src26[37] + src26[38] + src26[39] + src26[40] + src26[41] + src26[42] + src26[43] + src26[44] + src26[45] + src26[46] + src26[47] + src26[48] + src26[49] + src26[50] + src26[51] + src26[52] + src26[53] + src26[54] + src26[55] + src26[56] + src26[57] + src26[58] + src26[59] + src26[60] + src26[61] + src26[62] + src26[63] + src26[64] + src26[65] + src26[66] + src26[67] + src26[68] + src26[69] + src26[70] + src26[71] + src26[72] + src26[73] + src26[74] + src26[75] + src26[76] + src26[77] + src26[78] + src26[79] + src26[80] + src26[81] + src26[82] + src26[83] + src26[84] + src26[85] + src26[86] + src26[87] + src26[88] + src26[89] + src26[90] + src26[91] + src26[92] + src26[93] + src26[94] + src26[95] + src26[96] + src26[97] + src26[98] + src26[99] + src26[100] + src26[101] + src26[102] + src26[103] + src26[104] + src26[105] + src26[106] + src26[107] + src26[108] + src26[109] + src26[110] + src26[111] + src26[112] + src26[113] + src26[114] + src26[115] + src26[116] + src26[117] + src26[118] + src26[119] + src26[120] + src26[121] + src26[122] + src26[123] + src26[124] + src26[125] + src26[126] + src26[127])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31] + src27[32] + src27[33] + src27[34] + src27[35] + src27[36] + src27[37] + src27[38] + src27[39] + src27[40] + src27[41] + src27[42] + src27[43] + src27[44] + src27[45] + src27[46] + src27[47] + src27[48] + src27[49] + src27[50] + src27[51] + src27[52] + src27[53] + src27[54] + src27[55] + src27[56] + src27[57] + src27[58] + src27[59] + src27[60] + src27[61] + src27[62] + src27[63] + src27[64] + src27[65] + src27[66] + src27[67] + src27[68] + src27[69] + src27[70] + src27[71] + src27[72] + src27[73] + src27[74] + src27[75] + src27[76] + src27[77] + src27[78] + src27[79] + src27[80] + src27[81] + src27[82] + src27[83] + src27[84] + src27[85] + src27[86] + src27[87] + src27[88] + src27[89] + src27[90] + src27[91] + src27[92] + src27[93] + src27[94] + src27[95] + src27[96] + src27[97] + src27[98] + src27[99] + src27[100] + src27[101] + src27[102] + src27[103] + src27[104] + src27[105] + src27[106] + src27[107] + src27[108] + src27[109] + src27[110] + src27[111] + src27[112] + src27[113] + src27[114] + src27[115] + src27[116] + src27[117] + src27[118] + src27[119] + src27[120] + src27[121] + src27[122] + src27[123] + src27[124] + src27[125] + src27[126] + src27[127])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31] + src28[32] + src28[33] + src28[34] + src28[35] + src28[36] + src28[37] + src28[38] + src28[39] + src28[40] + src28[41] + src28[42] + src28[43] + src28[44] + src28[45] + src28[46] + src28[47] + src28[48] + src28[49] + src28[50] + src28[51] + src28[52] + src28[53] + src28[54] + src28[55] + src28[56] + src28[57] + src28[58] + src28[59] + src28[60] + src28[61] + src28[62] + src28[63] + src28[64] + src28[65] + src28[66] + src28[67] + src28[68] + src28[69] + src28[70] + src28[71] + src28[72] + src28[73] + src28[74] + src28[75] + src28[76] + src28[77] + src28[78] + src28[79] + src28[80] + src28[81] + src28[82] + src28[83] + src28[84] + src28[85] + src28[86] + src28[87] + src28[88] + src28[89] + src28[90] + src28[91] + src28[92] + src28[93] + src28[94] + src28[95] + src28[96] + src28[97] + src28[98] + src28[99] + src28[100] + src28[101] + src28[102] + src28[103] + src28[104] + src28[105] + src28[106] + src28[107] + src28[108] + src28[109] + src28[110] + src28[111] + src28[112] + src28[113] + src28[114] + src28[115] + src28[116] + src28[117] + src28[118] + src28[119] + src28[120] + src28[121] + src28[122] + src28[123] + src28[124] + src28[125] + src28[126] + src28[127])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31] + src29[32] + src29[33] + src29[34] + src29[35] + src29[36] + src29[37] + src29[38] + src29[39] + src29[40] + src29[41] + src29[42] + src29[43] + src29[44] + src29[45] + src29[46] + src29[47] + src29[48] + src29[49] + src29[50] + src29[51] + src29[52] + src29[53] + src29[54] + src29[55] + src29[56] + src29[57] + src29[58] + src29[59] + src29[60] + src29[61] + src29[62] + src29[63] + src29[64] + src29[65] + src29[66] + src29[67] + src29[68] + src29[69] + src29[70] + src29[71] + src29[72] + src29[73] + src29[74] + src29[75] + src29[76] + src29[77] + src29[78] + src29[79] + src29[80] + src29[81] + src29[82] + src29[83] + src29[84] + src29[85] + src29[86] + src29[87] + src29[88] + src29[89] + src29[90] + src29[91] + src29[92] + src29[93] + src29[94] + src29[95] + src29[96] + src29[97] + src29[98] + src29[99] + src29[100] + src29[101] + src29[102] + src29[103] + src29[104] + src29[105] + src29[106] + src29[107] + src29[108] + src29[109] + src29[110] + src29[111] + src29[112] + src29[113] + src29[114] + src29[115] + src29[116] + src29[117] + src29[118] + src29[119] + src29[120] + src29[121] + src29[122] + src29[123] + src29[124] + src29[125] + src29[126] + src29[127])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31] + src30[32] + src30[33] + src30[34] + src30[35] + src30[36] + src30[37] + src30[38] + src30[39] + src30[40] + src30[41] + src30[42] + src30[43] + src30[44] + src30[45] + src30[46] + src30[47] + src30[48] + src30[49] + src30[50] + src30[51] + src30[52] + src30[53] + src30[54] + src30[55] + src30[56] + src30[57] + src30[58] + src30[59] + src30[60] + src30[61] + src30[62] + src30[63] + src30[64] + src30[65] + src30[66] + src30[67] + src30[68] + src30[69] + src30[70] + src30[71] + src30[72] + src30[73] + src30[74] + src30[75] + src30[76] + src30[77] + src30[78] + src30[79] + src30[80] + src30[81] + src30[82] + src30[83] + src30[84] + src30[85] + src30[86] + src30[87] + src30[88] + src30[89] + src30[90] + src30[91] + src30[92] + src30[93] + src30[94] + src30[95] + src30[96] + src30[97] + src30[98] + src30[99] + src30[100] + src30[101] + src30[102] + src30[103] + src30[104] + src30[105] + src30[106] + src30[107] + src30[108] + src30[109] + src30[110] + src30[111] + src30[112] + src30[113] + src30[114] + src30[115] + src30[116] + src30[117] + src30[118] + src30[119] + src30[120] + src30[121] + src30[122] + src30[123] + src30[124] + src30[125] + src30[126] + src30[127])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31] + src31[32] + src31[33] + src31[34] + src31[35] + src31[36] + src31[37] + src31[38] + src31[39] + src31[40] + src31[41] + src31[42] + src31[43] + src31[44] + src31[45] + src31[46] + src31[47] + src31[48] + src31[49] + src31[50] + src31[51] + src31[52] + src31[53] + src31[54] + src31[55] + src31[56] + src31[57] + src31[58] + src31[59] + src31[60] + src31[61] + src31[62] + src31[63] + src31[64] + src31[65] + src31[66] + src31[67] + src31[68] + src31[69] + src31[70] + src31[71] + src31[72] + src31[73] + src31[74] + src31[75] + src31[76] + src31[77] + src31[78] + src31[79] + src31[80] + src31[81] + src31[82] + src31[83] + src31[84] + src31[85] + src31[86] + src31[87] + src31[88] + src31[89] + src31[90] + src31[91] + src31[92] + src31[93] + src31[94] + src31[95] + src31[96] + src31[97] + src31[98] + src31[99] + src31[100] + src31[101] + src31[102] + src31[103] + src31[104] + src31[105] + src31[106] + src31[107] + src31[108] + src31[109] + src31[110] + src31[111] + src31[112] + src31[113] + src31[114] + src31[115] + src31[116] + src31[117] + src31[118] + src31[119] + src31[120] + src31[121] + src31[122] + src31[123] + src31[124] + src31[125] + src31[126] + src31[127])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31] + src32[32] + src32[33] + src32[34] + src32[35] + src32[36] + src32[37] + src32[38] + src32[39] + src32[40] + src32[41] + src32[42] + src32[43] + src32[44] + src32[45] + src32[46] + src32[47] + src32[48] + src32[49] + src32[50] + src32[51] + src32[52] + src32[53] + src32[54] + src32[55] + src32[56] + src32[57] + src32[58] + src32[59] + src32[60] + src32[61] + src32[62] + src32[63] + src32[64] + src32[65] + src32[66] + src32[67] + src32[68] + src32[69] + src32[70] + src32[71] + src32[72] + src32[73] + src32[74] + src32[75] + src32[76] + src32[77] + src32[78] + src32[79] + src32[80] + src32[81] + src32[82] + src32[83] + src32[84] + src32[85] + src32[86] + src32[87] + src32[88] + src32[89] + src32[90] + src32[91] + src32[92] + src32[93] + src32[94] + src32[95] + src32[96] + src32[97] + src32[98] + src32[99] + src32[100] + src32[101] + src32[102] + src32[103] + src32[104] + src32[105] + src32[106] + src32[107] + src32[108] + src32[109] + src32[110] + src32[111] + src32[112] + src32[113] + src32[114] + src32[115] + src32[116] + src32[117] + src32[118] + src32[119] + src32[120] + src32[121] + src32[122] + src32[123] + src32[124] + src32[125] + src32[126] + src32[127])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31] + src33[32] + src33[33] + src33[34] + src33[35] + src33[36] + src33[37] + src33[38] + src33[39] + src33[40] + src33[41] + src33[42] + src33[43] + src33[44] + src33[45] + src33[46] + src33[47] + src33[48] + src33[49] + src33[50] + src33[51] + src33[52] + src33[53] + src33[54] + src33[55] + src33[56] + src33[57] + src33[58] + src33[59] + src33[60] + src33[61] + src33[62] + src33[63] + src33[64] + src33[65] + src33[66] + src33[67] + src33[68] + src33[69] + src33[70] + src33[71] + src33[72] + src33[73] + src33[74] + src33[75] + src33[76] + src33[77] + src33[78] + src33[79] + src33[80] + src33[81] + src33[82] + src33[83] + src33[84] + src33[85] + src33[86] + src33[87] + src33[88] + src33[89] + src33[90] + src33[91] + src33[92] + src33[93] + src33[94] + src33[95] + src33[96] + src33[97] + src33[98] + src33[99] + src33[100] + src33[101] + src33[102] + src33[103] + src33[104] + src33[105] + src33[106] + src33[107] + src33[108] + src33[109] + src33[110] + src33[111] + src33[112] + src33[113] + src33[114] + src33[115] + src33[116] + src33[117] + src33[118] + src33[119] + src33[120] + src33[121] + src33[122] + src33[123] + src33[124] + src33[125] + src33[126] + src33[127])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31] + src34[32] + src34[33] + src34[34] + src34[35] + src34[36] + src34[37] + src34[38] + src34[39] + src34[40] + src34[41] + src34[42] + src34[43] + src34[44] + src34[45] + src34[46] + src34[47] + src34[48] + src34[49] + src34[50] + src34[51] + src34[52] + src34[53] + src34[54] + src34[55] + src34[56] + src34[57] + src34[58] + src34[59] + src34[60] + src34[61] + src34[62] + src34[63] + src34[64] + src34[65] + src34[66] + src34[67] + src34[68] + src34[69] + src34[70] + src34[71] + src34[72] + src34[73] + src34[74] + src34[75] + src34[76] + src34[77] + src34[78] + src34[79] + src34[80] + src34[81] + src34[82] + src34[83] + src34[84] + src34[85] + src34[86] + src34[87] + src34[88] + src34[89] + src34[90] + src34[91] + src34[92] + src34[93] + src34[94] + src34[95] + src34[96] + src34[97] + src34[98] + src34[99] + src34[100] + src34[101] + src34[102] + src34[103] + src34[104] + src34[105] + src34[106] + src34[107] + src34[108] + src34[109] + src34[110] + src34[111] + src34[112] + src34[113] + src34[114] + src34[115] + src34[116] + src34[117] + src34[118] + src34[119] + src34[120] + src34[121] + src34[122] + src34[123] + src34[124] + src34[125] + src34[126] + src34[127])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31] + src35[32] + src35[33] + src35[34] + src35[35] + src35[36] + src35[37] + src35[38] + src35[39] + src35[40] + src35[41] + src35[42] + src35[43] + src35[44] + src35[45] + src35[46] + src35[47] + src35[48] + src35[49] + src35[50] + src35[51] + src35[52] + src35[53] + src35[54] + src35[55] + src35[56] + src35[57] + src35[58] + src35[59] + src35[60] + src35[61] + src35[62] + src35[63] + src35[64] + src35[65] + src35[66] + src35[67] + src35[68] + src35[69] + src35[70] + src35[71] + src35[72] + src35[73] + src35[74] + src35[75] + src35[76] + src35[77] + src35[78] + src35[79] + src35[80] + src35[81] + src35[82] + src35[83] + src35[84] + src35[85] + src35[86] + src35[87] + src35[88] + src35[89] + src35[90] + src35[91] + src35[92] + src35[93] + src35[94] + src35[95] + src35[96] + src35[97] + src35[98] + src35[99] + src35[100] + src35[101] + src35[102] + src35[103] + src35[104] + src35[105] + src35[106] + src35[107] + src35[108] + src35[109] + src35[110] + src35[111] + src35[112] + src35[113] + src35[114] + src35[115] + src35[116] + src35[117] + src35[118] + src35[119] + src35[120] + src35[121] + src35[122] + src35[123] + src35[124] + src35[125] + src35[126] + src35[127])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31] + src36[32] + src36[33] + src36[34] + src36[35] + src36[36] + src36[37] + src36[38] + src36[39] + src36[40] + src36[41] + src36[42] + src36[43] + src36[44] + src36[45] + src36[46] + src36[47] + src36[48] + src36[49] + src36[50] + src36[51] + src36[52] + src36[53] + src36[54] + src36[55] + src36[56] + src36[57] + src36[58] + src36[59] + src36[60] + src36[61] + src36[62] + src36[63] + src36[64] + src36[65] + src36[66] + src36[67] + src36[68] + src36[69] + src36[70] + src36[71] + src36[72] + src36[73] + src36[74] + src36[75] + src36[76] + src36[77] + src36[78] + src36[79] + src36[80] + src36[81] + src36[82] + src36[83] + src36[84] + src36[85] + src36[86] + src36[87] + src36[88] + src36[89] + src36[90] + src36[91] + src36[92] + src36[93] + src36[94] + src36[95] + src36[96] + src36[97] + src36[98] + src36[99] + src36[100] + src36[101] + src36[102] + src36[103] + src36[104] + src36[105] + src36[106] + src36[107] + src36[108] + src36[109] + src36[110] + src36[111] + src36[112] + src36[113] + src36[114] + src36[115] + src36[116] + src36[117] + src36[118] + src36[119] + src36[120] + src36[121] + src36[122] + src36[123] + src36[124] + src36[125] + src36[126] + src36[127])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31] + src37[32] + src37[33] + src37[34] + src37[35] + src37[36] + src37[37] + src37[38] + src37[39] + src37[40] + src37[41] + src37[42] + src37[43] + src37[44] + src37[45] + src37[46] + src37[47] + src37[48] + src37[49] + src37[50] + src37[51] + src37[52] + src37[53] + src37[54] + src37[55] + src37[56] + src37[57] + src37[58] + src37[59] + src37[60] + src37[61] + src37[62] + src37[63] + src37[64] + src37[65] + src37[66] + src37[67] + src37[68] + src37[69] + src37[70] + src37[71] + src37[72] + src37[73] + src37[74] + src37[75] + src37[76] + src37[77] + src37[78] + src37[79] + src37[80] + src37[81] + src37[82] + src37[83] + src37[84] + src37[85] + src37[86] + src37[87] + src37[88] + src37[89] + src37[90] + src37[91] + src37[92] + src37[93] + src37[94] + src37[95] + src37[96] + src37[97] + src37[98] + src37[99] + src37[100] + src37[101] + src37[102] + src37[103] + src37[104] + src37[105] + src37[106] + src37[107] + src37[108] + src37[109] + src37[110] + src37[111] + src37[112] + src37[113] + src37[114] + src37[115] + src37[116] + src37[117] + src37[118] + src37[119] + src37[120] + src37[121] + src37[122] + src37[123] + src37[124] + src37[125] + src37[126] + src37[127])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31] + src38[32] + src38[33] + src38[34] + src38[35] + src38[36] + src38[37] + src38[38] + src38[39] + src38[40] + src38[41] + src38[42] + src38[43] + src38[44] + src38[45] + src38[46] + src38[47] + src38[48] + src38[49] + src38[50] + src38[51] + src38[52] + src38[53] + src38[54] + src38[55] + src38[56] + src38[57] + src38[58] + src38[59] + src38[60] + src38[61] + src38[62] + src38[63] + src38[64] + src38[65] + src38[66] + src38[67] + src38[68] + src38[69] + src38[70] + src38[71] + src38[72] + src38[73] + src38[74] + src38[75] + src38[76] + src38[77] + src38[78] + src38[79] + src38[80] + src38[81] + src38[82] + src38[83] + src38[84] + src38[85] + src38[86] + src38[87] + src38[88] + src38[89] + src38[90] + src38[91] + src38[92] + src38[93] + src38[94] + src38[95] + src38[96] + src38[97] + src38[98] + src38[99] + src38[100] + src38[101] + src38[102] + src38[103] + src38[104] + src38[105] + src38[106] + src38[107] + src38[108] + src38[109] + src38[110] + src38[111] + src38[112] + src38[113] + src38[114] + src38[115] + src38[116] + src38[117] + src38[118] + src38[119] + src38[120] + src38[121] + src38[122] + src38[123] + src38[124] + src38[125] + src38[126] + src38[127])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31] + src39[32] + src39[33] + src39[34] + src39[35] + src39[36] + src39[37] + src39[38] + src39[39] + src39[40] + src39[41] + src39[42] + src39[43] + src39[44] + src39[45] + src39[46] + src39[47] + src39[48] + src39[49] + src39[50] + src39[51] + src39[52] + src39[53] + src39[54] + src39[55] + src39[56] + src39[57] + src39[58] + src39[59] + src39[60] + src39[61] + src39[62] + src39[63] + src39[64] + src39[65] + src39[66] + src39[67] + src39[68] + src39[69] + src39[70] + src39[71] + src39[72] + src39[73] + src39[74] + src39[75] + src39[76] + src39[77] + src39[78] + src39[79] + src39[80] + src39[81] + src39[82] + src39[83] + src39[84] + src39[85] + src39[86] + src39[87] + src39[88] + src39[89] + src39[90] + src39[91] + src39[92] + src39[93] + src39[94] + src39[95] + src39[96] + src39[97] + src39[98] + src39[99] + src39[100] + src39[101] + src39[102] + src39[103] + src39[104] + src39[105] + src39[106] + src39[107] + src39[108] + src39[109] + src39[110] + src39[111] + src39[112] + src39[113] + src39[114] + src39[115] + src39[116] + src39[117] + src39[118] + src39[119] + src39[120] + src39[121] + src39[122] + src39[123] + src39[124] + src39[125] + src39[126] + src39[127])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31] + src40[32] + src40[33] + src40[34] + src40[35] + src40[36] + src40[37] + src40[38] + src40[39] + src40[40] + src40[41] + src40[42] + src40[43] + src40[44] + src40[45] + src40[46] + src40[47] + src40[48] + src40[49] + src40[50] + src40[51] + src40[52] + src40[53] + src40[54] + src40[55] + src40[56] + src40[57] + src40[58] + src40[59] + src40[60] + src40[61] + src40[62] + src40[63] + src40[64] + src40[65] + src40[66] + src40[67] + src40[68] + src40[69] + src40[70] + src40[71] + src40[72] + src40[73] + src40[74] + src40[75] + src40[76] + src40[77] + src40[78] + src40[79] + src40[80] + src40[81] + src40[82] + src40[83] + src40[84] + src40[85] + src40[86] + src40[87] + src40[88] + src40[89] + src40[90] + src40[91] + src40[92] + src40[93] + src40[94] + src40[95] + src40[96] + src40[97] + src40[98] + src40[99] + src40[100] + src40[101] + src40[102] + src40[103] + src40[104] + src40[105] + src40[106] + src40[107] + src40[108] + src40[109] + src40[110] + src40[111] + src40[112] + src40[113] + src40[114] + src40[115] + src40[116] + src40[117] + src40[118] + src40[119] + src40[120] + src40[121] + src40[122] + src40[123] + src40[124] + src40[125] + src40[126] + src40[127])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31] + src41[32] + src41[33] + src41[34] + src41[35] + src41[36] + src41[37] + src41[38] + src41[39] + src41[40] + src41[41] + src41[42] + src41[43] + src41[44] + src41[45] + src41[46] + src41[47] + src41[48] + src41[49] + src41[50] + src41[51] + src41[52] + src41[53] + src41[54] + src41[55] + src41[56] + src41[57] + src41[58] + src41[59] + src41[60] + src41[61] + src41[62] + src41[63] + src41[64] + src41[65] + src41[66] + src41[67] + src41[68] + src41[69] + src41[70] + src41[71] + src41[72] + src41[73] + src41[74] + src41[75] + src41[76] + src41[77] + src41[78] + src41[79] + src41[80] + src41[81] + src41[82] + src41[83] + src41[84] + src41[85] + src41[86] + src41[87] + src41[88] + src41[89] + src41[90] + src41[91] + src41[92] + src41[93] + src41[94] + src41[95] + src41[96] + src41[97] + src41[98] + src41[99] + src41[100] + src41[101] + src41[102] + src41[103] + src41[104] + src41[105] + src41[106] + src41[107] + src41[108] + src41[109] + src41[110] + src41[111] + src41[112] + src41[113] + src41[114] + src41[115] + src41[116] + src41[117] + src41[118] + src41[119] + src41[120] + src41[121] + src41[122] + src41[123] + src41[124] + src41[125] + src41[126] + src41[127])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31] + src42[32] + src42[33] + src42[34] + src42[35] + src42[36] + src42[37] + src42[38] + src42[39] + src42[40] + src42[41] + src42[42] + src42[43] + src42[44] + src42[45] + src42[46] + src42[47] + src42[48] + src42[49] + src42[50] + src42[51] + src42[52] + src42[53] + src42[54] + src42[55] + src42[56] + src42[57] + src42[58] + src42[59] + src42[60] + src42[61] + src42[62] + src42[63] + src42[64] + src42[65] + src42[66] + src42[67] + src42[68] + src42[69] + src42[70] + src42[71] + src42[72] + src42[73] + src42[74] + src42[75] + src42[76] + src42[77] + src42[78] + src42[79] + src42[80] + src42[81] + src42[82] + src42[83] + src42[84] + src42[85] + src42[86] + src42[87] + src42[88] + src42[89] + src42[90] + src42[91] + src42[92] + src42[93] + src42[94] + src42[95] + src42[96] + src42[97] + src42[98] + src42[99] + src42[100] + src42[101] + src42[102] + src42[103] + src42[104] + src42[105] + src42[106] + src42[107] + src42[108] + src42[109] + src42[110] + src42[111] + src42[112] + src42[113] + src42[114] + src42[115] + src42[116] + src42[117] + src42[118] + src42[119] + src42[120] + src42[121] + src42[122] + src42[123] + src42[124] + src42[125] + src42[126] + src42[127])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31] + src43[32] + src43[33] + src43[34] + src43[35] + src43[36] + src43[37] + src43[38] + src43[39] + src43[40] + src43[41] + src43[42] + src43[43] + src43[44] + src43[45] + src43[46] + src43[47] + src43[48] + src43[49] + src43[50] + src43[51] + src43[52] + src43[53] + src43[54] + src43[55] + src43[56] + src43[57] + src43[58] + src43[59] + src43[60] + src43[61] + src43[62] + src43[63] + src43[64] + src43[65] + src43[66] + src43[67] + src43[68] + src43[69] + src43[70] + src43[71] + src43[72] + src43[73] + src43[74] + src43[75] + src43[76] + src43[77] + src43[78] + src43[79] + src43[80] + src43[81] + src43[82] + src43[83] + src43[84] + src43[85] + src43[86] + src43[87] + src43[88] + src43[89] + src43[90] + src43[91] + src43[92] + src43[93] + src43[94] + src43[95] + src43[96] + src43[97] + src43[98] + src43[99] + src43[100] + src43[101] + src43[102] + src43[103] + src43[104] + src43[105] + src43[106] + src43[107] + src43[108] + src43[109] + src43[110] + src43[111] + src43[112] + src43[113] + src43[114] + src43[115] + src43[116] + src43[117] + src43[118] + src43[119] + src43[120] + src43[121] + src43[122] + src43[123] + src43[124] + src43[125] + src43[126] + src43[127])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31] + src44[32] + src44[33] + src44[34] + src44[35] + src44[36] + src44[37] + src44[38] + src44[39] + src44[40] + src44[41] + src44[42] + src44[43] + src44[44] + src44[45] + src44[46] + src44[47] + src44[48] + src44[49] + src44[50] + src44[51] + src44[52] + src44[53] + src44[54] + src44[55] + src44[56] + src44[57] + src44[58] + src44[59] + src44[60] + src44[61] + src44[62] + src44[63] + src44[64] + src44[65] + src44[66] + src44[67] + src44[68] + src44[69] + src44[70] + src44[71] + src44[72] + src44[73] + src44[74] + src44[75] + src44[76] + src44[77] + src44[78] + src44[79] + src44[80] + src44[81] + src44[82] + src44[83] + src44[84] + src44[85] + src44[86] + src44[87] + src44[88] + src44[89] + src44[90] + src44[91] + src44[92] + src44[93] + src44[94] + src44[95] + src44[96] + src44[97] + src44[98] + src44[99] + src44[100] + src44[101] + src44[102] + src44[103] + src44[104] + src44[105] + src44[106] + src44[107] + src44[108] + src44[109] + src44[110] + src44[111] + src44[112] + src44[113] + src44[114] + src44[115] + src44[116] + src44[117] + src44[118] + src44[119] + src44[120] + src44[121] + src44[122] + src44[123] + src44[124] + src44[125] + src44[126] + src44[127])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31] + src45[32] + src45[33] + src45[34] + src45[35] + src45[36] + src45[37] + src45[38] + src45[39] + src45[40] + src45[41] + src45[42] + src45[43] + src45[44] + src45[45] + src45[46] + src45[47] + src45[48] + src45[49] + src45[50] + src45[51] + src45[52] + src45[53] + src45[54] + src45[55] + src45[56] + src45[57] + src45[58] + src45[59] + src45[60] + src45[61] + src45[62] + src45[63] + src45[64] + src45[65] + src45[66] + src45[67] + src45[68] + src45[69] + src45[70] + src45[71] + src45[72] + src45[73] + src45[74] + src45[75] + src45[76] + src45[77] + src45[78] + src45[79] + src45[80] + src45[81] + src45[82] + src45[83] + src45[84] + src45[85] + src45[86] + src45[87] + src45[88] + src45[89] + src45[90] + src45[91] + src45[92] + src45[93] + src45[94] + src45[95] + src45[96] + src45[97] + src45[98] + src45[99] + src45[100] + src45[101] + src45[102] + src45[103] + src45[104] + src45[105] + src45[106] + src45[107] + src45[108] + src45[109] + src45[110] + src45[111] + src45[112] + src45[113] + src45[114] + src45[115] + src45[116] + src45[117] + src45[118] + src45[119] + src45[120] + src45[121] + src45[122] + src45[123] + src45[124] + src45[125] + src45[126] + src45[127])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31] + src46[32] + src46[33] + src46[34] + src46[35] + src46[36] + src46[37] + src46[38] + src46[39] + src46[40] + src46[41] + src46[42] + src46[43] + src46[44] + src46[45] + src46[46] + src46[47] + src46[48] + src46[49] + src46[50] + src46[51] + src46[52] + src46[53] + src46[54] + src46[55] + src46[56] + src46[57] + src46[58] + src46[59] + src46[60] + src46[61] + src46[62] + src46[63] + src46[64] + src46[65] + src46[66] + src46[67] + src46[68] + src46[69] + src46[70] + src46[71] + src46[72] + src46[73] + src46[74] + src46[75] + src46[76] + src46[77] + src46[78] + src46[79] + src46[80] + src46[81] + src46[82] + src46[83] + src46[84] + src46[85] + src46[86] + src46[87] + src46[88] + src46[89] + src46[90] + src46[91] + src46[92] + src46[93] + src46[94] + src46[95] + src46[96] + src46[97] + src46[98] + src46[99] + src46[100] + src46[101] + src46[102] + src46[103] + src46[104] + src46[105] + src46[106] + src46[107] + src46[108] + src46[109] + src46[110] + src46[111] + src46[112] + src46[113] + src46[114] + src46[115] + src46[116] + src46[117] + src46[118] + src46[119] + src46[120] + src46[121] + src46[122] + src46[123] + src46[124] + src46[125] + src46[126] + src46[127])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31] + src47[32] + src47[33] + src47[34] + src47[35] + src47[36] + src47[37] + src47[38] + src47[39] + src47[40] + src47[41] + src47[42] + src47[43] + src47[44] + src47[45] + src47[46] + src47[47] + src47[48] + src47[49] + src47[50] + src47[51] + src47[52] + src47[53] + src47[54] + src47[55] + src47[56] + src47[57] + src47[58] + src47[59] + src47[60] + src47[61] + src47[62] + src47[63] + src47[64] + src47[65] + src47[66] + src47[67] + src47[68] + src47[69] + src47[70] + src47[71] + src47[72] + src47[73] + src47[74] + src47[75] + src47[76] + src47[77] + src47[78] + src47[79] + src47[80] + src47[81] + src47[82] + src47[83] + src47[84] + src47[85] + src47[86] + src47[87] + src47[88] + src47[89] + src47[90] + src47[91] + src47[92] + src47[93] + src47[94] + src47[95] + src47[96] + src47[97] + src47[98] + src47[99] + src47[100] + src47[101] + src47[102] + src47[103] + src47[104] + src47[105] + src47[106] + src47[107] + src47[108] + src47[109] + src47[110] + src47[111] + src47[112] + src47[113] + src47[114] + src47[115] + src47[116] + src47[117] + src47[118] + src47[119] + src47[120] + src47[121] + src47[122] + src47[123] + src47[124] + src47[125] + src47[126] + src47[127])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31] + src48[32] + src48[33] + src48[34] + src48[35] + src48[36] + src48[37] + src48[38] + src48[39] + src48[40] + src48[41] + src48[42] + src48[43] + src48[44] + src48[45] + src48[46] + src48[47] + src48[48] + src48[49] + src48[50] + src48[51] + src48[52] + src48[53] + src48[54] + src48[55] + src48[56] + src48[57] + src48[58] + src48[59] + src48[60] + src48[61] + src48[62] + src48[63] + src48[64] + src48[65] + src48[66] + src48[67] + src48[68] + src48[69] + src48[70] + src48[71] + src48[72] + src48[73] + src48[74] + src48[75] + src48[76] + src48[77] + src48[78] + src48[79] + src48[80] + src48[81] + src48[82] + src48[83] + src48[84] + src48[85] + src48[86] + src48[87] + src48[88] + src48[89] + src48[90] + src48[91] + src48[92] + src48[93] + src48[94] + src48[95] + src48[96] + src48[97] + src48[98] + src48[99] + src48[100] + src48[101] + src48[102] + src48[103] + src48[104] + src48[105] + src48[106] + src48[107] + src48[108] + src48[109] + src48[110] + src48[111] + src48[112] + src48[113] + src48[114] + src48[115] + src48[116] + src48[117] + src48[118] + src48[119] + src48[120] + src48[121] + src48[122] + src48[123] + src48[124] + src48[125] + src48[126] + src48[127])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31] + src49[32] + src49[33] + src49[34] + src49[35] + src49[36] + src49[37] + src49[38] + src49[39] + src49[40] + src49[41] + src49[42] + src49[43] + src49[44] + src49[45] + src49[46] + src49[47] + src49[48] + src49[49] + src49[50] + src49[51] + src49[52] + src49[53] + src49[54] + src49[55] + src49[56] + src49[57] + src49[58] + src49[59] + src49[60] + src49[61] + src49[62] + src49[63] + src49[64] + src49[65] + src49[66] + src49[67] + src49[68] + src49[69] + src49[70] + src49[71] + src49[72] + src49[73] + src49[74] + src49[75] + src49[76] + src49[77] + src49[78] + src49[79] + src49[80] + src49[81] + src49[82] + src49[83] + src49[84] + src49[85] + src49[86] + src49[87] + src49[88] + src49[89] + src49[90] + src49[91] + src49[92] + src49[93] + src49[94] + src49[95] + src49[96] + src49[97] + src49[98] + src49[99] + src49[100] + src49[101] + src49[102] + src49[103] + src49[104] + src49[105] + src49[106] + src49[107] + src49[108] + src49[109] + src49[110] + src49[111] + src49[112] + src49[113] + src49[114] + src49[115] + src49[116] + src49[117] + src49[118] + src49[119] + src49[120] + src49[121] + src49[122] + src49[123] + src49[124] + src49[125] + src49[126] + src49[127])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31] + src50[32] + src50[33] + src50[34] + src50[35] + src50[36] + src50[37] + src50[38] + src50[39] + src50[40] + src50[41] + src50[42] + src50[43] + src50[44] + src50[45] + src50[46] + src50[47] + src50[48] + src50[49] + src50[50] + src50[51] + src50[52] + src50[53] + src50[54] + src50[55] + src50[56] + src50[57] + src50[58] + src50[59] + src50[60] + src50[61] + src50[62] + src50[63] + src50[64] + src50[65] + src50[66] + src50[67] + src50[68] + src50[69] + src50[70] + src50[71] + src50[72] + src50[73] + src50[74] + src50[75] + src50[76] + src50[77] + src50[78] + src50[79] + src50[80] + src50[81] + src50[82] + src50[83] + src50[84] + src50[85] + src50[86] + src50[87] + src50[88] + src50[89] + src50[90] + src50[91] + src50[92] + src50[93] + src50[94] + src50[95] + src50[96] + src50[97] + src50[98] + src50[99] + src50[100] + src50[101] + src50[102] + src50[103] + src50[104] + src50[105] + src50[106] + src50[107] + src50[108] + src50[109] + src50[110] + src50[111] + src50[112] + src50[113] + src50[114] + src50[115] + src50[116] + src50[117] + src50[118] + src50[119] + src50[120] + src50[121] + src50[122] + src50[123] + src50[124] + src50[125] + src50[126] + src50[127])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31] + src51[32] + src51[33] + src51[34] + src51[35] + src51[36] + src51[37] + src51[38] + src51[39] + src51[40] + src51[41] + src51[42] + src51[43] + src51[44] + src51[45] + src51[46] + src51[47] + src51[48] + src51[49] + src51[50] + src51[51] + src51[52] + src51[53] + src51[54] + src51[55] + src51[56] + src51[57] + src51[58] + src51[59] + src51[60] + src51[61] + src51[62] + src51[63] + src51[64] + src51[65] + src51[66] + src51[67] + src51[68] + src51[69] + src51[70] + src51[71] + src51[72] + src51[73] + src51[74] + src51[75] + src51[76] + src51[77] + src51[78] + src51[79] + src51[80] + src51[81] + src51[82] + src51[83] + src51[84] + src51[85] + src51[86] + src51[87] + src51[88] + src51[89] + src51[90] + src51[91] + src51[92] + src51[93] + src51[94] + src51[95] + src51[96] + src51[97] + src51[98] + src51[99] + src51[100] + src51[101] + src51[102] + src51[103] + src51[104] + src51[105] + src51[106] + src51[107] + src51[108] + src51[109] + src51[110] + src51[111] + src51[112] + src51[113] + src51[114] + src51[115] + src51[116] + src51[117] + src51[118] + src51[119] + src51[120] + src51[121] + src51[122] + src51[123] + src51[124] + src51[125] + src51[126] + src51[127])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31] + src52[32] + src52[33] + src52[34] + src52[35] + src52[36] + src52[37] + src52[38] + src52[39] + src52[40] + src52[41] + src52[42] + src52[43] + src52[44] + src52[45] + src52[46] + src52[47] + src52[48] + src52[49] + src52[50] + src52[51] + src52[52] + src52[53] + src52[54] + src52[55] + src52[56] + src52[57] + src52[58] + src52[59] + src52[60] + src52[61] + src52[62] + src52[63] + src52[64] + src52[65] + src52[66] + src52[67] + src52[68] + src52[69] + src52[70] + src52[71] + src52[72] + src52[73] + src52[74] + src52[75] + src52[76] + src52[77] + src52[78] + src52[79] + src52[80] + src52[81] + src52[82] + src52[83] + src52[84] + src52[85] + src52[86] + src52[87] + src52[88] + src52[89] + src52[90] + src52[91] + src52[92] + src52[93] + src52[94] + src52[95] + src52[96] + src52[97] + src52[98] + src52[99] + src52[100] + src52[101] + src52[102] + src52[103] + src52[104] + src52[105] + src52[106] + src52[107] + src52[108] + src52[109] + src52[110] + src52[111] + src52[112] + src52[113] + src52[114] + src52[115] + src52[116] + src52[117] + src52[118] + src52[119] + src52[120] + src52[121] + src52[122] + src52[123] + src52[124] + src52[125] + src52[126] + src52[127])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31] + src53[32] + src53[33] + src53[34] + src53[35] + src53[36] + src53[37] + src53[38] + src53[39] + src53[40] + src53[41] + src53[42] + src53[43] + src53[44] + src53[45] + src53[46] + src53[47] + src53[48] + src53[49] + src53[50] + src53[51] + src53[52] + src53[53] + src53[54] + src53[55] + src53[56] + src53[57] + src53[58] + src53[59] + src53[60] + src53[61] + src53[62] + src53[63] + src53[64] + src53[65] + src53[66] + src53[67] + src53[68] + src53[69] + src53[70] + src53[71] + src53[72] + src53[73] + src53[74] + src53[75] + src53[76] + src53[77] + src53[78] + src53[79] + src53[80] + src53[81] + src53[82] + src53[83] + src53[84] + src53[85] + src53[86] + src53[87] + src53[88] + src53[89] + src53[90] + src53[91] + src53[92] + src53[93] + src53[94] + src53[95] + src53[96] + src53[97] + src53[98] + src53[99] + src53[100] + src53[101] + src53[102] + src53[103] + src53[104] + src53[105] + src53[106] + src53[107] + src53[108] + src53[109] + src53[110] + src53[111] + src53[112] + src53[113] + src53[114] + src53[115] + src53[116] + src53[117] + src53[118] + src53[119] + src53[120] + src53[121] + src53[122] + src53[123] + src53[124] + src53[125] + src53[126] + src53[127])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31] + src54[32] + src54[33] + src54[34] + src54[35] + src54[36] + src54[37] + src54[38] + src54[39] + src54[40] + src54[41] + src54[42] + src54[43] + src54[44] + src54[45] + src54[46] + src54[47] + src54[48] + src54[49] + src54[50] + src54[51] + src54[52] + src54[53] + src54[54] + src54[55] + src54[56] + src54[57] + src54[58] + src54[59] + src54[60] + src54[61] + src54[62] + src54[63] + src54[64] + src54[65] + src54[66] + src54[67] + src54[68] + src54[69] + src54[70] + src54[71] + src54[72] + src54[73] + src54[74] + src54[75] + src54[76] + src54[77] + src54[78] + src54[79] + src54[80] + src54[81] + src54[82] + src54[83] + src54[84] + src54[85] + src54[86] + src54[87] + src54[88] + src54[89] + src54[90] + src54[91] + src54[92] + src54[93] + src54[94] + src54[95] + src54[96] + src54[97] + src54[98] + src54[99] + src54[100] + src54[101] + src54[102] + src54[103] + src54[104] + src54[105] + src54[106] + src54[107] + src54[108] + src54[109] + src54[110] + src54[111] + src54[112] + src54[113] + src54[114] + src54[115] + src54[116] + src54[117] + src54[118] + src54[119] + src54[120] + src54[121] + src54[122] + src54[123] + src54[124] + src54[125] + src54[126] + src54[127])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31] + src55[32] + src55[33] + src55[34] + src55[35] + src55[36] + src55[37] + src55[38] + src55[39] + src55[40] + src55[41] + src55[42] + src55[43] + src55[44] + src55[45] + src55[46] + src55[47] + src55[48] + src55[49] + src55[50] + src55[51] + src55[52] + src55[53] + src55[54] + src55[55] + src55[56] + src55[57] + src55[58] + src55[59] + src55[60] + src55[61] + src55[62] + src55[63] + src55[64] + src55[65] + src55[66] + src55[67] + src55[68] + src55[69] + src55[70] + src55[71] + src55[72] + src55[73] + src55[74] + src55[75] + src55[76] + src55[77] + src55[78] + src55[79] + src55[80] + src55[81] + src55[82] + src55[83] + src55[84] + src55[85] + src55[86] + src55[87] + src55[88] + src55[89] + src55[90] + src55[91] + src55[92] + src55[93] + src55[94] + src55[95] + src55[96] + src55[97] + src55[98] + src55[99] + src55[100] + src55[101] + src55[102] + src55[103] + src55[104] + src55[105] + src55[106] + src55[107] + src55[108] + src55[109] + src55[110] + src55[111] + src55[112] + src55[113] + src55[114] + src55[115] + src55[116] + src55[117] + src55[118] + src55[119] + src55[120] + src55[121] + src55[122] + src55[123] + src55[124] + src55[125] + src55[126] + src55[127])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31] + src56[32] + src56[33] + src56[34] + src56[35] + src56[36] + src56[37] + src56[38] + src56[39] + src56[40] + src56[41] + src56[42] + src56[43] + src56[44] + src56[45] + src56[46] + src56[47] + src56[48] + src56[49] + src56[50] + src56[51] + src56[52] + src56[53] + src56[54] + src56[55] + src56[56] + src56[57] + src56[58] + src56[59] + src56[60] + src56[61] + src56[62] + src56[63] + src56[64] + src56[65] + src56[66] + src56[67] + src56[68] + src56[69] + src56[70] + src56[71] + src56[72] + src56[73] + src56[74] + src56[75] + src56[76] + src56[77] + src56[78] + src56[79] + src56[80] + src56[81] + src56[82] + src56[83] + src56[84] + src56[85] + src56[86] + src56[87] + src56[88] + src56[89] + src56[90] + src56[91] + src56[92] + src56[93] + src56[94] + src56[95] + src56[96] + src56[97] + src56[98] + src56[99] + src56[100] + src56[101] + src56[102] + src56[103] + src56[104] + src56[105] + src56[106] + src56[107] + src56[108] + src56[109] + src56[110] + src56[111] + src56[112] + src56[113] + src56[114] + src56[115] + src56[116] + src56[117] + src56[118] + src56[119] + src56[120] + src56[121] + src56[122] + src56[123] + src56[124] + src56[125] + src56[126] + src56[127])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31] + src57[32] + src57[33] + src57[34] + src57[35] + src57[36] + src57[37] + src57[38] + src57[39] + src57[40] + src57[41] + src57[42] + src57[43] + src57[44] + src57[45] + src57[46] + src57[47] + src57[48] + src57[49] + src57[50] + src57[51] + src57[52] + src57[53] + src57[54] + src57[55] + src57[56] + src57[57] + src57[58] + src57[59] + src57[60] + src57[61] + src57[62] + src57[63] + src57[64] + src57[65] + src57[66] + src57[67] + src57[68] + src57[69] + src57[70] + src57[71] + src57[72] + src57[73] + src57[74] + src57[75] + src57[76] + src57[77] + src57[78] + src57[79] + src57[80] + src57[81] + src57[82] + src57[83] + src57[84] + src57[85] + src57[86] + src57[87] + src57[88] + src57[89] + src57[90] + src57[91] + src57[92] + src57[93] + src57[94] + src57[95] + src57[96] + src57[97] + src57[98] + src57[99] + src57[100] + src57[101] + src57[102] + src57[103] + src57[104] + src57[105] + src57[106] + src57[107] + src57[108] + src57[109] + src57[110] + src57[111] + src57[112] + src57[113] + src57[114] + src57[115] + src57[116] + src57[117] + src57[118] + src57[119] + src57[120] + src57[121] + src57[122] + src57[123] + src57[124] + src57[125] + src57[126] + src57[127])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31] + src58[32] + src58[33] + src58[34] + src58[35] + src58[36] + src58[37] + src58[38] + src58[39] + src58[40] + src58[41] + src58[42] + src58[43] + src58[44] + src58[45] + src58[46] + src58[47] + src58[48] + src58[49] + src58[50] + src58[51] + src58[52] + src58[53] + src58[54] + src58[55] + src58[56] + src58[57] + src58[58] + src58[59] + src58[60] + src58[61] + src58[62] + src58[63] + src58[64] + src58[65] + src58[66] + src58[67] + src58[68] + src58[69] + src58[70] + src58[71] + src58[72] + src58[73] + src58[74] + src58[75] + src58[76] + src58[77] + src58[78] + src58[79] + src58[80] + src58[81] + src58[82] + src58[83] + src58[84] + src58[85] + src58[86] + src58[87] + src58[88] + src58[89] + src58[90] + src58[91] + src58[92] + src58[93] + src58[94] + src58[95] + src58[96] + src58[97] + src58[98] + src58[99] + src58[100] + src58[101] + src58[102] + src58[103] + src58[104] + src58[105] + src58[106] + src58[107] + src58[108] + src58[109] + src58[110] + src58[111] + src58[112] + src58[113] + src58[114] + src58[115] + src58[116] + src58[117] + src58[118] + src58[119] + src58[120] + src58[121] + src58[122] + src58[123] + src58[124] + src58[125] + src58[126] + src58[127])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31] + src59[32] + src59[33] + src59[34] + src59[35] + src59[36] + src59[37] + src59[38] + src59[39] + src59[40] + src59[41] + src59[42] + src59[43] + src59[44] + src59[45] + src59[46] + src59[47] + src59[48] + src59[49] + src59[50] + src59[51] + src59[52] + src59[53] + src59[54] + src59[55] + src59[56] + src59[57] + src59[58] + src59[59] + src59[60] + src59[61] + src59[62] + src59[63] + src59[64] + src59[65] + src59[66] + src59[67] + src59[68] + src59[69] + src59[70] + src59[71] + src59[72] + src59[73] + src59[74] + src59[75] + src59[76] + src59[77] + src59[78] + src59[79] + src59[80] + src59[81] + src59[82] + src59[83] + src59[84] + src59[85] + src59[86] + src59[87] + src59[88] + src59[89] + src59[90] + src59[91] + src59[92] + src59[93] + src59[94] + src59[95] + src59[96] + src59[97] + src59[98] + src59[99] + src59[100] + src59[101] + src59[102] + src59[103] + src59[104] + src59[105] + src59[106] + src59[107] + src59[108] + src59[109] + src59[110] + src59[111] + src59[112] + src59[113] + src59[114] + src59[115] + src59[116] + src59[117] + src59[118] + src59[119] + src59[120] + src59[121] + src59[122] + src59[123] + src59[124] + src59[125] + src59[126] + src59[127])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31] + src60[32] + src60[33] + src60[34] + src60[35] + src60[36] + src60[37] + src60[38] + src60[39] + src60[40] + src60[41] + src60[42] + src60[43] + src60[44] + src60[45] + src60[46] + src60[47] + src60[48] + src60[49] + src60[50] + src60[51] + src60[52] + src60[53] + src60[54] + src60[55] + src60[56] + src60[57] + src60[58] + src60[59] + src60[60] + src60[61] + src60[62] + src60[63] + src60[64] + src60[65] + src60[66] + src60[67] + src60[68] + src60[69] + src60[70] + src60[71] + src60[72] + src60[73] + src60[74] + src60[75] + src60[76] + src60[77] + src60[78] + src60[79] + src60[80] + src60[81] + src60[82] + src60[83] + src60[84] + src60[85] + src60[86] + src60[87] + src60[88] + src60[89] + src60[90] + src60[91] + src60[92] + src60[93] + src60[94] + src60[95] + src60[96] + src60[97] + src60[98] + src60[99] + src60[100] + src60[101] + src60[102] + src60[103] + src60[104] + src60[105] + src60[106] + src60[107] + src60[108] + src60[109] + src60[110] + src60[111] + src60[112] + src60[113] + src60[114] + src60[115] + src60[116] + src60[117] + src60[118] + src60[119] + src60[120] + src60[121] + src60[122] + src60[123] + src60[124] + src60[125] + src60[126] + src60[127])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31] + src61[32] + src61[33] + src61[34] + src61[35] + src61[36] + src61[37] + src61[38] + src61[39] + src61[40] + src61[41] + src61[42] + src61[43] + src61[44] + src61[45] + src61[46] + src61[47] + src61[48] + src61[49] + src61[50] + src61[51] + src61[52] + src61[53] + src61[54] + src61[55] + src61[56] + src61[57] + src61[58] + src61[59] + src61[60] + src61[61] + src61[62] + src61[63] + src61[64] + src61[65] + src61[66] + src61[67] + src61[68] + src61[69] + src61[70] + src61[71] + src61[72] + src61[73] + src61[74] + src61[75] + src61[76] + src61[77] + src61[78] + src61[79] + src61[80] + src61[81] + src61[82] + src61[83] + src61[84] + src61[85] + src61[86] + src61[87] + src61[88] + src61[89] + src61[90] + src61[91] + src61[92] + src61[93] + src61[94] + src61[95] + src61[96] + src61[97] + src61[98] + src61[99] + src61[100] + src61[101] + src61[102] + src61[103] + src61[104] + src61[105] + src61[106] + src61[107] + src61[108] + src61[109] + src61[110] + src61[111] + src61[112] + src61[113] + src61[114] + src61[115] + src61[116] + src61[117] + src61[118] + src61[119] + src61[120] + src61[121] + src61[122] + src61[123] + src61[124] + src61[125] + src61[126] + src61[127])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31] + src62[32] + src62[33] + src62[34] + src62[35] + src62[36] + src62[37] + src62[38] + src62[39] + src62[40] + src62[41] + src62[42] + src62[43] + src62[44] + src62[45] + src62[46] + src62[47] + src62[48] + src62[49] + src62[50] + src62[51] + src62[52] + src62[53] + src62[54] + src62[55] + src62[56] + src62[57] + src62[58] + src62[59] + src62[60] + src62[61] + src62[62] + src62[63] + src62[64] + src62[65] + src62[66] + src62[67] + src62[68] + src62[69] + src62[70] + src62[71] + src62[72] + src62[73] + src62[74] + src62[75] + src62[76] + src62[77] + src62[78] + src62[79] + src62[80] + src62[81] + src62[82] + src62[83] + src62[84] + src62[85] + src62[86] + src62[87] + src62[88] + src62[89] + src62[90] + src62[91] + src62[92] + src62[93] + src62[94] + src62[95] + src62[96] + src62[97] + src62[98] + src62[99] + src62[100] + src62[101] + src62[102] + src62[103] + src62[104] + src62[105] + src62[106] + src62[107] + src62[108] + src62[109] + src62[110] + src62[111] + src62[112] + src62[113] + src62[114] + src62[115] + src62[116] + src62[117] + src62[118] + src62[119] + src62[120] + src62[121] + src62[122] + src62[123] + src62[124] + src62[125] + src62[126] + src62[127])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31] + src63[32] + src63[33] + src63[34] + src63[35] + src63[36] + src63[37] + src63[38] + src63[39] + src63[40] + src63[41] + src63[42] + src63[43] + src63[44] + src63[45] + src63[46] + src63[47] + src63[48] + src63[49] + src63[50] + src63[51] + src63[52] + src63[53] + src63[54] + src63[55] + src63[56] + src63[57] + src63[58] + src63[59] + src63[60] + src63[61] + src63[62] + src63[63] + src63[64] + src63[65] + src63[66] + src63[67] + src63[68] + src63[69] + src63[70] + src63[71] + src63[72] + src63[73] + src63[74] + src63[75] + src63[76] + src63[77] + src63[78] + src63[79] + src63[80] + src63[81] + src63[82] + src63[83] + src63[84] + src63[85] + src63[86] + src63[87] + src63[88] + src63[89] + src63[90] + src63[91] + src63[92] + src63[93] + src63[94] + src63[95] + src63[96] + src63[97] + src63[98] + src63[99] + src63[100] + src63[101] + src63[102] + src63[103] + src63[104] + src63[105] + src63[106] + src63[107] + src63[108] + src63[109] + src63[110] + src63[111] + src63[112] + src63[113] + src63[114] + src63[115] + src63[116] + src63[117] + src63[118] + src63[119] + src63[120] + src63[121] + src63[122] + src63[123] + src63[124] + src63[125] + src63[126] + src63[127])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68) + ((dst69[0])<<69) + ((dst70[0])<<70);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h388e1b676400777fa0433d1630d9a15d84bb4ca40e82a4cfe68ab22a7e53727b77af33b847c5a47c37c190827eb77dbb7ffac6a7d8365b6f8b05cf036bb30bcc0a5f1666bbf0dd136279ee87b6086cda5438956fe87ae4676adaf45214ebf0e3cd32b388176902631fdac90567a39ed4287e8dd485a20dd82da1779ca52909beb9b179c5622bfdff378bff0607b6064235758dcc8a28c51cde94dd93f7153d38270dda4ebb92b97b6bbd2e637e277b6e5b528c9d3cb141f282c695fc604026371f04d01191e10c4c331facb6642661337a852f0e9f285dc3a28c01a8849b2cc26663fe4a93135fd34c1e496a51eee1c9bf8272a2f2b0b1aec438284265e79de64905e42e53d81ca8033c13f562a13b3142d2e394fb015ee04fd2045aca9d43661883fe6c48fb8b1a72e760dfecc19476a9965145837b5460c30e5d6246d69d82719ba9033572b30c408da7e395308baeccbb47f39d1a239d68db38c1b7ff6e1de910596de5066ee296541dc164e9ebb32dd8c4f925d52618bbf31969cbb2f86d0579fe5e4c6f3fd376246e9c25bcd06d657c15e476c075469d0e14dcae564a08a735a46dae7e0f63307f885481278773cffff3db4aae0e1d80c0218e981657a4a9f1df4a400ab3973556c68ad3c58872a34bdc4e322069eaf4f4a861051204fbe062d5246e6d1a520c27622622997f79d10734b1c1254305b5e94466a47e80f84bdb1bc8a2f8752907010e363b883f4f4374dbf5abad785671fbf0fc123108c0de49b9fe5639e8ede3d767ba03cfa446d5e1474c6bf5fa3873074f21af4c218935cfbefb3fe31f837e44623bcdff344b459accf0f35c8b54d6382476caf7080a1526234761c1ba39ef7d245a90cfcb7ee7e04cb2b37b938b1ad54824c8593405d7a690622f1bd316d627c46bce2cd202c7e9a19caadd9d61afaba32d800345bff29e0a2cd3eda14f19cf21e5fb1eb6a72c1bf024e45562d4bd1351d9e99c697de7deb8675751000360758e610748da80f565188918cb2cd65081e8074a957c2740c42d87cb48d69f8ddd307e4e0ee4a3e96a3fc6326fa94ec73210ef87eb4ea6f38e871d7312697299f6f6aa7fffb73068670a8ebfcf49b679c10527b6de3f5c842d20b5e2abfd78f8a973bed71b28cfb39b175223708b1a728695807a9925c6ef0e3fa6f8c23f5fe542394ef7056ed5ef1cdb92a14e3ab98854635fddc592a3046ff5aaef71129f6decdbc17c3c22fcc1bf480232a951bff0b9a161822f306acbc30f7b0b8b2f8dd61771cf10e9e20c870bc4c8df596ba8a7e7a2f6b3ae5365c586fb8f4c3e7aac51f60fd40dec666e741a83ac8c0e3f559ce559f4d6e027c21be0e244ed28d8442425952ff6af44c99e05bb1322be077917124d90398e0e9109dc4f36e425457035cc1e822b4f2a6137510ed31fb6f0a096c9e0de9b673bc5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd1e47831ea053941302da074758976384c4b43ccda8910bd29bdd0e01bf325e72b2c1a4ecc27cfecb9bb8e705d29d7f5953852f48c5da25c94a3a291c67d584a12cd442fb444b59c915733c8daa0bffa04447a90f4c6e812a8707cf2db1e9c27c10623f62563b9f5f98cb25a558682f36abfe4846619a6b1f57ce04c6012b982b84d904d49d6e5f1b09659ec1bf0ea1facc9eb6c91a54633403652cfb0c5f5449ef21117f63c418ed82cf16a67ff0c1d718a7c5399a62ee80f961f2f663e5686b647849d8ffb119480d63505015c7e3c35011933266780f938bf188bb68d30e08dc251b73f0cd7bd2ceb8d76829d7f3ddefd0c3336bad746d1e69e5a2f1f241914b5673876d90a3c1ca2065a607cf38bbeb37d14e21cf51acefc682d4f80e92d1efb936dd1a38d16be5a0bb4140b8b7597fdfc947029cdfde3186eb4b0695d03161614409e1e4fb9954ec33909d9372f4cb13761057d5949b6a0f9979e34f5c375d54ec7de1f8b2b92fe94470e14507c44827b40c924465302792604ea2d1be0759d453f88ee70d9b2f70b7e11a31503217902662f437f34a512d2ee9d7a3963d81664633b3599c05d39bf2941978f2115632cee147e5c3dbf851b668c1dc670a829e5ef8f9e451b6567879d56bfedd7c33f25ebeed3f9d9cc5f78993049af8185e92504d6eb42c83e90e87ec32aefd1fb9b87efbd1404877b700c44378e58eb0b689be5d00793b9380d3a197eac4872431f21e71c4ae549b3d409d7444d7f49a8950155eff6d5680265128eef4d2868451703862b507a49106ee82f92e58c3f069fd57ac992f504bde27aa7fc3ba98e620d358bb9ef0fa45c2715d322f3a22dd4e0a59a39fb1e034119061b97e0104b2493b46e7f548438de918ffee5460ac691c1f431a234fdd1f78f44d4b2462eb4cb86a943471ea0cd91c935cd65371bb556bcc0b54975ecbff01336b43ca865085091f56ce56a01b8d6932459aa566eabba2006750718337c816612b2ace65a1763ce1f9b9a69c0605f2404d0555612491b77ee622db7cee3abf62beacd9cf7486391dd1adb706ef1b5fb5e5159aa8e48629be01913c81b54b8aa9e62d8ec3a84c3e677e46d2035c84da06af5c711ab3108d020bea97c39dc2cee1abcb603967c0e0aee22c9cb5d1f2c64fe231d64271bde7fe027edd4d9abb65e910d9cc87b9bab318408bde0700649f72ab9bb7ed4cd36e79d6d3b42be2efa1f676ee128cf17f98d41a39114dd28b274f0439c46ee306706bf85edc628ea21c8a8447bdd38deb1df872e408555e45927c5fc4da71f9e018ac616d694ef47805d80697b9c683b8b8cf6b010e73add51485e0fbb6a777c5643709c5a5acd9d2a88ab3631cd332fa9a514d5451b47fae0e2df544ff04461a9ad2aa1fe4cad47329f80f8358b28db1d16c7264a5bb1ab2c64e9f123f34191;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hacd99edb31367013f7b64c938fed8c411e8d425ade7c17e36de1a0412e36391f8a7d276c0cf72287be0f47b9fe9b0ca7b382122dc02129ee9e924ff1b67b22c05d5b0cf08acdf3a5c931a43eeff120dd1a6da22f2e82895e5dc9f60fed6207bcea4b8c6c37bd117814f27d2f08a19d8db1ed96dac7f34f6d25114f5fb07f4e8cae51b3809b35492ec6a370db6cfe84e46d907516e72c99cc40c91b640d2df4e517ca6ba475967c6f7aa4f9884a0f814fb57b4b8351e0b32f039e13d45a7b317f05c2694ec1f41a27b03cf04727ddced1b47ba3982b52f50c48003133a6619dcf4bb730bf630f8fbbc34b31e6c3b6945f7d9765acc508668f37f73ada1eb69071fc86b74877599e72ea5397c7c3de76653d6c47fb2445d313722813082bba90076f65a58312d4c68458a2e1d8292ca4d8ad1374e810c0a2fd2ef891225ef3421846fb566df682eed31263f245ea7f9380d544a1e75d34a2ec35feba1fb045acad7085180ffdb54dd575e5e2097c4efdedb6e0c4bb7664f18ddfaabb3bd6a3d2f8654b28437b85d9a59a6264d962953b03c94410b4d47b1f15146c7d420d9f2a3a64050cd686e60aa25e4b6890951dd7e19b6d418194d318f026f98f0bed42d6183b15236519f68c43160eb1feca76b48e93b61fa52def6b90c9434a302662073171051f06568b375534be3908a42401e4360b8240637c7c205a66190be0390d39c4a8d80b4ceaac776bdad03abfbe045528ffc192719410826f0478df206975de3491d7282b1671e22ccfcb35400dca885a99a05d014065d6f67a4ea2e467bfa6e28a79c90e7d9518ff0be168bf8b0cd358c67d51344f61940561de28ea0a1079cbef092a890aab297ba201ca96da261c6c7d3d6b2b4daf4371b7b9e1cc5cba0f79542c38a86e97e1c56db0e0e085ba9b2ae373b972884577f7712c51b7cee0f09e602c66a0d03bff7a299027171568030ee39f0edaf287c39af548751c266781fa44f3cf1f6028b2318e51aa25389ca5604ae3d1f705fbb44de51c08f1dd09074a8cc6bbb326f04f924ac570bc856cd869c032d97f3b415681b5dd639704a30d8b73b72275ccd9713e7d2f600726a365b91d6052d0d3a5024a23a52d78baaa80844ec88cc625f19ea80babb7b18929d3fa3a1908b8152e791fc2734195d02a5bfe03bbb238a01b9522a8259f907ad2905789910150158d6f2eef8b39d7122e8b1780188625278ee4946f88c07ed293ca1f9d280cb7a32d33d5f34dc8ee6719bb3ac34167545acd8f00ad903e9d79b168942334095605146f4ff7de15020d51f0bb083e914e49762a6016f5d9a535468fb437c6504963357d2215001ad0030f20066c146368ab9c50f9d3581b8bd8d1f63c2e2f93fbcda5b23cdbdd08b866e1a6d0754c987f24af222fe21a88fba82c0aae15349a2b7e30a3bfae6e78e99306b4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb13d67faae6b7107fc599aa22c17f7c8e01a4cd70b5c076766963fcc343bb0e826c208cb418ef9410c5c2f694600d66e9c652c99c484e837986fe067cd3500a9e439754c7ded0d35e75f3b31605478e6571c01b7f7fd0434bb2801aa21f8ab0a2b6bef2b284e532f5c9db9d6f2d79d76154130de4c131381818c85dac85dd7e805b498544d6dc7fbe1335d3f93aefbb977989d6f77a5851d5e6f2c61e86c186c7c82677cb4eb7e9fa975c598ea0943b5dffaead523756ca48650b96240f19a46df90b520ba482857bfb4021b684a408cb0eef2e82e62e62764f9879226ac306d1f9567f31bb7891ea155fac19ad176282f7e5f7c19c8cdb913c8743e8245efd689739297fc1a756386f1b5181084785120aee3e933e92fa893f7eef54666fe6e24d421e93b1e258ed3c2c1ea81847ea90b1347f9b85d6cbd89fad4dea3ee48976318149152e903cba5d3362a6857c11b1c08972b3b9cf29424ae20e66471c8aa6ce12d4cf7c63584bf8f50598818440ef8b6954293bf2f7951183cd1d9deab03d4aa83c6c10f9585d809ab4afffe6221d68f7ece01d43518b733b582d25f10c468059fceb1fbfac6fe5a19b382267b2ef484c242f6d149edbbd5b2816e66070aabcad9d99495029c83526dfb6f1eec445d6e387f8453297a5173ab26ee7b3d83789e12f533404ab4b2438b61e814a82b3caad60abe77d03b2037e23b9bb06a08ec350a7738a9e8abd98d849c6c5c17d3a33c889ada59ff484be4cd808d0bba0743fc3ceab84a234bb337f05064e2415052caee6dfdfa21d95a74e5a1760a1a0488962a86ce44fcf6925b1761b94a619c7c853ce3002d045d297a1753040a58c91c09e5603a0bd95177dcb7f12ea68061e5679522d34d4f2ba02e5313a86c21dd8016276c1fe0973a0d374e8124c5c54659183629f65fb52d0a8907e28d0e2cc8b07c4120c6016d3e80e00df8863e3fec72edcbac366091f232b1367e5c010f197b6b061ce0e421500d31eb560e711728b88112c413257481ec3c15e5bc30ec70988328438514e1eda5d7a2d34ce22b9646281c80a050af032a2456eb908432684ce13aaef4ba2d7b1d3155aba16492162f60d0f426395d977ec42d7ef782cbff7f0a4078c08b40a0b0f7c4ce610456cc5f00fe61a86892d9c7c0e8d84e532aa72b0afc63c79d774414c2761cf9a4eadac3992829c07614c2ef56aad0795a175c25040c7a5b15ed2c6bd85008ff4589e961d8dd1784da2268f2d30ef932c74e902cb38b0a1b7633aecebfd66319d829d22ec8caac77a5e26fef8facd55fefb81d09e32ce3a2e83ba6322572fd9e0afe8feeddc39b82a34c96e526b451e95303a4021f0bb50b1ccff6dc4ab832cec11a93c1610f5a4c087b60af00bf25b91c50a261b7bf2bee4a6b5e6bf76919a4a28934f07bea7afbed33a73c04b2337825598d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h93960527da3f89a9c56c514f28f512899cf70c86175eddc5e1d050daed24bc5068dc5164888aa3ba2b9bd72ef195a3557d17ed210aec3e9b468bf095f504939db23890005946f061f437b81fec5ec334495bdb7f57ecdb52f4077bcda83f5fa5f5ed9f627c90af6c09c05d053410694c1ad9668552c3dcf7b081ffcd25d92dabd9aeb1a86b81b1ab1b22f1b38f3ae986eae40d2feeefe74eaa0cead0e4416a750fdb0bd314c8cf200a438c9dee3579cedc61533f2a468f7e086dd325aa2995506301dffd6fc5fa25bc777f61b13e717d58f229baa0c3d5107b2ef006152b7a41342671e96971ffece81d8a5920ef880a9d8af53dd7d20438b9d92dea210911190cfab769a3e7243ce4471197052b5c3aff5a6fa3fce828fba210ce393e5254f46dd74c7928de2ee360bcc43f92a7c070e33dc04c5ef9178a8a19e3bf566f993fcdc1dc63d1ce48ebdd5c6b71e825932a67863fb66d7e3ed5398b2eccae3e811f60aef0d70c4836e705c2b657bbee6e0361460cfef5d0bf23a5df01002fcf050ae5906f3ccf00b384e23f0583bff5fe68d1658d57725b188c51408bd370714ce34f39ed25e9f1199c5027131f37f1498bed7be5d3717f016aa45acdd41a6762d4345b62f9253d35ca65c9a5aa12b6b9864129a40555822ab9a34c91334e70fa7edb6409ae59395fd9b939eb2b1772f5393585d968027634607ef2efab0100683e6ea2414c7e79ec73d7ffdd012b0be1736689e35233cc849a43640d9da5b039a2ab632955561284bbe8a81accf9e3f06ecd6f88d8eec4f48b2a4a386c2a9091b4d48eb709244dc21a9f8917dea298b796de3023028a45b8d7f7cdee575b1550755e2a22d688489d9af03125a59d3d1a2087ed59da25b18a0354f220895578e06e059589cb0dd1774bba9d7d133e21c45b5d41e9c652f1385af9de4626b4014712eb48a3a7c7b99da96c13cf734ac606bde1a49d65da3def770c4a123cf5c5a1115a60bb953078230ebd9f42a27ae7afd5fc812947cd77b2ac21d347a734e2d9195785c73b9fefa09b02c14e79e157cddb282efc227c1d0f4d7ccf294afff6584467cc8c761b3bf4397e67e3372d5d9d15a2a314b632c6913274ee5c66e886874adf6f1d4d9bff72b908b1c0de76cbe3e52ad53faf957bab7fab42b6c6151d9939f1101046953c521e3935290c01e40b2b57673b1b88a5d4decdd8ce3a2ee152a80f3e35b102c02951fb761d87009f510753c51ea44d16a7afd7f482175835077642b8e01e2f6e48b445264c5498a613c24c4f2a882609db19d2cc353ecc8f32564c7ab9341d48a999ce12443d729a3b26cbbb9d6c3842b426ef0d6c3126c3a04e5bb11f6aaf1163219c77176deb5438df694950ada9ea75fc3cb9f509314050bc048207534a43e49de28e3230b35aa5d4ede0fe33791542e714bfe721da4bdfd9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7e0b895ae9ec1a05504d4d49b41d9ea299ec3f8e7c664d4381522b43b76297bec339c9314eac9eb026abfc7710aed7c8a542ec8525ad0a7eb266af4d33d73f147e3b7b49caf8b891c12d0319bfd99b635f8404a2339e792532be47a7f22707b0f66f6ab9d73387e36ef5d04fcac997b798f6804b1a408bb9e858b365a9d99397bae4a0db64fca6fc55c52e30df4b1daf4c12df2ec9a80ed610de1ced4d205f3cacfb82b2efdce613afd8e54b4f1c9d56f2a025b6e1f56a4e74f19e3f1921950fa90abeaaada247ec4d4f59bb0b8045ad221e78f38cbaa4c1614ed18693dfe8f89d96822faf4a3b0974c6bd3fc4a565fd25cea6e16bf77b7f53ac50c4c723ee7c9ceb0192480449080dbce0910b13b6560633500ee774a69cc08b043da7f80876a35b4baeb034be5998f4635115c2df59aac294fe47be8733a55432e80eaf14d0459f4d1f235c6315b282ba21b90001fe3f00968b48ddb1efc7fc04c2a0dcaea8dbaad237e834764dd0660c3780f6c1e90494888013292a8389f4ecb335b172cb636b20b8f899816e43181fb8a037745bcfbaf1e7ee7eae471a90ac7f750c3a07569178250028ea339f9322b1563ae896d3322c10eddbdbd0edd9c258cee2f35e76795bc405611a4d2e74c8fc52db1d5b2b13222289e24e48fc9b92c8c68e4b91e2b0a4127d70d5a68334870164a3f81d68c3db83dd03b4505717f24cb5fc6aa43bc203ed0d749fd7e70f3edbd68b4602de45b1c4bbef2a4037d770964c30c325be1c665c663ef9184277c36972a89be778503de5e5ed44ec487a2d10f6c7b18f72097ac67f89b56df3ffe10e8372ec3d0e982bb0e7e1e5853587c0297468eb8fcf09d4d610892f3be7d5bc5b088033b024a543f218135753d62c73972fe67e2fe5ed67576c28c2d5ceffe02f4c95afbdb4bca4a12c8fa6dd875f72272ec3dd8e1192bff68c1b5d3679817361f78eb1419f0086a724d460543e267f61056e11d67a8fab3a541431bfa9cb7b0016d21962d7d080eb53c8ed067b4728872de704fe91e469c16d52e2aba6153dd1a7d24c52162af5c87166c6c2792c205f2c42daf09eb3295c8873815849d14ee0ff490fa392da5a393640f9bc4be069ba49b5ffb47e8bb2ff47a525bcec695cada89dd6c5bea96e44878622070bc07d3e115bb15f36a2748e919c9712e2fd9575a13a016fa891c4f188be98384be556a8cd59b51bf77ad8b0e342ed133f9021f048b01c241120fdcac82a1ff01849407a5daf5de6b8550128cf301102f7c6625315b2548e71ea77b3dd04a6421ba6b8c8115a4d702c428450a6f47e3b86f71263f7d12c00e43cd5fac95f9be7a007d05de32703faa0f42edb3520677df16c997070e9b0f379c256381963add12949f40b1b0bdc4f34e00d29c42b5635ee8ef972144c604ce08f4c7a1c12e93bb5d615e8674a8ed5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h18e41757a8df5246816c82860913331b896c6e9d3a9f9d16693bf43318dfc9a9cc965322bc8bbf54b014cd5ae56b47eecfaf622bab1434dd591b0e991c4b8ae2c96441eafe189e87fcf373e00b94db9fe17345a5bfcb01acce701d611dfac773ee46e8e24e180952d9fa4c46545a7f35e239c65041a775f3c50545122399b599065173d364c58e6b9315e1f1d6c92e7d0ec1582af5ab121209c42d5f0c5270813de226061c49542337739218293546f6e0cf516a817a026253f6974dfd9bf450c2136ee8819216226793e976a607b1947f13c31374db379cfcbe0c6d5e4baa3f3a69bfd2ca3f4aab673fdb79e84c53894cf77dadbbaa95b937995dcb780fb24695dd8eca5430ab2fead220aee234e6bef1ec77290fc37d6f9fbeda9c635aa2889a70a1d0600b65baac717052bce475ae7c39d2f4047b257d676016771d82edf97b01cc8d6573f96d5fcecd52a4c27014e80e176d4fb0dd7da8c781934c4b4d0fcb6f9cd4d65734af347784fa36200988ed1d118271a8cb6e5efe2eb59bb576a0a82cf3ec4b5dedcebb4579a5ec296783c78e9f5da0e53f1899ef142aa5eac9869ff3842b5315e14a58ac40ed44ec8158031e57caff4fb8ccb2409078ae3e256e3a4e2faef6a2316387d1998b1b1a240f3882636a37c0c0a1e3119e2c25fd9d320036d5ae75266852b3d18de2a9fe59a34112992fb90c26785a01886b669e11ae44de4ed2404a4e7486939f9bb6dd5d2cf8b4fc8d122c72be09e4bb34aef3793a8412bf5b93050d0a2926d0aa1dd90d60c75912be51d40053583e54549af12fccd69c70174675e8f79e435e5a79a91e4bc2bf866517494073df0e05e0136e6c80d169ff722e4541492efd0b4124b70c1d6e224ecb349a21bc7202632b9e897703901c9674a4ebc951831fcf867442b40a1dcdc9dcc9ad26abac98ff099b7f2df6b1f61e39eee7c913066069c63e92ce711a6797ac11120392a284b208f8e5d0d3b3368210231c99fd3c27f4ba01c1014c92031c7ea5a845d6c7f3bad5eaefd2b24b98eff2ea8e0f2e1b68ab93d3d6ce9fb55021ec95f9df5d4fe8f6b2982ff522ffcca79ee07a1af6f435c3bbba7599c08fcda76470811f74e9bed7d51475445c341647ffcd863b616ff502da816d3ddd259925cfc2e3bae19f469a823080d19b1cd952de913cfad4ca90f3f1beea9eefb5a1eb67c5425725fc0ab6c4d8ac42d8ec080bf4d0b854a3b41c9f9ff9ba912e5b6c162e984818977670fdf752f9899cc378658692ef2519a50a51952a5b2d6bec32019cc8de138ca3cdf79b394608dc70fab0aa8d9afb4ec7a5c0d92c66f5fbf5a05ca7def10fdbc419f880f8db5bb471364cee3ca4a38d2a3e98723065addd498ceea9d2b38486f166f15117c10df6b9641cb14afc5093afb82a9b900d5e4d91a1611eaaccbc255edd685b90522adc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8b96c27902301e212413deb3941c2a8aded6be675966e52c5ceca54e5840fbd4c40df00a620843d82d10a0dc41c614150e064dd28f51c3f0ee1cb6aa7124dfa491265c8890cd215def18bc73dbeaba447bbfbd2db0cec42054beed322499f0b8a4162ca2e897fb8a899ec3a800413627fb98d5349d9a254d301efac64a44f2118ded7aad91ed4b23a3e0afa1d58a04f1f223d33b99be5b4912bd1a98481746b1f75cdabf7c8502785519efc570a5b4bb3941e743c9f014db0b8fd8d11da3c28d36a84954f097c351876d13498a2eaac3a8ace8b00d094e87151a2c79a31d17547862cf5f2e59b44d0832cf04f4b861fd60010a02a25b4329e94426c7b7a346881dea5bf773e5d20bf648ba473260bd6c4125d4f30af4505885e3e6a48ad44ecb91076f36fbcc29aa12d7abef86319c251380a66f239c5cfbab1b2ff9da7f68788ef6baa22e095cd4d1baf849e23ca95d36b96b079513c6ead5d920469fa1614b0bb966076ee61f0231ac151ea45031a92fc921fcced1b4a303d16db898929439e8778d3deb287fd784f1d0aa57decb32ccda3ff68be1eb8a237ff343c9cb78a9a2d10b31961ae97905ac3ef7a0a0f2355286f46637d2202e61cc187342a1ecd84d25a395df6900837ff543dcd012d50260b146203dddc372d7c91ec55810729a831a5429f7494e82c46b76cc1a23c62cbee55cf07c3ba32cfdf1136181cb61188fe3191d170a652cd8c369d7ffee12291a782c95652cc3e261857d92e766f872f89ffd652cf1857a34976367b3238f9fd10f83bdd0ed4ff25025725b2afe5d51113fe6ef085e39d07fde58fe92ed7f2965b50aadd89ee130510221a059fc177750446c1ae4af227e510655b4933dde71bcb635e669d0e3f8bd99ee67243901b9e9a96467e9a95ce1df83bd523bb11ab7ccabf5a0317bf489d9e52e2f915f8c0413b6879367357ccf8b6c469cd1bc27553af4b9aae39979b207e4c3fa896df9151d63e24b63b4186673e61a85be1738438c11020686d4ec8b918b3d7e89f5c8c8b6fa530b0b5ff4dd18dfd2d4eabbc6c61ae301089193154c7f119eb8f42699cae76e4d49b1374b294711af3daaef9516d2a2bb10db98b8255bc744c27c395af43f75cc8947416695dafc14e52745d142b835b2d474596d24415d7325a0d75557d39846f3cd995bbc6bd2c6c4df7aa30f177be11cb7b752c68bdfbf696f1209b8a8409223ff1d4b442d4d79f5e34ab741610dc2c40dfdf73ce73b1ee26bb5de29f76eeaa53d9be068c77aecdce5ba00219eaf8c1199aba82e18e36b5197ee91aaa17cc2da9d2a4889de3a77b9c96ac94bec96cf08e816754de6c95e09d26ff67c844d36985a7fd3210b0eb87e590beb0b17d6b31ff30519104a0b28bb40c0087e67c5366eefc4c775d08e3bd7c59a6f15ed29e9dd003974dc4ca6807a415a8e0f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h736db0ab136317fd57871c657a9b02ec0572822fd8f079e69dabf3f2b135ff3c97dc7a51ab8945a38ad6b3cf81cc7e8bca33cfea0ff37b60ff2046b57d8128c9f8d9d6b032542d6bcf208dbb4dc37d5a65eea849e266d943e9a32f74012df426af7a2e14b9874b57fdcc8e51188c88f65f2fa5135cb0356d802d5b911b69f3974904e04eac407933510488c0fb8618711dde370f28b5118211333c1946670751d9ba88012105fa6ba6c65a4821e1855daa66ad283f182965658abd11195bd5694942b60a97bb319059546655cec6a983bec8448cfb4e057094e53b6f8d8ac9a4bf7dd32f16e61320361e2980f5bc65c45af784abecfc3a8cefbd7f9f7a57eff72379ac1e2d0122657769b7bdfb495c73e7ec856ef2f1923d3276b7f6f14e0cae1afdb657170254b70062310a2eed47b39131bcd94aabbf14b4d3ab315d4bd6681382d7a65186d17cacf059753bef6e4c8bdbddee3c3b3643b41b3576663492f8f1336deb42584a0f344a2132c53b9182bd9089fa2cc611572cffc7cd94d68b9e6f6b8f05d458e72797eed9e08f13da239a8c59f11124daf7124c6e2f020c126d1b12398f713baa2cba65bb136d7b8886684781db595186e6e8070b027a3f58e02f12572389571539e6db3fd67e9d1199cfc42f16d422b610887156d9df20c81b3ed2ce3da1da41896dd1b8c384300e741448d1fd00d35d0902946fd463d7d03ef6a2acab4937b808bec57b5373f7ae6c233de10d2c7d8e9fe8d415f10cd4e80ab40c6f9d56e90048b655040bb87f0af23860cfe520f5ede2abbeeb33aea51e055440ae08101ca46c7dd24c300cd2e65dcd02c820ef37530f3b940fa3054f967ced1e04aced679fd5cb0324af07435053950cc4516221e90914b55427c71c2d527abfcd879c911082ebcbf2da9f755689baab0c9d1c3d609c7f5cb6f9b982378d0e2284702072861d192bf12bccab26af7620c1c3d3dfc4ff09a5019fefb001cd2dee7db59a46b849c0966a97f18f2374810b246362d7b1139c0d9ef5555ce1307e95c5ea14a5e34d3d0c093f43e0da1cd515e9319ea5b3ae04d5d79a99c945f7c7a03aac025707925406fe89df5332b378487306c587bfc7cf08f8282627dcbcc9941bb4ce60d111adc2325b33a7e90f761feefa9210ccda5212d1eda0bf0d245632ad7dd5534f9ae440075e3574e41657c2cdcc406801a9fecdcc1788a2a8119510a302b3de8187c4d992c1b001aea326d4fa497c1d3d118060cacb820a998b52f1e90a7fe820f6fdbcce1370e5076d8e12e5e89f7e192a768b39cf59da7ae919971aa6cd5bd6cd6de9b344758650cc41a5523a572c463787b85ca1a914efc295238bbf8a2747ef84f3df7177b9f6b0a8246df0dc82a42fcb91d8fc551578c973f40b14c83d90336cd40fd46469ac8d2831810302304cf29b3b193a50347076;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9c5d40e97b41c5250f14b5859aef1c2e54ca6a97230c860209a885504774eb6ffbf4edf8981aec764f80cb36d57e1f19d54092c643f2456baa09015c620c1a0e418df7347764b73c37cf28a2ea436f4ee2634264d3b041426ef33a229b08cf305e1a69cdeba94cf104fea95f3fc72ae36fe0bc3f22e64de190f701a607c58691acffd4957287af1f3887f30dafe4995f554914f3781980f868f2eb2e9dc91790190cbe444c033e31f172d21f2a06e99dd190dda8a54cbb3fab4178671790a715f8a800897bb3b13bc7b7f0bf8dcf2d39342de9f394f9d1ff39393324bfa9d193a50a8c3982792d352b33d234443f88c7e13ddca819b8489d24efa4d50868e8ac2332da430bd345e9598a57ff324323564f890cc600987ffe0b65ea95aa32a8c5f5f7a9604872d9cdce488d3ca4d944d44190ead898cf8d06c474de06ef1f1cb2e1614acfb6d1e43213220e77afa4495fc146a4f064954bb60ad78cf7b5d8ba9553d27ef4ebc77c70a212a27244e49ecce323db89f509a3b1589971a522e30cd75208755e513232e3c5ea5fe4c3ca257ac63963151fe5fa1c8ce07bf00dd1b2d7d7fc08afa0ff1e53109300b2f2946a07219125f0b9a45222ba0a7315c35c90d2258f6b7ad4030c39941a7a9c47835e11700529c94557504ed94771347a782962e25c85e4c5cd13012aa01891d119159b1e6d483b081fce67c8305628f0d9aed0685fff288368794bdbf28c971b08b3038862f2788a57fca0af10c04817ebf006d71ede1938d3eeb3668c53401faf3b37b3bffa418a9d690ec41338726ae28a3eeb52acc633a13af0692c26034b24c2f2a36f1b9b81241b4794755041b201c72383944bc47da0e79c20e40d59fbf990e380c0ca3633c86c9d7472453401664cf657cb6e22a371c6c3e1159847ae394f5350dd2a521ee80da62f95c804de79b39f2ec752ab3b5bf2cbd7eec11a3578743415a7898e962f677021c68ff98815088caced3323e7d9d692b06c985bab099366ab9f61ca95f505d05af3201e7b40b820cf5d9862767a053557a4751db864d084381a81e03f5ff3deb63b7abeab23ab93966a92430aa0d15e98261fc8a6ddcd1c22f0c20489eda6ee335ca4086a9dca12832ecd45b8e0a55efb4c5649d3bb2680856190dda287334c7ab781ae21d9ae23324e4a597dfa7be2af0658d2304b6819891451f668bd43cdf4638b290b6c34627a64d8c57b071c219ce76f9890bde0cc6a0d1184f2403238987b8ff01b1110311620beb5d7a4e2ec416146ecb2a9af8d5e05e17cd455cceb7a0ac6ed5a7f7ec5767edd274f36cb21acf5c63c3241da19708ca838ffd919400118dfcdf352f27d67c00535b680988bc9ee960819f4f7bd0220e1955bfec70b497dba89824bbe0c91b2c333e01311db2cd466a6eb34e6460567c4e91564602f1b33f25868e04b86;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4c72064f3b6cbf81d892f145293a9feecc16dc0e9f5618481b07859d6821016947c1ff3fbc523e58aa66086e85d417cd9d8a1349b7022eba05c44136c75df7b08add4acce2855b7a7f59128fd27404828c2a18f22abc9aba17b3ef2cf94d8e0d2572a169fb6c6b6c40ec6a9ee8cfe9e5b687c64131f52573ba864a10e2ff4ac9a89e6f44180532f8d547f340afa3d0f98ca64e97116c6d155d62bb91750c94ea75341179b49e7869d067577d3acd6401238c0f7e36cacf89e65c9992f35950698f94e10d21f59c7d0d9e525ba21866550c7b517a37eedbe0baf80510437fac3fb2fb925a95c1d22646d8862999739ddc9a1dc0297fe2755257934361e38165abb47c5fc6114d649b3438ce4f6057574d4f6d334f36aa29ff32994e98290fdcbaaef2b430ac57ff40b3c7c85c2e0a71b40f90a72c05e141810939e71bc1eef19360d0abf779031fde91b5d91906a567af4b3ec29994e8bd79c7d742cd70c092b29fba34a85db54e2843d61a9d91b9316aa64c9854e0f552bb9a957afabfcaecf4e84900cb0bc9fd24b97dc28e4067b9a00d8aa113abc1d1aae6eb5cc17c0b5067c863e6ee13c97e6115791767cae3d5269329c4c5ee158fab33fc9c67737e470e93dc3615c92ea913d202de9bd648ca37c9dab099b202cf31e515fb9a9db240f7964c94341f6748db3c95bf673b4780479049c1998ab2ae2deea13dacebecb01a94e8055da76d9f58587374441e1d4547ffed6da0890a5a0c6ed4b0b816aebaebab3af6301e76720a5742ba87534f760f8bb3cd249285f9196428ad933334386a987d482abad3f355fb0e2f574a0c77f2de69ee88ab620185944e80547e98b997f1d4859339cfe833e7630b5143e218f69fad9c36f4d33746ad65f298782e9a651f22d016639cca5fd14ccf1bb5ef7f2d8b662f1ec4e035b9b183f4c848767158b57e2fb36a5b3c5ff4ca9d50b3742d41c53539af1d305dd278ea6a34ce16d412aab61bae7d70a574e0bcacd313fdc933e26bc2d0ea41ba3e6dc0232a06085b21bfd493d4e667ea9575e561b1979ff0d3015e5e565ad8472a03fcaa2ef25f8521f422aa6339399affe783bb4e754bb6848a287b83a1bfc74942415fcceffcb2d80720b29f24106cbf52a9a25608980d9304da461e728972ed23bedef0e2088965fbf61fad80b9d01c5c839f9943df4f5b9189b98dcddd19defed5f0f19441603b9d88ae0e7d619ef2102565a721fccc176455b4c0b495789ef47984f0aa6f05c037eb1f653ea5c0fc582f63384db2b6ce7520a93ee0e4bbaebfb5a1a18c48b3f882cb1a40a8926b12c70eb6b9c4918c53c97d80d27a189c27057746d9cb97c5f4ac74e5e02212ff78a80cacbf9aa7d94756b5a24bed407bc4c6cf20592bec324132c62270bc421cb9500eabf9fcc80bf01565366b663a9a2bbd934b1f7a3fe414;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h56f5289332cbe7bfc1327b8abecd44aa657fcd7b3f1b7ea7f26d4b8800b2680147afa809402269536c7254641641d6125028464a7b699a3c53022d0b7cdcf5e383993e82671d78e56c00eae9cf95a46d1676681180b066412c53086d9cb73c76b53906807ead4f7caee36560762a7968de66ca1db27172a55b961354cdc6c1fd56795a04209affc528496994ff19448dd08dd0d4c252b5c87f7579fdec87d8f8be1cf4e36817e5162b26223ef47d472e708c0015c4265b925eaf33e96beed3e47265fa629eca2385b422925228b2ba45a96d4a07baaf83bae704bdda0fa227a8cbfd57e4a092b7130020738306fefd02380710380ed868388b962b26196900630868b22fbf855ab70f3a7f941dff0089e5fa73f603d1a1a5b1801fb512172948148b82d980863d6ec13ff8219a4e014d0ccd6d3fc7f61dd9a771cade472432c48cf67363e4e5d2675fb9860a53bb868454db1c6960d195f46d5bc551ff4afcdfd7f1492b47d67ce6edb7240461ac3f8c29b92c57e2f0fbe2cc6eef1474fac15befaea4edc2597d48ad0749a11621c3a20abe7e84bb41a003e377cb9e5672b65711dfb3dfe60c751c95c68c7893eec37d65b848842610d8ca1e668fdec800487c1b2e27f24d8dad28dbdf384c011c8f38b6406869cbdc27180dac31b169d6077583c42a0cfb29af952509dcb89888581c637f9b3051e008b1f95114e2acce331b7fc08da29215cf6b3581011100a261785d4cd52f85bbbfd3119d2696bda6dcead17a8eeb708616ab1d172430292dddfffba417868ceb6bf4d75ded876719ff28b74d7668af69ee27d9074d80a2fb91d2d19ff91d9ee375f1251e0ea9a39e65396a327b044713b8294e31d356283c6e42546d8f3695f3e560cb855ce077ebf18b76411cf7f75e078f62a9c947ee1e506661df4300b1bfcbe46009b72b9190529aae18bc180e58f0fc9a00e23de2f2b9f7651941f9e07b49fdd79d4c792c32409cf667d2e1028b170ad1faa31e4957efada16d0612f2ce666658c0a521c2aa3ea831919b949a6c9c5cd72a1ce5ce6a324d2c86946125d11df09a46bb8881f354ae6b8dcb242ba5a3f567ec69564ea096a4f5e55b32837fa0af572f82fbb36493417e2ff6f075baa70ee1f5877e51c87f4e381fda000849ef2009244ef9d901200481ef1eb8e7abd17e1a576c4add9ca005b7b50982cb55a7eec961940c15afb1334441958c6c0c0ad65b5f7b355ce765c0ccf6030d39668eedc8300bc99d3ab14bab693c944e8031d5c8058c99d85a68224d6e47d9762bb25d96bf329bef4a59ae4df297f250c2c82960749c8481565be9c639ef6af4dbe67d84cf690b4c41a7c448487907b9640dc64d95d7329586d8ca3f5f52ba7b031ce8031f0a93c349d931ec591db8afbaa06ae677c6958ed6e01a93374228e131de0d0ed068760a4e7ccb;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h6dbb5d0c5e421df6cd052ea5c62f0cc39dcd4b7168ef6f0de80d97f2e5ba2270ebdbdefad48bc96f5dc3e60b950216a234ef5d956d1a8b74150c31ad02681a177232368a33cc3aa617712c00f24f5754452fcf4c0616a08f5f27467c482a285d85e13eecca4dc746e821dbfc22edd8c9813cdce19fb99399efff82bfd390580daf76e2c717d530e0e18cffd4c7b50f9f169ec4047017ccabab32089fc868e34875cbe7adef9fcb06dfcfcfa21d47738db6c22212ba52880d72ab0749e15b0493cfa75bb9a73d02e7a6801f9b58739b5723069bad912312b71a8c448f17f50209f62ca41aee619b2e9bd49b93e47f5f50578c463fd9d459012df621291c724c0ea2be43e6b422b88ddc5be5ea024628c55de7244d7a535f7ab67eb4545dd005c21957c77592d356280e65ef777d69d6d875b244e138a99c184c1f52662070d622ae63d90ca942db11c60235ce57d15ed92f9c49e4512d0d952e101bbd118cd790569b0d778dc92d61851dc764d7aaa74670ea6be41fbf32e1c5941e8322e7c332e03dc2b2e052a464a6bf6214f7390d7eeda0fc24524f240bb858ba7208965d14aafb7fc44d178239a5a58d309f8ec338fe9174f31bc029e3eaa7c58ab4c045c4e78f4e1a7543ff040aad3dd00656d5938c266fe45006d41c31679f963f232560c017fe2e09c226f824c55ffd1cf4b0d3e8fa8b2abd91ec3cea9906db9079648f440b3af2a53b2da6684e2cb9f06cc8f66b643a2deaf6226139473f8e86981a037143b0139e79306d07afb595fbd1e89a5770194691d17d75e532329486e49fa2584b103bf086e8ea7e1676b837f70a1a9fceffce8be5b41d6949f81b2cda1f701819afe62498620f67cf4e940028c0d302dbe909259ea7486a8badc52cabc042a4361b04d109125217e53e9c10fb171ef9e0837219107097cb3fc44f21e600c1c6cac5f90959166f7d04a289725abcf2151e2da57289e950626fccffa831ec5e9aa6d3ea52513f593b42c038609044b91b923e6ddc85e29a3ca00e02c5a317d7ed0cd04e319414124804b9cf4409589ee5a80c2aa6c94ecb3903cc34c648fcf3b74956fd2cfae8ccfe2fe6c55adf13768598f1ea69aef8f6b381d1bc26076d4d9d6aaad1e273586dc4591f98988547db98961cded5b30d1cd6b045186c75ab2aeaf4456c9b2a2a6b43bcaaf2322513451dae2d1325470ff3d4a2438ed17d7957e287adeca52994cc956187b9ead0387853dc058f235457c5a41f6cbae16982c1eeb7642933299ddbb4d99c50d6d8a04385a847408e0c47cf44b91d97a8638aff1b00223b3c32946f72018a609e46fe05285c02f578e6984f4ffae4469f86904e7038449db0e72f550f837e21187ebf5080959472aa8d5e4f6c62592ca54ef99c132cd5a4659e0cfbbd9888dc6f28fcb03a8b1af8bd4b144f3bb78d60496d44b7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf7c979893649030ed1c3fbc8f6c133498367520aab6581d3aea8aefdb2240def39bc9d7bf5a6b52c9fa713373b496dd3c0e111ed8e574ef778b143298b97c29cb48e5d4231a778be6134b4716ea49c60db8234f4fe976047429cb00624545db04875fb6269836bdbb118984b5c3e3982bb2bf3ac3367bd3db05e56c215725e8e69e2f64c0a13c0ea191cb48b23b3db2b28b06f5a1e0ff28984b798088874f58edac247463a7e53019b7ec761825c22eb07f4e7824eafc6f420feff6ecb0c3cbe833ac7cd19ca01ffd14fff9eddf77bf0ee866edafd105fef8615165bf4231876bff411847a194bfa16e6b46988f23d984f37790b0767efbec7aa70ed5332b4e88f1986b10ac391c8f1cab8aafc94e14f1f2c5547ec6c7024a2201aed0b61a6d65033f517a628bf6d4e1dc3bac4d795b33ca939b58a681a90f22146516cd3bf588951df6a2f3abc12d3ee79fa1875f2a816f7b5efa6dadee93ddaad6a822fb45eb90b2674a9fef16b80c9feb37689618755a96bcfb08f2d05a84df93a895b4320b97f5921c823f895b77ead285e2933b513fb2dafca3dfbd234a1589be05de8dabe7b1abd9e6ed6a657f2ac4ae2ffb5d07de9d730ca5fc8d6d45742bd1b8ae29c7da8a58f8159dc1183a901eea06c6a2a759b5324da3878b9ee1570ae500d780f499b139097dbd4f1b63a0d709a7e1149f504735a025e37c980748c7b4f5e6c14ace17cce8e9df79620c2f5523aaafad3c92f673c06c109da5cf36073c7242d3e1309e1da1b713e5a2b2d0bb7f8117ad4c52191e76e0eb333981e687b500979aa51bedb492e5cef9269e12fc1a51329d028abc77f412ad6bb52117d09a7ca8a4306c511e753bc191aaf395299b6591de6b6f1bf95ded73367a9628cc1a4d9449d37b0d6adf4903664a6fc00efae34104094a5567e8038ee278329d5f35e737f90c7a94f0ce52128751ef0da4096efd7540694780fc450069caf08a3feec80cc6682900c0f6f1f55206e457aed66a2a788486fd7340378afa726479f78f00e29832f214c73f6c96cb49d710ca7284de11cb832be88fbffcf22684716364e18d20053e022aef762772dbb0ddbe6f874daed036e7843435fc73f44e396452f0f3214187630b610b8ac8c5d1a5190ed853056104db6a570cc7a7e5831bc752dd745bd489138bd1ef9c68e89d834ca0a2a93a3f3b4e8c319ae2dec536f0aa4972cd0ae38febb6f1959b6f387152e198d95af43f9ab4e77da42471f08b7ff56a42a5ee90b9a54e36711d6d33a87b20ae0e15f40fed0e8188a52f1245ddfbd4d8718cb76a5d3e9b3e000cf06853f342c6d084480e6cbe91ba183ff1e71dd57960093d323f6779feb4a42f4b1fda64ae880d198fbe431ef87614811eff8167dc73e6ebd900d8d145b6b99040ad81820b235cb5b4d37cb7b93698eb74ff6fb74d50ca8b7d9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb3d249601619d6018f2f52ef2b82698f822a9a67f0f0576ce6a0b03766ff82c0a655796521810ae9e6adfaa04bdbe07c4f1bdd5508827328017f9b685ad524634662500a8eb7061a4454a9e5ce203fa1dd54791ea6dedfe9c1f2e7f3f8fe951d301a383d85e129944680539278234ed2f0e27b46f83bb81b5fb7ca43e9ed315485f5d78e9d2322e5c2c4c95e8875e090d478a3db5795d43dc7a729978729aa618ec5c0811fa85efa79de9b3b2e74d34fd227943482aa9f86967bc67ad71cd87dda37770f18ee9527e57f6afde712af256139a79b15c506734844667f04af2a37b8dc0e1a5bd5b78d80352af8abfc24e66809d16a1dc56aed2b8801d140808067f7bb71cde90e76b67c37d230502a326c984c50e151788a9b6e965f169542834cdb37f22ae5b483748e6d21ef20fdcd69eb4c532c7f47cb2d0d98240cf481ba588b53756e775fa6b8f5cc9be1e6ba2eeed2c35d9269c12da2b41fb7b95e3adefb7054f6f6a2a09e369ea4f4c739f4acdd71f14d2c010a9b817668d2d0ae6cd758adee5357f7555d5bd53d9ff5e0a5f8a3168bd58286a382a33edab9be0c51648a2ecc70a2e91ec766e979e0437c1f7d46bc6a2d87c190e347ed5f6a7062b2f6d78d883d50218e331c3b55864e46d71f04a1fa76cd1a0dd5258f31ef4596e42ef44d638c6bbb998cc74a18762dc29d42a507590d87f82fb45719b7d2682d2ebfc8ba7b8802b938b1b063c30771eaac2a39e66db57462c57c9517791a8d8dba44ed4417030de3d31985d3aadc35c9301a41b6f3d7abaf53e62e8b8a17bd4bb934fb5dccf784d66049de682ea3bbf5b9415959b06d604c60da5bf4b3f40d7ba8dfdb35bf769a52ed6331d65babdb21776667c50cbae64e6d7dc8e09e8b3bb0cbd1aea03163ac43e8d3ab92aac915e17656039f735775386b8aa85d12f4c3706bcf57c5e748bacb258e4daf4e1c983e7dd5df4d989b00e25d524973073f67521c156335972d51c97c402684543af84bc703c8c052f2f54fad0aeada38274f28c43058c6d9eae26db26727600c833e38e67a7eff34889bf22c7f0746e0ce10076f4d8480ba9b3666ffc7a62d562e567c4057559b014ebdc9f070baba362839718b486a9e5a072fd5565a0ae54cea0f7e6f9ce9edab866e569de9fb0982a80ebfb56fbbbb57f17e720d7e9864e4882082dc7fefe0ea133df536e35a4f5679d244c9ec7403a410f52df8a364246817ab302358fa563f101ce595cc20ea733affd756953491e57fb5b689d852d164345859f9b47fb962ce907556ac658ccf0f53697d8013601a902cc38f82c144879e158e75a0b99be8f348d3378a6725f0890976dc9a0a736c7e31fac7aedcd26ce9d7726f4612d54b53569543157affa29bb3d502064b1baef87e9ab8028db3ff91aab467d2077b039f6b23098a1109e502a55fc6bf58;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7bff991dac6234c7a5f13d529739a5436414f3ad936b725b0b36fe0adbf6d14dd88a53de84de8bd6cc685442797949055a6b872929c8feef78f2dd2a4673d59ab2358498d3f2ef696f70b8ff82b3fc278bd1e87bd23b9dff77edd386293a453cb66aa9212dd5baec65a456f2edfd20e6567db3ffb292a7990983d54a457499f20a872290d5765b503a774ddb463e7dd92a5fdbc54b092c2b33dbf573b407ccf66a8e6ff3378d8a097ff1a1893c15f87cf25758cf67e8ea0a8c3f289660797213be4025e7b4bd352a0d50ac721a74a25b4a82f5f43c36adec2c0a480a444365cdf011eb59300074fa2e97aeb097aeedbcfd636e3a1d915aa5f6bb438014756a96e402beb38b12a0d2679be1906c73e0340a3c3b1aac7ed0aee5996dfb8b3ddfbf8f1a61aa2a19044af733becfacf8464633bbf5b73d86888a79b7af6e4d55ae75653f114ab380dae2aa871f46b0d5126f92012dc285da2fded689aeed7ef18fa90faa5fa580bec2e8a21c4872837c29b6c5f17d9b7f94e882cb51da3e6203c14927bdbb20558ff4870947cae972b4354c09e9ae14164c6a17a3ea96fce21787e196450b8881494c004633b2d59e805c4df34f2e6f6fcb3ca563117fde71c55db81812470853f99833a0a61dc23a39ee3484002a20c2c997c890a56eb17d989d32808af162e1a8513ab141c16f4a146bf85836bc895b4b91e38d30a26097cd6e7b0d36e448d31556348021c21d93dc181e887c905593d296ccc07fe2f9fe8b5678ced2cd57e8acbe2daf342e85cd6f03e0f5d4673dd38b4efaee54353276b4dbc36f520f88b3bb2d1810a4ad3effbb5e8b0e923c2fd6546d15b068cb53e9fb8230fe12053f4d69b8cbf0899d8d20118acf40d216cc44545952e272af9a676967e54279c0eb8294d1966c08ae1ca40d63c07b9e74948e1739351a394927c9b3a081531359551eee6688e3496564bbd2be2ec5096205ad1a5e51d8fac41d43b704fe3faae07d4da0a0a1211fc1fb3677f7cc24c8b3e146833a37039a553977c90291e10da0433cb6dc40db7859ef521e6c6acb713c2e15885459dea76c8f06f8d8d66b9ee56363abdf1e240be27f85b8823c4eb41b71dc7c1b1595b69b6e5bfa860043eaf058dcadc850f78e0fc6b699647333fbd9e3c785acd689b1156fc60af71cef0ea0225f132cd6ac04705388ef94dd06b079cf369e8366e71334a47800073f7427e4d6cb40a318e7e88c0c631e9313cefda1692daba6bf1ec52c3c6019142eb79a4dc4a2066dca4dc03a52ac1726e57ac2ffdf0781347a8743113314b59d12a4a65e61b03a65ac2ea9fd203511d0e51ef440d797b35dd9d12370814f8d87c7e7f34965eb124e0671c887d97d2e532af37450e73413500e9007a2c121af10f966906b897e1e90c62521e49686a73b54b67f6addac3a46c7285bcdc79a604b8c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8cb92d347c5eae8cfadf432e374fbb300e04335f4895f85cb4e8d8d98f46d4b7169f07b630faf2541b3f7865316729472c82557a1b13a55b9f4cb5c0c02629ace2523d8aed83594cfde44de6e656033ab6a54eb6b71ca374e5439c70a5ee6f2edfdafece9e203d5aa033afd05fc5246c63a33f3ed5d6460be0b9107c40d3decb3ce330c7d86fffbfa97c6fab0159cae88e620f68de12e3034a139328c84072b61b1ca062a3ca845f04513cb9c9529f0852e1df71d73a78325a19b2cb58698b6261a923da3dc65207ec1c0f64c15868f15be705877b17636e97351ea3d73e557073aea7b7ec7d360ebe015f665d245eac58223599b1d948c721a5f68f59138203aaea0c840954d31107b365b095139f864ad65b41933c6d0cc5adda7560463f7bc5b0a094f716e34a536669e104d0fa47473b850028c59b16c3c32afdb9e952d9a8f16e130d9585ead01581e11a9db793bd10ca998e5deaf76548bbee5a5c92c3a8043142799d01b2ae1b193469173092a21d92922e49236021ae4d4772c2b9cd06c02158859e45f70749221575fb80fe9759874c7846d9174e74d33d6903eb58a0e6879a5b61d5479c33250c9debc78226da7119eed365f40af3c8b0368f987c306786ebd322ce509e904d1dd5f34db77e77feff35c13d507ca54dab22a55610d140456485f41718d3e05a4fcc8686e25b669e9e4330223cf334b4c6227d892faea2267e85a1ba4b89fe1e4a99ae17ab06c83feabf2353d6e8bb863d6594fe5f160cb0b0f3719299765b921a920cb8e2b5b9166dcd81664dba4cc19377a0e5b254b8764dc18f518874925176ab00f6ffcc09814101e9f6d447eb5cf88e6920d2b6a7b9f89c60643009956b03fd26330c12160d0e378fd1a8bf662b3fd3d7f7553e59c4fdaa5d5d199ff05033939a951b42941086ba723842312a0213a7ad38a1b6f79bfe2df37ea20149fb88fca4dcfb07b996460cc110ed132f3da9974c95a2c92b265fe4c5a8f1002581b2daee52aeed6180823d9367eed1228836f9d427f101ed75eef2a0c2bca33134cd42a85e05897fb88726e14c682a04401c0ed02c2dfc5c91bf7d01512f43ca5a9adcc3b38e918d59d05db169e4d77596165f70358f380026bc75e550834314d3bc28ed5ef2103cf37f2acb3385a43df5eb0a95bd90bebb6a4ddff776c61f4b03429d31e7ffa49c50cfc8514b88210826399a50ae52dd0e6e054922089dfd4c6f3b44cc0570af02689cea20cfeb9b5e4697b06d474448a33320a965404fd691f2758b81ca9132824a36449a49524edfc4d2e9f3dd842826a2459c27db7e10db6b89fe0067e53b8e71c5a9de00f789923fdad3dfdf4cd543d8d9cd49e0bff0ae51cc7d4bb594483279b6fbb75cffa7f3d4d85a13d8a393b6ab5deb8799f54f2fc972730055ada1dee256bf986857e97e6e7354947170;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha8b9b85b382e191d500c27a524617e50153a59ac95f6cc858b179fd696fbaa0185a6a0b3c6a32ce1f49c7f469f2a7b31bef89e82abadbba0a92a9a4f08f83c354dd3fbfadec033a2ee77ecc26895a798ad76df3ef7d2c87661867a6ca559fa68f141de969552bf9b5e274fcd91e7efce2ae46c4c79dfb1d0387bdfdd9bbfec22b08634888e8f34b3f7563d0c8d009767010e2e4483ee4ad8b4269d9a2d1713068b8fd6652037d6b2459e314777c349274d102881745572b0882ea2850abe3d9a7f550c70a45a4f76262130b3565ec2cb65d84b2df2a51e23c25fedd02e1dec55cbfd06b6224931e10558e54954f0dc0c87ebcc297ba318f754f6634bd040bff4e5ef092bf051715498eb2c03b51bc674b182c5b45358acef0e5d658d23e407d84ab2bc2e6cfd0f1cb50c23abf54c1047c224dca1130b6b0f8072163f6a392b850d2c639cc20f0e84aa24fbcbd50872c760ae12fbd884d9145b16094aefd0631d34df93527a95774ce7f20f1458c3619711cb0e73d977f7df663c19e173789acc6ac31602ea5661a40980aab670474fb4e2f419b413ccf6f9371fdfcaec53ef27a5b1a8d3f69d83d39ef9226350b8e15561ec56bac74fa90253de8c5546c3f10b5c2cfe2ab725a0319823e225434389c12e8a5834aa4f3f9bde071bf58bf7ccaa43259d21997f8fdbc0c7ab7f319a03ab597cd0f350aa4a002e401d16028f4f222df81a61f0fe1d55810dda38ab50ed76d38f720cd0cb9fd91d873fedcbdc012f6b16198f7da3a36e1314ea7fe2709eaf5ab279cdee211d2eeaa0591b7016fbc733e5f77a0d4c7beddb6c48db08a101bac8ac2d19c73238a686e3df19961d13baee0185bab14e14fa6b91b03974f08fbc64b232ea090e4a493159bf6565151da3e9862c32cc890b5a6d3e6ae627c524bfb9e73bef9f2f1ccdbc4ba938e6db61263e073f3d8a702b0fbf70ac91c55fc48d82a42def7d18c6b3b8bdbc594578d72f4136f2f16fef15ebd383e18a410923db5ab0979d7c6f5b6bcda9e0d5137a187cdd133727417433df26088910c59726679bd74214edebe2b2809f65af8e41b029e98238d1462b11d0fb2170afed268658dcac0993de0b370cf349b9de1902e5912bdd9df7537b7afe624cfa505c268caac9559e0cd2a83c64f42654677f5ddd62cd3aff7858b6e9e7278c49a8adbbd3997e7969e7ab043a35d4056376823518822979867ec014437bc8e1af5e9d60854f0184ead81efb98419a2dcc88d63078b68b9d8aabcc0b0bbbc313fb78731c9d4e3713e5558c04fe21ca2eca7b8c9e8655dc1d561d0259add530b5fd5018ed41ebf23eccb0913ddd2a88842fb9dcccff526c8b291a9053dc8ade14b2c6d550b24629ffe7b6f81cf9df6b479fe7ccd9c1fa9dbb5a94f5e841fe71c24180117a6dd75f51b383197c593b6917c097881c5c9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1e4020c7808783ace51f217fe0c06e9778cdf72049af564e95f46adc651c4f2134d195851698b665f93c893c613eb6806b6e17cfe829653d1e55a2e1096c842d97805f75760de05c3d1b594f24dc60fc2876f1dac91bb772ab9a16bed2761f82de98647a414126cb887d5978928c8379bef5ac3f4a4d77bfaba7da6d017ded482deef046e03bb05bf4cfe02c58c3a067cdcd208d9e415e33e6a2b130f11874d8dd2229d3eb15f4b8491088359d30ce1fa946b9003774698d4a633745f96e36cecf0f2174293fe0b0685ad3dd7bdd1493eb809469ea6539a2c038de513878c023addec93b2114d8d6e66017c3d495b4ff3d487e091ce5755a29c4b6737575f38ab8587e7ab867baa47ac1a1eea3313b4bf9cda6c81058584138ca2d1f454b291cfb4ee4cee55bf73e39f1668db4b7fe7d75df76c8499ad12f7065867863d1013264db39279a0946834b71c8e678c0f3f1e7d4792594670f979864eb9380bfa7849de2df36543da1752dd98a12de39c4f724c05d6be990ef9e2e3fe3718861a0006b192c516bed88916ba221d43eb1cddde02012f4c67d495297d4d535d99f29afdf8cdf9316f024f6c7c1b37bb2255892b50a7dfd2cde3b56a64dc5b8eab31f0bb223471e1fd28e91e62c0548275cff954f213456357f2505d39604a52e25213b9e0b0196cf98ff975c45b5a9f2f915fd028a6ea0da65e9be3d5609d3f6aa0c6345231744187d92c8d5e893cc0bae304968c537c4b9d1f3a18476690ce2d3eebfd0bcc470677ac0e80b7e8d0182a0f0ea60d3cb3c52422db851cdbc5a2a13e5f741e060884e28406b3191adea339d66c63b2e5d91ece67f61cdeb3eeb2fbaa89ed981ed9ae3d411fe3c24c78c7d689e5e54eb7082eda99236e22f55da8ddb2f55a81e2feee14bc5f92881db3626d9365405c9a6859ace101f47f0d1eef1811c32f77422e4e66e5d1e0dc539a813880cd6bf12b83c57cec4dc35613925a1d5fa7c68835a1869572e1e2aaf01861b403ba77a40bc65c0514d0579fd2e19e6a779a6ad1986fc5edb83781ee7844cd602581774be18fae12373e5565724681b007dd0a5e2389b0df9208bfdfa9c2ddb500357080a16e3e08f80c6d4ea059a51d3942a83cf9e8d3a9a13c28e7b95d1a03467847fc4d8e503b8b202fff47ccf3efe7826a25d5b084a86ccf7bfd47a60fd8e8615f365cabb37623afa40db7f5b44719f1597038fe7c74fcc3ca00eb16040ededa863c8a7b6e397f53516cf57b56ff7adcd3d6a3855ab75f32c1aaf9a7f44fccaa742cef6322eecf30f60ed1b55021e1172383393c1fb57f6b5d3545e6fa2bf94b6131b89a62b47c4d98855547c2e2bddd22d9dc6c3fbce68f9c55f5f9438df58d337e87dd88b013eb5ff9a23ac7a0413cdbcd7535b151966ea0e0692602b4131d3fc85427e609120d4845cf09e2fa8fb88;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc82dd0590348e00bd12f728bc61bfd2d0971c88540d2302176dd9b7c466ddb43ad0eaa7b3c3d340150343f9c419fad01c3319b6348e2281afc77a2d51fd819e094c44adcfb168791cb5839f22ac2f0d3b00e40cae32d1866abf2f86435a4dd1208f3db18fc4f9d40dc988db1d4e198b33c8ce99bbe0cc0fec5f3de41a921a60c5ba5147e48c3c225ff5e9327267a12d610f5d7fb50d43f5e4993a50b762145247043b88736b1a38691ab5b3b4426c9b9cf867c1906902e57bcaadb590907d8ab1538252c812062e968abb2395751db15e6fe143812d09901aaac30fb9053d078d42970323958b7509a6735749264e6394ea0e08acfe0c16b9ed6cf947e8afd66012e3496f627cf2e606c655ab86fe9356dbca4c6d1314a195a37b3551f458cd652b5303249b55dada3e3860dc5dd81c659c1af10cd770d82dafddec23280b10d936b0526aeb947bb08ea47750de4348fed003156ef15e4216e98387201f6238a97cc88257abd7c5e053e148431ff44ffa0876fd4f750b6f286ddffb364283fc5b285c50b3d3cc488190926cc7161d733c0fe3e4f56f79bcd4d31300c4759fd1d61b15dd92aab3518a09ef1226efc946630316906b09b6cb890a077cabf92ba3444991c524f8bde8408dd5ef5dda260ab7f4b49d7605b27ba26f27d35f0ad2c2412b434770be72355a6ee0ddf8e0e92f23dafb63a5866b1f9d912ef143cd9e5262103b5beeabe7bba246437958adac0eaf5e12ee25d511beaba301f406a1b8b02068683b4c434c130aa9db76b86fe5415c5afef58db02d72357fcb034a58797080acb9ad84d3a1f15516d4a92d4a445567120895bca4202da4bf703f4a1a16deabd352e9205a182a47773453fd281f2734763d159f1bfb305b06116ce8a47b961d67ee529ac463439bab1c390f70c47e61bb52ef15ca0300aa44a1eb7db4212cb62ce614e7585c7c6b65a1cc7f5816b5861d37302f6882307d22ddcf01fcea9c6170da2badf158419e9dd27eac4b8b8203205555547eaa672f5afa49eb0fe4815852eaebea8282d96cb57c7e03175bd8a614356a53cb73a72f148cc3a537159d8ca49d413b31f86d827a50f539647b404fb540edad95509fda1ab765a59f1ff03904f7651a1851b41fa92f1ff6206ce99e08fbefc5c17104ec60c5192ab1e8e05c31f69c4209ad26898bb95e17c398889f1731cf8a91ac323501ee12c33a898f41fd34b46384d3bccf07921f2b347b4ccccb8bfa70a9ddd96d5036554044541ccf394531ebe4aab26a65c3f0e8aefdc9ffb2a462ca7546532699e1ada301c595f017a144ebc844d1180aff68a052291aad4863c29ab45d787813c56ae8a04b3ea5b403d153fd10a8ec7a73808b24be5c0b9ed51b3c5c290299df3541477044f7ad085004a6cde147d8b4a39068fa51458fa36ca467085cd6b40b50905239ab035;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc4320e7cbb096913b5f54cc1df35959975230d89b953b0ff53bfa8b25f0df7dee237ad818b1e747d4a0ff96e0f660103fae145d15fef57811cf877543809c71368d3a3b454110cf4e35453862c19e7188a1294a94823ba6847337ddd1a628ed31d60d898a1783e7616baa5200c78403eeb99e2cb804f4da5130d9e306e068795c08c22770958e7e0a9966bc5360e29eebff9d885196ba88c28ca165a1f7641fe9244ec6542c46f5ff6489b850a64a9c6ce580f527b46b08ce6c68297aecf4c3ba73c760cef53035f1da61038cb8248f9e58d5deed19149148272cb806671e0bd9b4eae12cbfa2eb5060063910c375ae553ea1d8ceae53fd1abf1f438524126303258a1316fdfa7c1423f0a0df509ba352be8177086e595c3342b1faff10b0b1be2124854550e9909968b3ed4ae42be3ede1e3813516e8742ef59bdf602da15bd8416b0c96048c624e8ffbb79565e0d5ab4ea2e991e52d6916976d02d27f5a2cb023c031936a9ff5ac33bc30a9be816d616876f7b2c4603320a9984b6d467347dc83efa71d85e496936e818d600fd572cd9143c7f4b052305b60add6f8fe05ac0fe05172cffac94e5555c9e3a4d05d14d8a896de8c87dbbc3094399a52a7e6828d3a7e34e39c5444dfbc036b70c71a6bfc534a2211636dd107c2b6e597addda0fb0d0bdec0757442b58250446eb55fb1cb1cc0e476e7bf1c5286419ff238c88dd8910e5cef143744f4c5fe24b203209ae4a99cf2a330447abe677ee5a4598cb0c2e0161ff67645dec5eaff04e6b2bfde3cd9a6d1bc511b42414f42041408616282fabf750510bbe4cfaef080f3f99d746dc3558d322b21a1cdde3904bbc253361f74341646ed0d86d772aff6ffc55dfb15fa2f793691d0669df5282829664a341418a626ef9430a593c8f52b3f2a8dbb7df26dea8c62ee6aa4c4af3f5ee2ddbac9ef884a0b44dcabb8db3d9d3b28d4592273b31f29c0a960a8ce06535fc85a9a256e0963a6b9ecabac71426bde1441c03f2dac16477b57f1561c21d3a7e8521b71a36b1d50b7603435ccf30d34efe416b01acfaccfb59ac08eb1807469c1fbd3c8c021092c2873880df323ceca3d23210c32ee3efe8b1a223f746d7ae465368c8a60cf321ac3dc1592e90ccd2e9534feb6ce96d7d03a093bf98fdc2e30ed1116cd3cb79dfeccfd8794a1bff07efbdf3d89e8ba16bac2e83f5c0f9d687afe5373c235bdc579aa239f37309fffff2f0878d9d82f9abe56e320bf16cb1c8461d2bc4c350650b8aba866b2a63c2e541cd0f731bd24ab9ba4d943c6dcb696d7beee68160b05d6fbffe2d4a397fcd4469460ff0a55577cfc56b636e4ce687e9c20b11933dd1b25228494b505c013cd95f15fd5fcb4b09e1ada1089fcb015cd833feb0302882dc9ba783a1694a2f517a789f7a4ddf52f4fde43352470cd4d8b379dbe740;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hebf12f63b176a89183e0078dc876d1eae9f6dacd5457a915ccf35efdea548fed78a08763cbc90a38fa4b0acdac52aac9d4398a73f8dcc3dc4c2976c3b84f5903d64688f1cfe58056e6e39ebc90210efee236f29e67fa6b1e03b972da02069989141cbe3b643b43182aee9b801270d0dc2faf8518202ff28707d21d6d514b790c7760be50fba91ab3f6326389d4b2ef6faade9abd1d9f73560317ab0a22cd004203c57573a15aa3c589a40ce7277fb6b68ea6f16db6e8a40c3a4560a755ad050cfd4d7b744e10b0267c7b7b2387ca2cb7d5a724c53aba8b797391737ef2e09ba09877467e3688fd19494811ac2a44e0119ac0e55e254210e42641982e0baa3a35af73cc7be3e7311b0cd69c37f71ce767061eedbcbb0a3b78965b7bb5c98db853ac07411d9699737b330d4c8d7a0debebfd87f2628a59c32a24b1e473052c78498ab680b251fb508e7ed180b059d98b647dfcc1e4645505eb46f9821f8560428c19505f30c1acd13dbd3180f0daaf42c5a327b7e395473d975667c86706c5e8d86ea5a31d1b748bb6abe696d1050166c5fd6415e0e0e8286d207b48a3a4bf26cc5d786b395d36863a67ce4652426a592d3cd5b48277c350ee22c0d53f506956e299b16a3ab8d790b57c1bb70987d52a5589556795d52f98a5bc3b0832d8582573aedd9713305e1c2c635596cd8c12e9f4fb287d76f1afad344ec6eb13bf2b51f335f1d3e43c64b809bd0692e15dc7720a5c11264d469cc734c4ab8e19687fb4349456478340ffa20ff3a44659c90aec0530456b3ced66c80d8b08f2763dac23e398f8ae5bb175c1c75d2fd6c29247835b12e31d457da60557d558695f801211610a0bf54bbf024eb09b4ad644b632c25f065d2166b333e6aaf19c9ee9b1001ffe12e18ecf74a05cb1db1f1c80a89d8b12320da243b1e8aa208f693bda041b8d0cc196449ba0f3616cb35e02198f7e32b0ba254c0b5d687d143eaa0d852e7c013d023bd1e9127d1ab657cd012e6bcbc2d77c0989769a2b3f3fa7cf51301b151ed2b8e614a0a0f2f9cf122c73e568b9f602842497bc9576903accece3a876ef886a998f4c7c642ed4663c07ed20629ba62255dd5c0c8bacd8270f8d30f88a005cba3c643d83e19b413721159d66095886bff14b55d2363cc45874ee59a35608d2e927a5087d54d64c9df39d77ca1805c83f0573f631e02329e5cfd24bf2486519ffc1bc2fa3483a0db3eaa28dc2a6a3c220b90e8e5c5a0616cc9c79feef280977bdb581e69e70144030085c208df06d5f5e43e9c75aeeeac6b248db8047a18916b88bc7de1389525124524c6eb75cd4ca07d53c1647b7cc82ed1c5b087959a52e44abdf40a7bcbaae9f4706fb55cbabe3b05265351cc1ae39bf57ccd1e60f535b16edf1ff9f13ab15ed459fe4aae1a3ab745f50f5c96fc6cf9257ed8372ebd98674;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9d34cfa576e0581a4513b5822cb2fb5fcf3672952b98f3d8b9eeabdc76ee403c4e3533476018b912b9b055a03553b838c92f06264acef18a7e66c5326e8b3f761b7ba66801c47ad39fc5e92e6b03f40fe5b871fee85dc4bed09aaca7064a3fbb177bf228e9516bbf8ec80c597b524cef802351edca6aee95792802fc31e9e8125316698de88a8805cbad81e80074711676093e40daa904aacfe43e0488edef6f9f5e5d81b1cd7b52da18ee23a35554b29171498237c8d74d4f29a7dfccbbdf99d8c7b9079190873acdac6495208a14e19ded9f8272455dbe383fb30a408848d6952edcf5b540295f654300210c48ba9c13717a69c003ad9b834579ca16d9794d37f012b9fa85e304ad75a0becba5c5a8cae44eb856e5974354a33f37a68e1c35ee20a485011179b77c6338ee0260a9c53762ac8f9781910400ee2409b93c2fab55f1df53f1ca6d46eced6c68cd6c8639a540b321640ee5bcfccb72c5ec569ab782259766d7e58d13acd931d184f506ac9659a50f6289988fe631caf5b510ef17276494bd30372ac21e4521596cb286aac4a978824abbb84f8f8953f048ef179bb4b9d45da7af98f085ea221bebd02af295eb944f9a666b0ccc66ef822ba9ae301fb0ebaafc8f3416d17a60851f5fa98477c58752f4eb1ab0817c02fa083b01d7dd1a5e9cfa1170ce574f2bc727537930efcce3e8a09af82c8cb327350c219d974d5ca34a1c4836c04edac1ef7978e4f5c8354f4637afd667b7c190223c2019632cbdaa87d24cbc74511851ff0a1cdd2d711ba2bc1b47e8fd29251a70c5f0b8f06523ef38f2d4a55b86a546822c8b499832e7f668dbf7ccd05ce7e64857b8fca893bde1082b8deccd5b35011f320da530865675c162ac528ceb1f4c8a59d2b87da1586710928c1337a9a7e36a2db2d0337cf5eec966b95981a2f7cc53abdedcb032661cd325fd3f6adbc43fa4ce0715648cf0f16e7c1e21efabee351784e8f81651d3ae521e652f87436db22f81a663c37aae12c4e0c547a99283250893763b2bb3d604895740952ee750078d4489060cab82b609ee631c19493746a7f8ab4d80e6d727ee0891a8e2efbff631e02ce8fd3c355a726ee206f1590e89d81c9d33f6223b78df8a9ac42088634a390a38bd863b7f7840a0a23d444505a4aaf2366ac32f2a5b53402c512011649dc37bf53dc6a2be2bd9f3fb8d9d7f4ee190831810e1fabc6ea07f2b70f4dbb504fce3481a1942fbaf841311b4b361c9f5de7a72dd30195ee54cc14b4613e44d833911dc6daa185f001a8ec3ffad491f2b07d0427ccef61229bfc6e62212d9f5f2f819acf3eb2573c02855f3da0875b8fab563e98e76b9c5629aac0706182cfeb021ab3a64d608702b96dfa2e239bd1b1e09bac298b8959b8599f9c9b195df75ecba50177818c0585fbf36791f69981bc1a1f713ded;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4a6b8cbb8b8e9eadd312ef88d43c0dc4fc875047ee116ee93cfcd08d7822529a7f485b8771fa61eddf652f10be3b041fac397417630e2fca2960f948955295e28a635a51f3246e901cb22afd924c4a4e68abb4482420aa5ba26932249976ae07433d9f4c40bfa0565f8b8530d64f4468ba98ff978165bc8cf4b52d406145d2dd0dc8e8dd9ddd90637d17711479692df2d6fdbae10f6176846910db2d95df62d8ec18e16c1364e48216956258c0316d9b88f30b2ef588dae467e74d92be81117b01017957bab08dcee3392151401dda5ff46dc81fdb382dcfb09bd7ca8181f21ec7eb0de0450b9c61467a094cc01f7b71ec7d5e7c23d5551dd85728b6b465f6b3b055c782a414b38b4abb600a08c9d528484d08d153d29246b12ce7f56d351c052b849bb83d20f82f24cabe24b2a9b00d84c86f034384f01d4f746571600e582c5790dbe89db52b6137ba9980722cd056283fd6299f3c8659018409b8e06b216eb6816c5107c1a66c60f6d9028e4603857b77afa4ee08f355a04c929ae63841ddc7099d1e866940a2245da0eb5b1e5e6b1414aa3976a52e26b9000c66b309adab3a76f154081c0d1163a80fc5a49d708f6e237e1c0f22e4e3ce8496c7d5f13ce935cb2428fffc641158b01ddda0c75b85a1c1aff5569f5e70e715be593e82cffee10a9b68e49e9a260bdf0113d99681dfa2c1bb767c6c332cbe625857d79d220f836d68b8deaa114c0d830aac75d20ef25021b391ad828b70e56a36e064f6d2e7103ed5d350767e57cb82c85beb914dc5db555716e0ec01d01487876b8f45af2c931ccb7b8494d18dc155527722a9e348297e68a878744edf0fcef96f88c5f6df30be428aa88abf78b28e02f16ff28207d553620310ddcdccb6e4e3bfe417acbf75bff0e04d7e89169dd08c7f2ef4c17e58e7490c875b345894734cfbb1e35a800ccc3347b02d11ef315dcb54228229728039a56686b77018d089a41a69b1c873875f62734409107c7d42cf2b862ff318f997e399df6d775be252ecca0e02355e3a2dbc5024b5029695827ea313f8a230a7ecab2b3250106849d3a6639e58106d4b661feb19d73d26b757ff861fb9881fc91a4c3fb9ec69fa47ae09ed4defd0bfbc65515f118ff71add3112b28a0eb473ecf8dc574d0dc96d49ba2463abfdbc16df6f16cc6e0c339fc665e0b5310a7f8569ea40f13a6c2a01d2ce34ec89257833204f1078abca7303e1200b36a1bbe9096bc5c49501de5b58f03c412969f1559f2363e57f3c1ed5ecebce3446575568fb2cb59864a4026f307d24416010e941559eef871163bbffc5c5a8af18e004d323c06a93170d586b6dd9d93ffc60c263f44182e465a6e783d1357c247e66d6095a761ace479fa99967e6254951712278eb4639840da846fed26af1af4b672ff9c14b1c11e7ccd18b7a838145d0f9dcef17;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h36450e3d2b4ecdf75dcde7e045f782924cb70ac4a5a9c8ff332d12bfff58157abf99f01e7afab4942ca059b44f0750061afcf32fc02b8eca8bb4ed87b6e51784f80210ee417e513a07b1ee1e7554d8ead0317af812664460f21ea4176ca1bcb85bcd597848583e6d382afce88230907f2c90265a0a88b7a8afe8e4efe0d2cf0479a2dad5bb2a910981813a03227ceec8160d0b7ee5c1545bcac9d57be949f41ebb50f14ce8849eb2dd844f7b4ff31a1385d9609ef4919725bca7206dd217a53ee9f88a374b25c6a69dcae529a4a8ba4a2346dada56085cd98e6ab6caf99d4251f6c9a2a8b01c241292ff5d3c796ff30cbdaf7dbf053b2f81167e13cef1beb9e08c230c6729f12aab090ea154fe0066c4ab51c6bdc3bae8dffe5c10294b7ab5661baf1eaa0be951e0a09dfc0a94f2b1708e999543a998d00f67d6bb92e397e6e08851f9fe758d2e1c1fd93ea655a03a92e779af2d3ffee7e63c01365d8a2f6ac34f2dbfbad05e809409b8efeb3f77e4f7af2be45d55492070cd9a730962650de3ef730c53c4be961a9ed8178fcc86541ec2444eef309fbeaaa0953aa5d1d212c8b725c59d5bc74beda4b8e61e7ee15fc430dee86b08cc5e8578ab803015f34f00b2795cb309e9660399207cf303d87a3848af01408a0938a73612b87bf5a6bb8c273f4719389c7db064416026d875d7e2ffa5e77dac6fe96c09ed5842e43800f4ee1d01c0b4935abf68367eccc808166a3556165bc4f819cf25af3e92a9e98c20a6c85173e7c73b9af160d335656ac7ff501dd29e717a09d956e6568a93354597e46758f658fe617f8bf8c16a55a25687cd1fae9daea8989254e7d8e94fe7498aa6a07614ed1f52fdb502582685f5debfec4870b8c89c5c63a99dcdeb1999e06707a8aad8bee61a0a9105617c24ae83fa3eeb06b091daaaf2a179be49c911f0f5a87f916dcacc44e2c29ce57e38d2ee124d3154d15410e43bb697e644790b4183f6d351667b352969aa314277b00e9feed96efd030e92a46f5c2c57ec1d39cff50596a2fb8226fa639b8420d8cb956326cc6e275c557c81ec6816c14d57ecfd0fef951dc5a8481cc3c99ad7c898435724ab9cc8d39624bf69f974917732c493fe95a0d6f44312263dd79763c03e749ced1f721f15bba1886a4c8e2cf877b69c9a0f63cbd449a67469c9ea4ad9b2c8b0d475a5a66daf9434034aacaf71d93978a5496313464116059f9594f52dea2f3a26fed0eee41a298f5f48b1aeb956e18c5fbd7e7b4d61900a4bed25c65f79bff0a67297a5257bb643517426edcdce054af17099525509c4f237d7138674fd90a1a0ac0968bd7a56ad57b9e0b5b1518a9fc98c83a050cfcd289e83893c5f24bb7409ff8bcee7057ab018ac1e6578857b8a2dd6b41fcf4f92ef68d6d2938791f4752a6354b749d6089a53a23ea2b8eed48845;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h86fe82cce8002ec80ceb6db69cd4da37dd84a08d9f37a20aeac0583fc030fde8e0b20041f2420ef3f75c894896ac86ac6e650e6ce6a398f42f34273ec970cd60f746bcbe982d7bd40440d370a3e9546a9d61ea9d098a8848412c5d3bd41d935216ffb4cfef92702757cf9eb18426356e07ba35add7fe5174c51a3473490be00e0ad1b612835c629d8612e3534720ea83c7f0aa956e3d5dfb4b874068872f72130bfa488369f0d4bc02df26d0a6586c0df01ded40d5f3d9a1e13d069cc71aaec830895bedae5588a96e71267c79fd3cc8f3840c5ce4a47eb5d0ed0e11383335e45e7e0e3abbfa733e23cda2f127746ca481c508965b1c62b6a0805dbd561630f2656fe6a24f1c318c0d27143213cfa10a07883b14580c8cb2bf9b1df77bc8299f6112e01ec9b8916769baa0203bcb695e250c1a53c9bb0bbd235dda7991c78576f04a187e58bc7a84f7917d9bc77d329dc8c09b40ebd29b2b7c8ccec8c4173a6c83aeefa164ec2ca6e4d1fb0259529638148243c410c4bb88ee2fb6d5baa5058a066c9352add39d3f4a30f89855d0380e7ec2f449f6e6eede67db6994abe65466f1dfde972148a9f12bcad8e3dcf2ace94b8dc03c3042962a1ef2906c8c5ce65ac66299d6e97ab7fe28fb63fc5194436f17439c71f96f7c098dd4781316abdd840b25c05494e7c9478e16376512eec94cbb3020bf37489e581f9cd8309b3ab13d28adf7863c8f59107f19f8137068209ca044f7a50de98c5ff63811240c5267a889f8e6017348058b42bfce625f98c15189cf13817c590718df1eb76fcd6f1eb22d239c547a0c9ad5a5e6dfebf9d9769c1887e0503a424191108107995320951ce5281c7fb8f093835d0b6a32755cc1cc989a195025930a9f896ff2c2c5768eed108658c3d9a59091944d744839209f96231b1bb3fb1816809e98bb18f539d01ac6c702d88af7a224a91e9153178de25c74a0ea643c32b15963d9ceaf4eeb59e26ba96c38c1634f57191e81b877533d062550066eb956a67e41dcb11ad288aa90d29509dd6580e732efc051f5ded3ff9321744b43ad6bf9625ab7ca93899fcbb7e2be32f5afc77e7cdfb7cc4e9ae8acd2dd5e46b00b17b367a66a4cdea84ea2ed3ba8f53485813e86eceb3c06c6c002c1057520f8b53ebde72b96253c6ed6da94bc428cdeb8bf122753dd726e3f6f26371426a214f48bbdf40f85fce946eea5eb44e481a97c768e409961250ff4f1772a5646696888890ed93f3ed65981f60aa606290b276921fc12a0ec56a7c4185c69682b05f1813c8f4972f7219267860f3330de0501c50e87164a4e88bc99953b6ac94273b473e8ddca4fc9a9e04905e33d0af55b13c3b4fe0af6497acd2db064914a72f02deb21ce1594821008585a246977f862325934337e4309211b8e9ac6de0546f48620e5475f582bcacaae5b3a70;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3bd8b558272ac1055b6674563da936550ce734c424e1c80ae18432bcf416bd79ba9bcbe6b42ef95563793503b3a410932db58b2d85a51217dd53c22c72df2fe449034684037948ad563be8767c1f5fc3e7ef5afd7178f2fe14c69d14ede71314a7f86080f7e40c776027b774a86dbb88317e9724a3cb8f5223d8cd974412e2c06e28eb4cd66b85c1224a7b53256ab0e319b0da0afdc1e65ee592793eaf1ba3c84d24b24a38ceea95bdcf7e3657dcf675f655c93b672885c5f961e51f20f4cdfe8c82022b63b923f1b11ae78a5ba750930f24cde9560da94162b92dbfc62dbe4d622620c0c2e7ca156726c092372fe879a77823834659dd76e6d621c982f9847ae9e838bbcc6ea0a92858bb967c250edd75b3687ea8de041b25744396ecf1c450f056195701377c654640fd03577a1805adec405d705b790dbe33806251b38cb33b14a0f508d3c86e30eaa0b49c66fb95b872ce574fa0e61ec25509e3b1090d98f0c5e343a0ac5247dd43f499425ead6112ad760a92c356dc3fee30f34a072ceeb6381c7dbcf914a36b39c80adb064976c2d031a5c4cf32cfe715962ce7d6d337c203fcbd2dc346b13b75773160583183c5b548e7813df96c55f4b807357f88157d151bd944bd1c2ecafb0efd482e4814338a2897746d7830027cfdb863359190faa5bf419e5f3bd03b097dd7f7ce19b3d32b057e152f4ef923b7e4465ca24d7c10cbc74723223816185a35b3580b58ddc5b160b1c49a19ee5c4922a158b3fb04e30136bb113285664451bffb27cd4b3173b0d47a7bc9a46627ddfcd289504873cc668c3ac67c0e4ec33d8c960cda72fa85cc480ca81868c6268822d0110431d3f819119c6670d2d4af9ff3840cb7926ea83de2b2dc31daf6c8355384e0a36adadb031ad913e896f1625f2fe24d95e99be1b3b8e21353a84d0a985138ab5111a38d97e750956b03cd66135de0ab046262765dcf77d71b291ae2ad87179b4093f2f6111a87f564ae991453875a617c4651ea3e0521dc7cfd08cd259514ef7477b6cb1add992d66ed2569ade8a0251a35e31b8e76860ea8f8f7bff19da0265d912d6ff29aae933272189c28a68a0aa1740a635f5d224e09f7e77bab31c54950b6a84486c4fedb03bcbf4a666123e78f7309deea7b6e499cf66efdf5a40f65244b34ca687f14e50c1a2c09918acf2cb9d319e7a1288e57d9e703c7f6499e7c079b17390b0cef77e6ba07daad7dea33f10d6059d623ee1df13996f4a1fc309b4f6184a4420ca205b8133162c57b00954e486fe70eefc85d08cdf36f94b38c8b179b44909011c24e94c0d6c40e9543f88c7f31dce2e459862b5665ecd495a49a86daea1cd2c551ffabb2e44902e85950d19c0bfc1e2361545188910b4aeef5d052a81f04dbcdb6b1c2be618087444b86a260ee919fd2551f20ba516a33a73f5845349f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hafdb232d823165166c6c808c3b6a39cada6bccfc6a2d709a1276a63a1e7ef9281cb6b4e492e4dfcd6bcae4398ae9bdb86f61f0ed9df4e103a7f62418a6370752d80f1e824dc0ba9c1faa4ffb22c8d8fdf534f32be6ac4abf0c76b009bafba8d4c6998fb302ba5dc3d67a4ba067faacf9e0c01b598cbd3c312b20f093642c083bcd3f9860b371e7de9f61f4d9325f8eed94c3ca722c76c0db91b6880f2dda927939de27355622c2b355a8cbaf611af3dbea68eb6a3bd93c264bf8a71213a1a0f03075fedc2283ac0ae6c9077a045e7c0f206352cd3c3377f7d0788fcebf6ad0facf98526d289017be2c07e9bebb2ace60ec8ea5d4afa1bc6c9c6631c95c0f42517ec05d975f9cea85dab8ac8056e6ec0471288956fe09f40314a894f9802ca7ba9461d079fd8395aa290b279986392743cc62b62660e22e9c8aa7c037347aa0a4202685708193c1523e78981a3a073be107096bb972f0f90813d03dfb83fbf841cdf8c0dde53e814cfb05859b0a3b03a66ac5ac97c4ddfe97c3c9b4ac97e7850f722af6cd74720fab8777abbe309908195831aed87635abea0f322ace9c9a3c61e18e6b6e4e5d49d519aea447ada4a7b785b13682f895619ca24936c5650ce2ab9f701ba89967faf3dd1eeaf20566909e8066acc253e772fe04dac6ebe5e4f4ac9312367e8d3a8bb558f3b1fa3f3806e75a2db182facde3fa57d27560a606bf4001949f906f4a469114974a462774cc8653645b6ae321fe2bd8cfc694df46923dea8b4567a1ecabb238f927b20c267cb44a6e7168a6dd6b64a3dfaaae30052e5fb26e02b8d648de6b85ea4f66927c84c4d60988fe476f82ee2b6849561871a7f5ea49452cce399bdaf6c55c54495f8254ad63d09a8f08605c451ab095bd3c6c7b32e7aae5deb5a1e14f60c83b7b3810fdcb2178753307c7377f7f2d64b3dc18f78feec92c8acdf8e34ab2bb377273665909a879bba9f87d75a5df7e2658e474fcf3cc165df023eb0045e0be1adc80a980b8b975d55b9bab3397bb23add8f5aa92d970a026342c119c7306ca92ee9934c248ccc576ba356c593e96883bf1432eab7a7ee914820e8e72ead47f11a8744589f4a2420d30c23e9bcdfb345281d9c2133fc6ba31a3fa636c4a7d952a291e7a2021b066650be0f2398029d7a4134821e70b01318fca4741b1a2b9134cb38d792bf2a2057fe96a435517f1b0dc3f76ce77166d9b3064319681b0cafb3fc55057d908e07e016b81b151d33a42a11aa3d3c09876e8f061302da868b3e1019927aac35da558ceb2a4f052e9427f475a270a2f201d19be65a6b301bfb12b688ac84b2e832619a7356f427eb73cdf70c60ab01d40e2dfc5b10ef6cf89802c2c7076fdc52d568965d2f391ce00004cb5cbcf04333eb7f9621613d17671166781326696e83a6d50a67a0e0b601a2c08710bb12990;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9afdf80032cb71e4f132984acf3161196584fe0397a6264cf24e83de0016666382c1c342414a7ade6c9b3c31c5f140184552aff743bbfbc617450cfbf69c1395ba5d3e7124d2608386c8e17e88145684a5c884cd5ff09e67814cf488e36390898bc27bb9b83f90c67db03e4d6332863af834b350acc213ed1cef50b2a3f44724611b06dd68e8886ce3d856e726a8ad1178b31e98feaa8c72b03d6b290ceaad51bdee65e770c68bd4ec3e815df03b5daaa8372beba1c2980d17c52970ccb25847216a088f60112a2e8dfa39a4e89a945ae5a9884e095b6223951e77d84d791a5dcfc01e8bac18ce61ba8c58443c914e54e8944b9078270562f57102d3baebb85bea1d88d53d0412c9b69450df6c39f26d24e46d5f2ff6fc4933bc5afeaa2118a304d02177f9f51fdf8803855e921b220e5e7739c8e3de0499bcc8bf78c0cebe6e0cba241cc2a2df4ccd2fddb4855d89a86ec848f9ceb82cfa24fdcb26c7075015dfecb0f0a4dfe3b523c8a2c09f812c96029176c11beac272b12ea5f90d6e122139adecbd08a0e36e87ce97efe343fe8f176b7c098968fe6f36ee02e7870ca3c95ac11416b22fd708db39f3982b182263441dc8e7e5755cfef0d68e0610a68b8a7fd0636e413cddc3848a1750c30189248dd7c1070c213e702eed142c8e5411c061d8066fe44ba74d08c95b9f6985b2261260b70ca69d34d6dd732e880302914b0809c3bd29b6a9859d904d48826ef93ee1eea1d4f8fafb0e47a936d9d6d2cc0fb36ad01f3a59cf1a1077eedd20ad8906bf204301f9714cdf7f8241aa840aacdaea8ae27511461741e94af2c1067efbfec6b9f2ca6f6591674c608d78bdb8901c49944886e955b561550bc5dee8fda9c8e4f4db0aa7f978d93d09fd874ba3e550ea376f0f00907cd69ab87ef1315756ae5674f63b2dbbab54b01e69f7202775316484d6ce129e75828178be852985de8085aa64138a7ff41fa7087b117642ab217e6cd99b768a429b586e664b7c52c9f4a2eabd0381cdb3469f7e4a43b5f14292cb7fa38a8c7bd4ba5ef9bef49e3f455fb686fb50d860bddcccc204c2f42e7c9030317ab960c3996b1204c0209fa0153d6c32e71757adfbc0af307548945ecd92eec23d50a0d0e8d86189e7a82e2ef5cc8b0a5c147e30105a1e004a2d2b00276112acc035f57dcd02d35a8d950f2dcbb82cd78c777d6e81b9a6020cbacb6e2788405e2fd25c69a312412baee49557f3e6d9047c9a0abea8d181b9d1ac3363011872afb1667159d7e5c703abb6bb1ec6ad062f137fa0b689df538e450cc262c466a721dcbe21a37b4f4feb2731a2fb598f4425986260760ca0611399b42f9e28b0cb137b8fa8c34fce4f255b7654864e6ad59649984e4b887e4c46a063813006db6b794c34bc9aed90fea7fce1f4029ff835169756308206f7895b874b385d47a7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he62934b83f447171de25178ea67aebb9a854e65c9f8af105fd4c634c1d527d23188253ce8ebc5e52e05ccc8d6516beb7cc38dd1ea0d0c3f9bdb4b05ef511425bed702f1aa7fc8c8b3a3e47e1991ab74c97c456785baad8439fb7edffe29b5fb53c1761c99b4918921b5a03a42500159ff4027bc40baeb52f46a043a7557693ef27fc8e92353c1fe80f0dec1a183b020cec212905397e26de370c4df507e52acdfb77c2fdff4997366c63560622cdc5a261ff6d8be3c3e9e36ab32bd10fcc640e21f3edf0f560ae647405a067da957697af5ae45fa55dee2bab9020b44eefc42fa23f2470ccc545d1669cdcf1545839badef3bbe157668389d4dea287a7c5417544c37a8076cb450f05b5e353b694e1eb53a1046a2281130957ac87d1c2ba17d3a33a4e6d7ebf12e3081d947dfa199195a0747845cc6286c73ddf1736eacf8120e3a67024e99a591f6438335ea0bf4787480d9d2207f6cbd40aa182163175cebd547d8303b8eeac7ce4b5c4fec6957b5ada1738b845e166a2ac15386997207554149331dc9003f92c3729da8f0c954b988693b489e49275acd8ce18c3ce9f8830e459ea56ec462e0a7e176b09dbd974223f3f2ef92b0d0442563cf2c0e3291e18e94154b5ee75e71e8cdb99068f1332065ccf7ed06b0dfbabc650dfe211d652a23a9ad49e777877d512313622ed2e816b8ccdc0739a27ab3c172c65d715a32a7e3d4bf0e71a3a37f819af5b44091a71d9b976ef5203e978ff9bfe490639d13b57feb788cb6a4804c17384fe9e51a611ebb714b518c875c1ca11ed970090a187dfcd6eb676a838116fc5aeaad3c25862b833572d6053b4228994f02566d8a76c833ca421e123790992bdfb236410c9c64e2379fa1d6101439106105efe1e0953cbaefceed19cdda4d4bdfde1faca657340598ae5088d92ca050cfda2262995f0fc1081cac199820616ed09510ce9c480bf268f3c4f42c086be006909a96b7d485a366331b7f3aa05456e029ce06ecc16f12abbc18c7b83c477f7cdebe4ad66ff387d43d2431e0b195df03ff0be6b76327aaa4dbb330cd636d7692e272c37a577a45389933d69ac238f8eac7477521e4e743c2b35b78b173e0c4f55601d8360a88dfecac1e81e6d19af72ba4f87b6be9aae9dbc4429386b4475e98a4337c2a038b49fff130a32d8274c50eeed320dd4debad63fd8a4338c1853016cf9e4eb355ca6402cb2e25582b7f469db1feffc0c1cb1c3f5e2eb707306894c0534730d948b88619175d0df17004902a619ead40d90699e789eb0c80088333b24020b26d601122522fd5bc5b27494b9017d53fc8ae8f25f388709d02f2e97ead132020c6a4ea832d460fdaa9ae8d718194267a948dda64909379f408160f84869f6fcff5f79b7442bdac8c4836cc829c85c5eb9095959767af9d393231ee8832a3b9b120c110;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h97b5176d00a95a95d58808c0f62735b78f84100d9e260b4b52ce5700a228c2fe335a059e22aad5960a69cacf731376c4f94958ae0145d9939dcadefcb0edeca9793a88bd55fce97c6cb23a9a140cfc984391cdcd89c2e679f84c1b4c341e4533a1ef786cace179725ab36bfd400ab5ca52eb9e5fff8518925addb2e1e1c8543b5d501be2897dd3b79067e0dc8abd17822d80cc9f25dc5ef226c7b3a5696a7224c1668ef5eef7e89eeb81d04b49100ad102ce008175a2a6391b7ed41543a6b35682f35cb40278147e703c9317a064b7b0b2f0dd9eb0e39b9e6dac69ac2685ef62e4a15edffa366f57befc7e01016655306c49d492dcd89570ed3dc1b7ac957985821fbb23891b2356eae7b3894eb553a362f2a3731c81711882cabd24defd77a50b88363898fc21d3ea5d18137508ee726068954a2cf89a73af03d906d063675a3680f81d735a8cc0929b4a84a9ff60609ace91ac835a2f557f6b186b4374794e3fd7ed025d77f5684a1f916b4c7f0b981cde58bd7fd789953d31bb6d425dd8cf17c09c3e4496e3265ceb0acdd2e36eaba562284349363cf56bab4166addc257129bebf87afeb9bc8381a6134768689044ed1dc4abe22cd508aace996029c1cebad9e3d284d563d0b362874c74c21d7e110a4b79a55b985a08ebeabc0b783c8ebdc51adb03c5647b3a2407fab26dbab6aba0c4a089151dbdf08349aca52788868d578ace7aa71a1f4933a9ef987936edd5ffb9890a5a631e0e853df1c5fc17bb2a46f6f83579c4f8df2c65fb25fad4ef814c74eb2e21ccd06820f2f309a6e5c819e9c0a52eaf3916d0c98904f4b22e4e14cbc2033aac0f342237487ee4844251c425ca1cba51f99280eed6793482017fee52960cc144b628020f27401d86e286559e90d2e389442e8d0734f728b2216d853ec24da50c4eef0770388ffa283bdca9189ea40020f689ddbc51660c6fc53315ceae08ced28f5d4cd1c8681ae6336c7e137b9072e15e2a00f7e2f11c0e4b9ef3e1c743d8112721caad2904b5fa136e6fe30bc0b97ddd999ea8ceaf5d0cbfa0dbf492df0127c6945758d9bdf3d710ec6297ccd2cb52133f682977a448562f95f3325509affc0e07782b42f3d2489dbb50fa0b8d1acc4fc4f8a2fafed129e514f90d5b026abd295a5aea843cf70b71308f3aec4f05b3c3deba2d88a6807b59fa357ffec98c8e3ddbec4e19b299d4159ea9b2d788e9631a7b35057666b7e1d77c3c51b8f485a96f1de172c7237ddf7d5af0029b8abb1e0a8f4bbcb84242572ace1603a69c2e1b7a0f09f8bd86263ca2ab3359f7dfdd8b1a411731e71355fe2a172416e909d6be41d5a5a87e6b0fcf77bd84e140152f063dcc7db29570b6417a15b3be5a9ba13b12e62b7351e22d2bf53cd5954197cc9af75a195d4180081625f8f67766e613dac765ae3bda655452d4155;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'had0cbf77227e373fdbb4d430632ad704481a4599d5776290e48a15fee9bcccb60bb6197dd1b07af9c7abc66ae08e9efc0a8f459bc49b99e36f9fbcdaa4b5fc2dee68e0c381e40486626aeef0dc2b72c4cd7660430fa11f317e356049e9517eb795e59e995e82acdb1c7064cea571eabb6b86f2c5855478a1f148ae39aed0e97292c97310036f58c86c4d51fe4b105503af02dd6c5dd9c33d86831be8c1fd0833cf27e27cb453e4993ca322763cfe5a973cfe332d20b7fd15655ba83305a0d987cb7c0c65ce179c57bd73e91aeece0b1994abfeecd387e03b337d951f073acf62b07bf09ff3260824760ab9d8b8d8d72c5381ee70c3512320e37bfde1fff53ac1412b76abe206ebe0be57f3f9c0e3873265a03deb9b7c2975b2efbd051b32201fb9eb6c215ee0740cb9dfc6508366aa898855b1f9189ab4899d2956570c753d10d38afc39746c0f06c38f12df1ee70433eb65aa0c1bec869f339eb887705345c28507b3fa97127d73c1d701ee5b93dcc2b1a9664ae8cba9940790a00931fb3a378a316cb841e4716a22f66cdc65961de3757e98b70b09c80c6bffe6479583f65179a912f04f6f8b1baa5d637a20de987b6aedb4d9191f8186cd9edf0884b94d99effc700d2895334866a41e399f2fb8c8484721d55091923066b517446010f1e57f026cb14522bcfbf8ed11b35258be337cd904130a1dff9ec140f279c0e9f5090b69e9ad4463ca8c6b845029946a14012016058ab126b1a02432f8e5c2804c4fe6fd8b6898723fc6f8fd3f76506351f88847d019df4f5b57c61c177143131de629913e0c3082bfe3d3f54e26280d8d1d3fdc0e78c0119e7a6ea77f44621247faaf29f9937c44aafa9061ad7a2e45e3400a200e2990da12ef44cdce27f581f1be9b44989f903f0821a5e84c2df720eef9c3bb1244cb139a6d7a7199cf0ae51f12c4f3f0ea01a2278e681534df16360974fcc6b8f419328bed0c39cf105e6d30a56f3b9d91a55f2a898d0b44ced0ab6f2de529848b7f1f84df5033c76e80eb993ce993d39555f41e86216cda55911fb90563c3b1acc4508ce4ec2c227700963ac0f49bcc27cdb7befc2366c2b3d6df93898e8821b12b6122a273d157f42b91e63b60a3dcc5febb90db220ab56f126e15b0464986ba78c3a41119bb8307ace731f9eebf5b0ad24327fd614b2cdc9199a633300f7e288ec0cdf24edd09e19048491e660c42183da1b10a6281d19a600b4e6a90e9ba7a4a09c472b3caadbb75601d97e2827ecaa4094ea24e570d4d6282fabb349fc4b8712fed4e7d02726b57071942c2bc36791b41c9e9365abd40cc8827e4583e25d330c97805e43423b8717388ef03e5c3dfb107d4f161c0000c79ca8130171c4fb102b70c7e8f3b7631f42f0bb12f25a19eba09f6a26d8cd5da47699474e629cdecb40c527079cb59778f908377;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb88af78a7ed367b76444f6ef7451855726cd397b5cc93afc785501a811cac329401463a514d77164da221f48dadc5b77dea4a3be0c83ff685df689911154edaddee74073865105f49cc524d3b326165105ceb2be4b6e73f713c0c484222e30e26d7020103f6bb388f115487491ff3cbf2445dac6562f20ae3494515898effc9ac7aae9b72e54da0b4afb7cac9281ed9ef67590e97e570df149108fc919eb1461971217743bd5563a50bc29d1690f6a61857eb2dc514cae0e0c92724f161bec3a14ab2409bc4aaccb7c865e809c5ae365d5dba8dde5b399b858f8b3d6a86ca13022000672439aa117932f5edae27d5bb39707d36cf689be25ebde7d9295df6b3f1e960f87a658907b3e73d71685a26506abaa8d703f26c52bff9d0a70023b985ea5be391deb502fc33a67e38c2be6ffc2a9ce7ca16f9bbea2df6116f4fb64cdd37bb44f8f7c8a149fe96705d22c55c0b67b9225fbb45483c04fbe57e4b2f282b8fab9b4f7cfbca93d879837fd2eb7298521f32e352c9e44611c5be64a3b18336ee4971be8c2bc8ad7ff60f589f94569360ded1b1e0f0b41fe8fc56a44296b39d4daf29d9100b7ae7ce204edf9c9071e8c2dd343ff9c1468fe4008a8b2609d01f4e0b7c0250fcb93cf565240a8fa65bfa42e77dcbb16f669c9c0ac68473c39cb161e1c2a5bfddc6a91d0d45775c277eabf126a9460ea9246946e182e776e8a0b52cef3c985efee367c6a23f11b3566db3cba8ce2fd1a2f351ab4da3d4a27ed325abff6d2d74b2542b2b66a68c9383833523d3ee50c06dbdbb25aba3777618b77d140744755bfaf5335bc8cb16857193b4bbb483d2b15873d0a0cedd237238d14642a8bd3a7121ea54d9e64b32754c4ae006465fb962e9fbf203101c1b81c8b54c67d11e73a184eb65d4118365586cd7ba2f5457674a59c215c876be646e7dd0ae4bb4b120fbdb618a1284da94c049262642f1e59b5bc7627fed581613b475d0070b44cd7149ca638f8eb3fafc5c018e79624683360fa9785156f0db55978755c9c62dce407840b3440333735e4cd757f85829a26cc0de5524fc9d4ef31a1854ec1e76db39f637cfb62b221f2d1ce85cb18cc62eb0acd973de00fccf82572e49e6844fd4cd4658c746a9a37ee4dc399c89465533f7ddedac6e68f6a0604195299fb17f7da2b11fd742275d51c0464322f8c2a77dbde6331f922a53603160481fddfd04c28c27552702cc8ed5908c5474219d6b272613a1b85547bc1b7da1fcf7874013be0a44b03172e567ec4591a804f2d0ca273f5529e313610d073d9d7a1078f37d66dddd155d1dc66d4cbf70d0e5c4d9a732f3ac69c5f6bcf706f0728fb46b33ae7b5accb0e48410222dbf5681dd2c8a69f852dc23195dcf9940461aed405cc8f0c3234a48f228b3130aa125296f6a49865fd869faff57bd36cab572a4639ba;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h776f3d6ef7b04d1b0cf36b61c21f59d9bf53a355dadda8fb77da552c5b60333dea15ac92048cb1fc16588285be2b8415075a514917a6fccc70da568a51b73f704f783e07f9f63c1f5a481c7eb4459a388780cde435d9bb26d6ae5fd35817af667f0e3f4241ae00e27b4de332acaf07a4b7537f38969d40f28b5e7547c6bb47f7492a317f0702aefb68c8423486bd0ee1b65a1b4eb13dfe1bfdf55aad8fbb1a2684d002e145d20592e1760d5f14cd443ab0953da606e79f260d3d0c5ba138752ebec6f4dfd2fbf4584455c9760da0ce02f636250c3bad1fd08e351d6e4e57b98b2ae150705c4e2394dacddc2104c57d52f6c4e997ab4163181f62b9f0163e7de02906584e782e523817ab274e75caabf18ae621bb4b89a00b52dc2e6dec15975dc8bca892564dd2dfc3db9fdb833d55d13be38ad3dd0ad0e6127fa3aeb023dfd6f13d319506d1bac051717ee424af088613aa73fb609093b55cb1b04a2c85827b9d17c9a50be296ce5c2da7d0f9a8cc884960070dc71b1bef1f8c15e3bd795b79d6432e9e3f996336d25c800b6923535362d8c9bc8bc7d9b9db178be8eaa57d64169c5b3abf616f14fe9b394720f2d8d6a18b3a22bd8495bb022d7c02ab339195d6d0eaac2c74bcbe98a46671f67b194dbfc762a7de31ab396de0008e1ac858b32085c2ceecbd430f2521006a5c372f9f39d8787daf8b187b7a7ba0f8b386fd5a21acce6d6938218cdba4ce1b9c6dbd72667047db1ff2e46a13d97b60f0f2534e59825872d0f5b05ba66f4d904bb793fc2025a3fef13ffe61ea92f5f5722b1200abde797f4ea9a61c0233b5e88101de637bf2584bb357cedfd71e7c32114ae2b4f5740d1c51a257ac5051d9306b474e64df41f09405e29cd97532b0791fd5dd01bd53f7b10e58766fab42a57fab85b621e02c593471e5d855e9d764f80907eb469a56369bcd9f44dd4896b5d4e0a48e6f303ff91a3f3e962ed90992a35625124f37165f60a8b6e7a57c6541a0d54c9c4eea8c5d7352c573e44b56bad28317df98a6a53eb448176811b944513168d043657129ef5801f4794123f58fabb311b358e3c516c327e03cefb56ec0cef07b3c95976e2ca7d13a2977d4a5cee02c59b59ae1bff971e14ec00e7f4916c038c2a4dfc8385adb233e22f2b5059ffdb38ffa198a1f950140a17106ecc8f91c0104e3d545bba27fa540a206e59d8f5e6caa3b3be4fde203155b33a67cda9bbd0553317498b0411e1c33b5deff8f67b9c2ed67229f94de3b1e9e94d273bca39c6862e8024fdd87abf293eebe0d8acd28cf34b32f97ad981f990f2960de84938d7b45c09617f9f046788a4b7ba71d0b100bb88446ca9431007250395ab094089cd24401a9d183e9f1726dc2580b18aee39f45d286b96e85d8457d685d9ef88b6b396fc6cb6aea047c4452d0ad0737954720b91ef2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h157c4f27a64300261340aa8f246e68f1e338abd938a558fabd073339038cf2a98e08a8876425375b2d3682a095c219b2d91c841f76385cb4094a3761d2906513931841e4f39706fb19c6beed551d8181a5130ba2decf7472f70cfbe24620a81a27865b85de9f460aa5ba94d5128143632dc0592958f9ae5e92d310f350bbd6d1938389243e88a3acb2668cf5a24e6c6ef252daf988f04bfabfa428b7a9f038c9c78731b400b04c253bc6baaaf9b8fe454aee2c0bcab78b6ac7be7a410284cc9d98bdf38d07438af12af5d57d4093fc20ff81f617f379600038df66ae03a8247734159c47e687cb55f45a741448864a98b7ace248ffa0dfbdd3083b01b7fabfffb530c0f37c9885b783c2802ab00096aecf49c2d0b0820669a4b0c66606166c0d756eae01363e3ceb4cab289080902421421b7bc1e08bb5de43459e7f0172d833c5879d260385348ea947185ca75af688ca6d5d9a2566a8d53b6e9cf1d18de57b8e0286f005c7b6642d04a9c17df5afd22eaaffbb94bbf35c5b15020ea71fe16dc2d7e77384a9f58a91d11d2edee6ddb9a5c5243cf27c85ae3c007feffb594635e08bcff929f69c7848459ee1ec129ceb7eade2083ca3f52a672d6ed6d09d897d2781eef34f4748d9235dfaee8cf57437a8cea3cc291c0b1b3f3b4d1808e219b9d6a3dbb1efc2805e24f591c3bea445101f019f551026980646629dcfe3b1ad57d72d806cae68c16b0d610782ea79a0f0788d2d3a55f42ecf3c07be6ab5ff94ce76de9f59280a98d7769d8d89e45a12cbcad0443e87905707e2a805583ad6e5b36d2c6595e0a2a0d17f8a6d655d732eadbe2a1d9aaad3f8aa0b7e6210a125b8614aaddc3c6d57d5093841fc8215470d0ca70240cfa48f32b912671e99ecbe2581b9a96e5fe0f582acb862deeae93aea7855ad3bb3398d4cc1dcb05ae0303b204ddf130c7b13458c4ddbebe62892f91b72ba21ef8fa72d3090162a981632c793e29df513f558550f7561738b47427a9c7aa276ead2cb2c39950146c1d8e570d1e5bb0acda8579c9ee0873080d6a6e861d455057ba6991c77011db93e7b3bb4ed2b16614aff1e32f1e8471dc389b12a2ef3605a3ed19fcbd7355635685b20317dfaea0170a448aa8e24ed896ed9f8977e2369c58c6f196d4b40be4887566a1e16a8ce0e38108081b1d2dc40135441d7141350b2e34735b4a4852209c40e3da0c8542f94edbde9c10ceb8ea2664ac948d634bda3212a0a0a9957a210f4bf0638eb06eabd03d83a116dffec9b62f63976fad65a963264e392872ad247e7e7151aabbc8163ad57370eacaaffbf9ca87fa33c64e5685bb062c2f1551763b7f27d33ce7aa6920dccc5ac91642edfe414ac9f1be9a14bb3ab80ec41031655f5b0259b7a6eeafff18de339fca505440a8bd0cbeee5fd3d5a06efb76bf572faf5834e22cc7d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h589ddb02548539bf7b9105f0535864b58aced7732bc3234c46a7e7358843967794bf1f69c53dd44f1ad5e7423507b2f8dd307c20f21744e26b89677cf299fe97cd9ca8df3a79f23ed9a9a96e867e673c09f7ddbcd4d4a66d7017a50d88ba02b683baf6650e8273c76a12632d1c2d0c74e57007ab664844891bc018d1232c554f0781dfca21f8819d8948ef1c1d47d1fafb395654ea1307dc2f7344c5185c1c4aab92164aa38221ecba150cf4b6c4aeca03c8e759550553b208bf613a14d8e5337aa53d44220f0c4a056d9f8428f3c5a136c39548aeb62458daeec5435dd9b643ee7e245ecfbeb3831ea137b2bbd625ca9078c1d1bbde3e7133429b9ceb6835868de79107b96d4fcf67c2251db35e6d8fd6d6e3bfa48dcb95a79f00d30a7c889ecf967219b3a7e5d8c238d48bc2388c6bee2d6b55af721ccd8aba99591a2cb7da426c507d11ebcd03256e630996638a820f506cba4b761305faa689e3f6224dfbda5501352dfdfe02d4519d74ef0c4b08230e0ab684920c5983cf3ab176a47a02e5f6955a2801f5aad18341dce7a9b0b426151d0c576e8088238109d1922a2dac7e86510fb487779f7532713d213af233a0182de6a77248a692d92bb2c97f79fb2240759b36caa2fc1198801d7b498a72096e6a56c6e83557c9dfafa9440d57c4c751d2f73dbf240873ddb592fd025c48cc7cd0c96506c441d8d3ddcca55f8c1a3348ac16f84d29c8d9c9027dbc8b28811e81248e26dfd1a046a6914da27f6d0588629d57dbbc4479ca1c605a8d308d45bb1e1aaad2e880a1cbf742d08ea5443c3cdf503274709d9800363bcf818a9add886961157f2f74e8e781b077ad7f3eccccc86cfe7d28d985df75a63b1cbf56385e4e2b708b86c5079b6410998cba6fb806e740b79657f5fa486ce274773b22b8aba6e8cc2e44f447a5d94302f3ed41dae6b9b0d0ad7bae727f9d675495bc10fd38564f63a5683e88cd31a8068cde4b72d834d14a30bd72e6be7e0644e705698c1af2bdfc8a04f75de82d95f9e55619f8c5255875b98acdaa8fcb7418c1db2b53f5f8c01c8f837d8f679d9318f2993fbd116a8d51752e48f6d9da39e946a9cd3323b18c370fa096b5276cb7d04ca4c38a029862beb03334dcd871a32a87d8c56aab192ca8ce69016d735ab2ddfd046a025a86574cccf0956079287db8456947b7928187b56bd80d09b87d9e7d74ab04e4d5bc60e39cf93c63ae85cd94e9a505ddbca6bf4a3a581a22974597b9d1f8fe4cda67c65acb719d71c25b2468256289bc9f992a2aeed1b7e78c8fb0ad29508c90159428124fd6075ffec3c90a4c79780902072308bd85c2ac4a4d0dc6ddce3342e0c4cd53d1b90d3a78ac2a499068464ec19972838bf130977f416238608822ec60c4d603d7c37949d87c486c650501b0206dbe23fcec74448d1d7d3112aec844;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h90a32e9fa64d2cfb3cdc7dacdc4355720ad106c3fbb26dbf3c23757b3d294fce6ba2070deee71997e21dfd536a4197e942868040cd26a02099283ee0cf05a8e274a5e696cd4a1bb90571b576e5325072911b14665d17ca5bd18f103d73f9a033bcac45e0779903f75f6ddf7ff3796d8c7722b987909cb9551b579877774b5007c65f8c763b34d22b2a5a5f417f0a8bf4a1e82b09b8777c1c9b710c159058b8c271569ce3625ed7fdd3ff78336ba9a5a2ab6259a626461c14f57df6099f0828a89ac0c2b498307ab9cffd03fbcdffbfce519e68e58bdeccfe5e9dea6874e61648091e9a9c84d120bcdd2716d3d397e0c6006fc50923309a7282c37e4aa7c2fd8509393605dc55c3900b230e4d845aa3fa7c7830c82892ed5793ff17944c6b33bcad25a9ecbcc94d28beaa187c8865b11f6f4d05f1c4ecd7039bd996769840513f8b4e9b3e6983637b05f8bbc4079401f63a6272f3441c2931699fb93e3f18a5977691d17005690d7061f1666cb433f5193193b022a4eecbd9f4080d02fb9f1dfcb01afecd644783c62c2606df99afb3829bd6a687d2becbf7e59636de46bb073d1f7717acf66191fe134a781fe1dc9b141657449fdfe107a8a138cf9623300c945ac3cca4a86ed11dac2737cc8343497eb5984c0df71ee42660b771f468bf23635923d7f377ce9936b0209ffca65b34776a916092bc12abfab146218a31e0cb7aed1a28f4ac7aab67d2075aaa08b9a37bbcc2ee076fa27b9b82ee9d028f21b6a114faaacaaf80375555d7aabbd9550e1e995645ef1ec68bbae5298541a0901ab360aae6244c172505ff3d03ddac76dcb6506fa53a290d09d4738a2bf2c75a18725ee07a6386e943528bd707e6d7bfcd8239a1d15aa25859fc67871be505055afcaae03a812f8749f83aa093fb7baff0cf06733d94e3684e9b52a031a262a48d4bb5dd7db08d6479be548ce66f62f856f8a23e0f1b3303ff8da2bf03ec9f7de226385649f33cb8033874eae1e0b6bd8aafd23cff79dd96a2868c43f314727d73c1a25c842916a5ecb23cd36bbe466e2ba9ba80b62bfd1d86542e142194c8f581df58c28cbe859ac143dc42e444372cdaf57e716615cbb372dc1b121479b2b7fa47d9bf7b2f8c936e29bd7c911c4b60a130bbcf41291505152271ae4f084e9693ec859129c370d0675b7d1717ca75d7503cecbbf2d9ea5062524469dea59f7c17eb45ea2e494d4c46ff3138b0397550253d62107db35105a93ad5239618db8e71211db670197532a2e56df43da45c59a4d55c22d4e292574f955db6fe03635f1a878695d942039f98c4c88ab2a97f68cc409f486bda8f6254afe3892cca788262b27a6cf5495a397fa05c7e88578a0322f6af325f92e16f2f97ba8726fdbdc6153528aa6cf3ff22d08753f0702697bb53a771c4ae5bbabe2046bb2484b5eb0e570e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h95ce418b33068adc7682f22bbe3ab6133fa1ac40831d852f482b017742edd37b17a692eec55ed24bd0d0343da7afd8dd45f1ec91f133aed132680f35d59ed3d95a6eeae51fb3ce9b959e2f1af3b37953244b3d290a43ed484a2971dd31e7ff4997baff8f8e13b6213489966e342fab7aec7246bab0f0e9457edcced07d98670873cdee03fe1f3b4edeb23112d2584b777a97e2eaf1f2975d7e1895aa34b6f7110c5fd840c380e261b6427c78f15703bcdfe376f325201d3900e8101d9a060522ced47e649ce5d04eb0d97f66f44e07fc3db24b7921d343a276409bfbe42797e363815879cf5caa3ca27d96d5631d7bccc622361d7bd3e9d2d3ec8e0136812d5c33c020d7e0b66e644ea6c04930c410ac08b3b19fd67411e63fafc8278a14d7961d5e7156be9c73e34310535df0477dc8f2ea58af856725a136d336d914d4f38ed4abdb33d843ac1f1513fdfb77b28a5f960e1b5068ded25cf0971f47e6d3378e487d09dfff93a113ab3c62bc88175c097ed2b213afeaa60005f8b8e8804bc0ad77c1bff766549cedc71b685ca8988d87b5c9b91dc34dd848837daff20646b750a051476f61e7b7f3817141d831165b114d308d44dcda7e0abdef7df9d79650f6875581c3cd33f072e2b84e7bc8b506d84539938117139af62e114d87e4ce8a289e1ce9e8db586a14393729c1894f76270f6fa7d261694ee5433e9d5d824f717d6992734bbbacc42146dda3087c9969a92acd6ffef4a7a2d827b63e88c36b69bd2942f6a524612b0ed0a705972d000b9fa616fe97c4839ef2f792b4c98bf4bfe554affe9b98d43de2cffc308729916f4638dae83d19828ce3bf73f3a4dc22b33c04cfb827a1921912ffd84ec728c26d3d45454560ec4e4e916bba712e37e0cb54bc1be8d2a1710cfa236912a23e5d77f5d136a82873808a90e79acdd9c3d0d2992bbe0a81358cfdcdb460076f7db072626524cec78987c44cc78e6e30a95ee428caea0c134383784fb60a6ebadcb07b799aaf2367bae41b2c743f47f366054db53e25ba57f8a7d9a13209c535cbf6aeb06eb52e7e0ed8c8c488694a1288915d40bc835c2f98517789c13e0dc4232d2fc81dd3eac8a9032d86fc2cb5636b8ae28bffece982f39bfd53fbc51c99a3d26663392a7aa9700b80cdbe4af4f96e1baa86b11826f22aa3846b0eab07b35025d34422cac940d3ee8e6fd5169ecd99096ebc6fd7c1b321fa3bdef957aa0d908e2d395bedb45da580125a1d601bdd8912501a5bae8d1998098ef43074a0e6df068e506745129fea73a1c34fde7f1e3944d0511887d6550067c71d207c6ce08247e14271bcbcdc384d09a4f893fab3c72e6201599af7da93010277f59e6931fb721d0f16fe609a233eafae781923a2ac603ad2741a2b75e5133f442d5b57f0434435f0ad8386e78222e79532a171a43508f295;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h76e27c5ad3e5ebed08e80aef88fa9189391e23996c2e61a971a3a8f13939ba915cf1ed0540df0485013174a11b562f12bb5727e7bdf81c408f6f9cdd958ea2b5517ef3267c6bdcf4a4946f9c368b16d631e751c366151df3db748730f5d50dad184d9aceecb0e3a33968a90173b0452e6bbc32a95cff8586915f823ee9ed52f76a08aa17cb5a0e54054fa85ddaf828cb3a44ab902e451d4c5729a0622a1a375880b98395cff0e5ed64d3f2a32a6b36b884256a0234021c00544143ec439daa7f34014334b16d460319adf5c5df7f63088bb9379b4497340e16db97256f60a517d4e2c0c75748090c10632006b705c2773eb19666b2b90a5cea98c4efee9883f0d37984e2a68a89e4407717d6267d928b927f3d1a3a4830c24464c671b99fa6767fb8c05bdf8d572d042b2ccb7e79754f4c566c90ca46f1e419aa134403cf0b67d7730d09c2014f003a350e249ad6e2e24fc3da0db44aadff816c967f38c6b4d20c00beb4405b31f8837a817e943522b912b26d653d57f462c8134b9ebbb096ddebfba7aad96007368031e462692957880a2548b6f88787de4fe5178f60f907e55a7d18b892dfab9472370518609f55e20f682e4237e86824f33f42920dfdf00bfa815f90bc65d243c3e71626092d743b53319bb1d72a1a183ea2d03bf7d88ec4da7f5a90615ce2acbbb63cd115246a27ac7d51074ef4a926778bcada6ed6df895c0b1ace03d49bdfecf3e1e2e23455c7654df264b89b21bb360616d286da91a210765ee267ec4cc11f1c0719c97155ac328f9087d4487795c05d1005ae127bd5229d63dbcc44b70f8b573c08af9f6b085fa70d93556c486d700849357dc6e5fb755b4f6be9ee0f5bcf12ef7a55ece14a4dd43ec478c7f093c0fb6d7c69dd5077f8ade0bdc01ee801364b8e34962329bc020f9715c1e4bce9783082b2ad9c9402835522efe8d82a605a9fc5ed50fdb8e7002c0edc6bfcf6555df8b3cd43e0901a6d659dd790d2f9d85fd53b5453f8a473d9b4036d29979ec513c0f8b94d9c8a16e0277c2185886c6471bef3dff894be28988500affef4efd69b3dc9d0ceba493613c50466c5220ac03ced61968a3621bb6ced919aef5dceb58c9243bf65df920fe7b50e8db0c6ab918623aad5fa63dc847bacd24a0acbc1f8a47a3aa3388785f1427b9973c22aa9a8ce54af2408f44eb0063e2a2695b3a92ce701882483d3b1a568a81f24f02fc0dff37b58c975a4e05c481b6c088cf0fb2f9944efc601a8aeeabcd1050e0a3cd54c629de5dc3e1807fa5cf241e9627093492eaab8df2e7a8a5f9f4f735b06dc3214c0e454414e09bfebbd086d78c9aa7bca8d33547c3506cfdbe74d2d62f8cae3474c8966b0ca28a625ed22daef1f5a90187c895901ef7b2381b7a12848a849217802baf390a20ff2af606d772f4989b503b08e16db595e7fd3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb18a902d526d6d5c28eb41bc7a7261f6ecf45f3f018fbc7b6d8eec254589fb8103f86f7a0afe1822324c426dd5f21a26cacbd5ea715dd95dbbf3fbf3a3b91052b0bd5dbec7aa0d046b4729b8c09cdfee8a186982afa4a08bb214786e85f280e3cd7eb076ba0cacee85c278f98b45834da3bbe04b9232fcd6f6c3526e0792852676d990a05072415ac19c2d33d1811d219aed9f9ac578f4ef8af40a94054e1d2a7c04a15f117556d8f6bebb0c35e7598fe18f1d45599d302b3c11f16bf6fdf16f9b50234221f1178962633b3c35dab2455351c01634167cdddd008cce6b68e018878e9c9e3fc8df1fe70812b5c68827ea88372f5a6e3fcc5a153e1dd63f84315efda710b5ff78090102b9072676f64ee298891ef8c7f966c9d430bb385efb62bc8bc6a99f419a4da5e9bd4413eb013658aa2d9a2d0cf962d6ddda280813a27875aa8391492d59272fa72f5fd33dcc857a51abdf4d3bf1462b43e41e28ae09d4769bdd5ae76bff7f10bd6a7b34d4f607d7b9e1f07a46e0326a27bc1ae57374d780ad352ae6211c566722e4b0939a5ce85057c57b8ebd8ddb4dccafab83f3dcefd498e418e3480ff74f5a3ad6f44048ee9cc966f253c6be139f3665f14c8a85da9b064cb1e5c173d77a1626653e0f6334b2c64b59f325ecd7748e12074a8896db34532098db1fcd56c1f2a1137a98442d8b49ccf5bf7f2a37b1033f117665b190a02ff043fa140cf697b5e1a355e09c2ffeee3346fad5ad48d279c4f7a4abb36bf199246fd625843046d7f3d3fc0154404a01e37d4bb1a31a1c7f9ba28aa766576afee073bda63387ed520e397cc3bc16e689e4d91c46c286ac22ebf64eb671468593fdbde7652325b3f680fbc6e1b014e6fd25ee96c98c33ecdbdb334e76a4f55773835eb319e35b9230e6e60f776dabc85707c58e2bb007d2ae7198c93db0aa7ddae49eedeb6694205013964d38831a4ddcec6b0d25e22f9bbddadc5ba11e452bd71e96cd9b6b9fd91cb4aae93bb311a720bd9356520a1174a53ea48082e8a4d8bb3fb1022e315e4eb380af257d16e32c2d17bd2d5e6a2a5c3abf41a5807f0e2fc19f455f5679de3e6d3e12f2efc0c59c980ec56807bbd46d0267207df9e788e27835d3aedc6b283c483c59925b7bca7f223bd3e23a7c964f61334fd896615850630f8905875474da6cb4a4f16e592008580eb4ebda5cc930cac28392fe5ffd8c021fd169462b2ab105b0706ea567d153dd5a08694bae8a09f3802ef5dd422457b6b9de20c96ee761298a54ae70d46fb56a89f7c74244cfa624faf03d539a577d8fbff6db0128dbe985e2c9e8409734ce9f467a7b5f72240606d50f150162c483e93875d87b0d6f846583d7ec5a9e93d61e6c9c8c80723cad8a6e19bff89b2f17f8f901ee587b7dd775ab2a4d28818daf4bee3a8017222a51e0130114fba0f2d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h35aff8f31325122ac2f9e02ced4494da5f5f045d42d85d519e0dde83d9beeb97a13b96a42a41d325eb84d4c2d83494a0e59735aae139585d0b06052e691a02fef60a3848ba4c5b7e832e1efad9c052743b153ed8fb6aa27c664b7470708266b7077e1161a296c9cb5821781a87df5706736b571b2dfd2d21c911f87dafd1e460e739314eac92a6240dd4afd4059d014c9a842925c3833b4ff3fefe28a0baf0e123faeea2a879796cd04978b753aeac745744c8e4ffdd6c6683a027f6b85547956366483154ac15344c4498609088a87631a3c26f0db1b36d6e83f85d50feb5b97dc0e8641a7e38799dacd58d1592acf6d7fb4cc0b827ab4725aa9db7f238be0c5d28a00c1bfbe5de331c9a8cf26ba738620ef2c8f2ebae3fcd273e4b7247ee3cd21ad10d805ffcbe1a127a9bbc9b7c3679e8b394840242e52d56c4983c28b890c903cbece54ea89acf2243ee817fa4cc1d5d6ee3e8b3f6d87a67e2a1e191eaa946f49ca2d8187e3416073723d514afa11434922267165ea8f5f67f96e010e94fd28b4194308f0f56c6e9daf355280aff4d34c57010c306b12332d26fa506daba01b95ff9ef40dc97f3514fe279f39bc46a952e51a0002315b16c3fee2a9ccacd51173f7c2841aecc6824789dc43e545385b66ac622627f58c6e6730f72483f6c4a9b11011203ff2e9134ffdaf494577aed135bb4a20b577992481923e90395f8c4951fdd5ebef7ddc65e3ac0e33afc99a50d67a207408e22c28e1233bd1c8808bbccb980ad960f8c04c5999cb7938c2030d1a0e37bb0727fb633df25d2ddb72629cb6fb053f6e4e9248fde4590bcb109b29ca27baa2678c7b040ae20598e2bea98941bd97a3daa6159a46182bb4eb69ae32957edbd04ad67cdd515ccbc4c5a16ca9c236b9df0e2682be86481bb9f691c4c3dc6088519291913ab5556f83138beb2b19c4cd8d975d427fc118c2797f9c6c0cda39177425245581d7269ea1e1b4707e106e15653e606c758067fd3347c7b91668fba57bc060b08ef1ead06205a408b734713d3ddee07343e2d5cfed51096d79e6603c214eee8c9cc66faadd534c9415859959b30cedca354a7b6cfcbd042dd3c276c983f2d1b4239b0efb8d0de8bdc2f15c072f505848b5293c43cba851ad0439c064774c7bb5774f74f1bb50c6435ccd4b08b7f98ef020c05f92a0fb96ae12101094d10aceb4f9d27ce00f0324861e45224badcb54db9331e81c24ef6668ba2de4be7e7fe24d8ee063c5c1aad7504ea5a14bfec2e5aa19e316bd8e7c93960b0bb20f7484f089c1f9acf4f055cbbac3cb46492b185977f4869a0c594977f63af9c311bfc0f549f984c222990cbabf3094aefa865c0a3a5695ddcca3879c7712622a075be86105f07d18582910f654b35b49a0ef52ce8281ca2bb670522523565ca394b771fce4caa41d70bbed52e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd55de377deec4e816c7d2f1f98f07ae9fa359040b3fbbd658b899e577094e18b8a3a250fc8317aab26d7ab4f0f20cd137cc5a05d855871ce42794915fb6463281cf9e2a6fc4543bc82e2f54a79ef2639610a0dafb9eb8b51219f1dcd0a0c76a65693b2df9e92c47a1a017723a67018adeb55ec5f4a859b40d857a06bee83065c4444c212e616b4dadac2ea34b5b888c31bf2ed195b096b4f52d8b91303f6811500cf494b2b2d3e2628732b22ceeab39f2d0576db61983bbe04b83aa39acd39e5cec6cdd325650bb16fd6927a9940071daa800e0a5fa669cc60b65ec38fa8d5314e6410d0f92bc3c465f809f27495805f46da086288965d69c47b8219089d6f8eb90bd0877966d30c8031ab3a570817b5798b72252ba5008f03778d855b954207561a52c5585519a1a4a4db1d3801906e6467644695d2a0b92afa93c1b154b5df16d879b9ad97857c80df7f87df2927ab796dd6c187ef7d949ecd92be3b8dad692f89f4118cb7cb1522f6e9f1b92c2d130e81b3a20f26fce3e6376bbae851086561e51f9cf1d5527fa63e866ef393c51b5bb1d6d98c78d71942862ec35aa14a719b95dae28377a850f10b0fc98ffb110c35dd12ef2ccde12b131a1f9557fdc5d7368ef253148f5c24c3d0da7aff5c6aeeda251b39f77fcd7eb2133ca5b6315893a06169eb8faeaa197aab28d623c5c4c89e395cf2e2ca81bfb0c3b6296d3ec3d205339d23d683172b912449e84c8784a7610aa06b7604a6ccef7d4fe27e08d0f4d9d124deecbbd0df581648285dea66bfaf6d2da75a9580034f4d3362831164f3cfa2c4c6d4a1fbc6f1266abbe3484d14b0714a4888c9c04b03dfb845f4bae5b26ac97e052280515f22d581b6b6ebebdffa542b11e659eff3a4c3ad364323b3c94daaa30ea584031e5acb5db21000d1be25ada0375d655938a5cbc21aed9dd5f0ef8b5117340ba11da38db45a9d0be69d1b33dfb5b774cfdf444ccb5482aacbf21b403573bc8c7b8742059463b9843040b465ae48fc88c501d1107d5b3786934537b5714ffb914040d39cc401d4e84b76169b9ee485ca7daa81dbcd0f969eb3d4f305f45a896a9f9371a4291df4a00918ae6fd04baa4e28573b6eb9a65139c6951efa1f2244a7ee8dba841b96c21f988da5767d18dd1ed8c9f7966867bcd91a5f643942c4afe0f4b0715d13309c3a41dfe1b51cc55162fd66cec28043367ad1fd2e6ef207891eab1ddaddebe241d884fa2dfd5e2d69c6bc2382c4d14124d52a4822686fb501d6e2030b9593fda3027070d112ee7ac86cdd4e7023f67a3e1b5cef339c0e678fcc38c1f1706e35a44bfd4b73279cb24b8a2d8dbf59207f399e9109fce497fa9d3879b09baaa7335eabdc56b1bf618258b2b229438cc4b6d698a2631a6bd1ad2f453b4c699235cb0f0d6807d2987417926ff2c2c25d573324f43f68;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h94f93fda0d1cb093e95dc1501bffb9498e339aedd9ab43bc0a7046f56bab2292a2a4b4b83a34dd25e020add440025d96162f75278cc804d6f4a8316b43a705cbb5a107d4eb2b5caad4cbb28aad7808c98ec3b67dd2c1739f9afc1c80c1ea0fa4bf211944e850aa98f2aae636522563bd0f6a8ca4bfeb0acfc49293afc1c38ae1a044fbd18a798f5f8cc8dd3e95f67687d15020a29d2268d5e10d3cd14c6029d1a915b018fdb369e6973f116ebe2d1ced57a97adf37c63335a67b652b3492afda1b019ba16dbe697856255ba61e0b0e06f7cdda9aa329825ba1a0702e377ab00ad0daf47af09f1d81f9a692733d5ab38ec85b7d19dfbcefa3b4f0fba7a5280544d2d48abbcdef3d61a7da77ba6bed80ba413d20a3b1e52b4c293a4aedc15c098b820ba407b6fdd318c4371173ef472e674bcf2d4fbf99c1103161d8221f9c80b4d7f7ea049709fbc265ca0a4f40701a184c8ff08c1ee71b5a13059a506a7a1288b7f728b26b2eba883b78b7dc3061f2f1b480abb28b0f86ab5a6e750d4ea00f76d46519d5a3f67f431be43af3491124035e6e4bdb30df06e87595db924bdff1a344f82054af40d2a3488dbe0fd4b875c4205d755cfa6c2e3792f5f3c1df033a017326209eee8f120196968cc6a74111a8da8c1e77f456065069405a2351ceeccdca3ede2e86b98c12aecab5c4b64ae5cdfc8404026936dacc89437238a641643e0aaae15edf748ac0a220d99ad4628600f1650eaf107cc3054083b9c354d14fc4a22b2b7eb9c9eea2bf2022b970b5c59758e83aca9cec8e4d43f5e34d5f9a2018aa2af70494bc4428366a1b8a9f8d97d815791be7fedc421bbc2ccd418194004f94b74ad2a5818911ae9f3a0d43ee063f8f1ca4a43bd5f38fa23f991fe9a680ad6904843798ff56df5d347324bca52311c20b504b90c4b8a9f31444b0939f130b9aa0c71ac308d804618495a90c77613a4e2a667ddb8894d7c1d47a68e249432bf854ee0d66530c37a51ae73be2668863e09acba2dd14a8ac7bc5ee1a17d55db202d402e6c3002fd535a7bcec7119153b8c89fcbcb30b4c9803f76fab76fe76079ce08f0245a31c211c3a857240dcf9eb022c4c192cb5dd6759d21ae9325dd1f472b6081f7aeefc50598128a44a7d0ba8ff0896607524f417de001673d35e586981fbc7b75ae73038b1e9b7e4e959648dc34636ed920ecf825251ae6ef89ca84e5fb1b950c8d86943eed22a185a50df3e805d14d5668c838227b98a643d4062da2584b52623736dda499533e723e672d74e18318160639baadeea71d0d90e684cdc0b83d79cfa04f930158c21013dd7be8ca2fc5bfe79c63d91aea1eef3e5d8029e9afd0059a51ac74f155fd6fac522798f211730dcd40b511a0c8e68b268d5eeb7aecfe64d13abd9e1c96dd52b48d26e2a347a0074c2308232b74ce00b01878a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3334bcb370ad987932fa1e813c5c737ad11658df1cf5005ad64e0955f64f574007d13fcaa63777572a33014ead0573163bfe680e1ae2f7efc81b307c0b9d99e6a3d26600a26a21df2341426b967a5f4e618206c48bd10e90aa4cdd8f6d4aede879ef7e9857ec77ade30a877afc3ef42ab97fcd39fc55c3bacdfc7af48c50f17a0a2bda0543ed42d9aaad12b0e874952f88402a3128bc9f829536a4ba520c43d3c058e878807048fc99ef3ac8fb7d1a5ffef425d9178d9f5403a22570e4d4e1c2439ca96baa35aaf541b20cee6f84829ad8fce839bedd758eaf2a4c2da4808ac912c367c87aeb7251a8ba4d5ca69478d7071e31483fa5ae57216aabe8cee08707058c4450226b3823bf6bae336eb5fd525ba9a7f188ef6430a98a0f428cb7cb2c174283b7d8a7f79fe2b02d139692797273b6de2931100098dd15d92f4c84bab49539211cf63f52adbb933bee29eb95bd17ee1a213aa272b0e9867a7e997e8fa52ade311629b970d830a4d1d7127d8f9df1e7d36955444d2059f148a720746afdeb023503120c0d5f23e1a2a7be614755cde44b8ad7533bc56d84d8c7b4f91890a85fa00c5910597105c618fa03ec23a26e36656b891b9bf66a21d9ea8cc29d6fbb8eca29ee1dbdfe580ab11570c27d8db1bfa413f70400db48384eb0f1418e34b0b8979536c3293451d60b7ad630df71758c769ac65317ca0cbb16ae8dc992340c8a8e0a04b302117add05032429012e82071ea7eaaf03fc83b9861f0f4161c11e50056a72c05eab98b88a402a70c9e145528a3a71a926376f5ba1d1b32129f5322fe398104f6f1db7bccc9c4f817b3e84c8e8e6cc96b52a592c40ba6f64b67ce1c7d20f65874275de9d077b443298139e70b2677763df759fbdab419723bf51fce83fd691e518be42452a8b1757d4b7ca59f8841f4b1a11521f006d872b0b05c8eb4c71d382b248d82d6b6554a36934795864935e04493df822d6074bd8e6f7bd36803490c2d2e84d50719fc4888da2bf7d17d754686a893643e2d6cfd76fadad4738767ca8b210653cdbef15e80e8ed6f87a5002600123ccabb8b227308bcd32fbee69dbc5489a76d089f632a9d18689f588d3ef74b43780659a910a0fcbe3b0830ff3fd2b7b8f53bd7e84d5511f6b2d3e293e2d43b13873a3565762e89541d7a42ee7c8b012b20dff9092e3ed73e3d7e986453ab121db143345720014d09e0353dce4c6fa0ba41e9e6bafd7d6ef6f7378647634c4606817353afe5f76a7658cce83a46efbe761a1e05c91a300550f1665d654eddc0bf8d36f8851d5ae638fce0c92453f31e8199bc2f21b88d4af8fe48a00b384ea303bf74c5a9465c16f8434cd41fa9a2c3481ab04740eca2c122a9d987f73960385f76c1fa4e0e4845ae55558bb2de0ec75984cd65ac2183fb45908ea51a62e45e9a69a0f143cce07a5c3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9279ee1f55a4066f8c2aa75a93bab4dccbbfcd2c7729226e82e830fd409a64bb50d17cd823d25dc0d6cdaa0d947749b6462e7b6b1b3a8380d34485951700244aba4174a7c1fd92940cc8f31c3adcaccf9ead7cf06631957efa61d2ab43743f17bebdc69be24e0e3f4e7da2b45f25ad0e4f9a838eda826b5d2f81d5681f7e63f1b0111326b71b2bceab6b7474cd31544be0da54345d8fa3da4659bee074895e96046cd81d0392b047d4a496c82fc8e2051e7fbd7e8572487a766e1618fff97362510c699098c0e7203f398678b6ad6d0b3cb880e21049cfee4942601398430feaf5a04154155255def28cb1b8188d002aabdeddad191afcb2708a10a6a2b9bb8c135a738338b0b2d8c70ebb120fd20c247769b0c2d7e0e6a84bb792bb19d3c709016aad8207b71ff12c6a7b8333353d568e50039ca301d0b9a1819ec5e06bcb2799d324a8aa3f53e830c1ba1ae9b99811a4ca3de4bda80f032965ae7a75a86a06f0f41831eb07b282170454e4f582b0bd24deef3f8b981bb8afc10f71d0da1c138bc6c940242eb70f4624fa86ee6ac4fb55ef88bbd2ad468732a7be18df6407646a69064bc1c8a07097001c106baf9e065fb3ee31eb826f98aab00178802910c7e6e0d561444f55a4f02e8cdbe2f9359feb3f2aaf3a00cca1fbab03f86dedc34b20f5963eeff82ff8eebd6474040c7b1d3a241dff9f12cc28d4e4ed3d93d8c043558263e97bc4d2bab5f887bcace637fdffbf75975523a1cbdb0cd8e23bd2040a0037808b6ce22b6dddc83cfd1f944577c8749ad52e016f83e74fbc3d0312e86f16dd34cafa84fe7ff7f7f743aa0a6cc9db408906d67c7f6a610ae5d0bf708c741100c8322fe96cabb18c81926862b575998181b068851658918c3cff19bcad4b7113477c091707f782e2c5e6fef8d1fb4ea7fa892b377c673b499debfe3200e44bcfad8544501e584543630a0b0b513863f29786a9455f27c2c6ce66bcddbf10c2e1e29eb81d60a3edbf5535804707c6bcd79aca03db1aa91fb495e3a8fa828ad7ec38a19f06b6f3192bf1c148ec903383b47d5a283d705cf5730c88199551b9f7be7e2ec013dbf3e92e39be96a956383814408a3d01ca61eff7395d9052d1bbf4a9d924d2c5654bf1e59071eeeceabb7965374456f079b44f0410af08091c30b4eae31a695981343a8e1c1c09c3db748a2251ac2de8fb43c5aea3cc2785107968c1e4dd463139c92bb62f8c7f4eb75903bb67ceb8cdbd661d43cdbd2fd2d19c8c5816aea261ff96c4b3b3e1f460920d17eeea3fa8e8640252d014824bbeb989a00104d38aeb397bc6cc6de8a3d04ddfb482e0ea99afef03642e269d0f98819d557c439f0b89debd026c9c45704c309132b64816bba00c97ead4dec0721a0afdc33ad7cca92f156b2cac6b15484b8e5f968c3b290c0920d9a83580d147271527;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hbde5b098d575cf238671520d1289e21ee03d9e2cfbd52c19f4a3d7e4cc5b8304861a61abd669482ecc8fdbf388a052635ec270e0347bd10941f20af691a1bd8b78123734cafce6ad06bce78396669ea69ef2b09563cb366c41ce9a5a3ef248aafe7edabc2ff50e2da06247f635a504f3f65de14c4c1a2e0e42954b1f40924c0cf4b6d5de08382afa27adb7cd4e98733070e4d57e38d09789040de2c7c7ac6cc4528f557c1b8b875d937e5aea186b50c3b4b5d933e6f58b4cd9b910987e681d538573d39b342b66b8c3688016115018945678354c1c475da4a081f667aa5f294735617494f6f13ff4bcb165b3d6cfa5603e0253c0fdf6309e3f1ede6ffaa67ff05296e714d7ea49087cc244e34c782ccbf0aa938446cd51a9206aa8e34ef6018dc813e0307e64c1ee20c3296050cb895a2919cb3aaa7a9b300ed0ea7aa778a07bad46e74e6adf2255ac74d5f9e9d5a9cd1538e0e74ee8b8ef41b46d6a065db4057e0cd820ddb733b58bac92d69ed1230b7cb661bd21121167317682b7cb70dedef9b3e875e44830def813683c905dbc896b57cda40b66737a6b83352383d5103a9e563e8dcd5ad74c39b6f1a0d81a9f07040e25edafcd5de1b9072c1dd9fa35fc36c41a2205da2866b738e1bd1f7d055d643b65349a536d17214b80b72caa798b5bbc12cebea6b390eb74ab7905d986f21bba50d848ef9bd52aff2f414fc7ac52bcdf38333891594bbb4ba7d2b8747b4681434aec29cb2416f1dac5cf354d885805182a2a9dc32f289469b42e7291fbdc8bd88e6dd5d5f620ed4b35c9e96859490360b82615d9c2b6f8a1dfddeb49f9846bc4da9b72d591c4dc76accbf187c4529e2acccd4c4923c8ee020da2ca5a916715ea472f286807c869e39b9766f8b301532c4ed8eabc884215da63fc81f40e4ecbcc4ae2cb728fc238e6f69d2b487a475c939043eadb1f5ca67fbd1cffda347b7abb92daa58999fe751717d5f098cb49ca705937b7781c874242c0c305822215798046ee62108038579abbbc6ccd8aba6892840513ebc53fc5b9ce991ccd927124980320af12b46b9445e8a40976a5acb0ac388f52e487a59b9e7ec7d08dd71dfa080abf72c7115981b39ec4382a11deb047e715bc923015ec096e2c2c74e1fb43838bd75895a5326aa058688e5257e8b9b1253ac4376cf97ba27d8effb1ab76791b7a1c0b679dc0d4e233e0597a8944dec0a86071f6131977c4f3c746cf3c9d55fd37fb4c639cb745bc1b6d3f54e73e875a33028d41e9aba5bc2aea8fea21923408f20dbd4fbff5b853ab7e141fca1542344c40a8add2242fb371f7ebbbde10a7c9a609aef934cf320ff3f7aaf799c678ad50efa61da5f88c065e1dd66b0e5031266c1e8fab38adf4ba5d678b07d3cb95f60f7f3c99400fbf5b727538f7dec61ec829d7bc992b25f0c1f35b15963db;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3b898c415ea19e9bf6d5675bd1cdb75d175e1a755af006086c3c5a7cce77fbb78427e711c266c845a984021a216e91863940a4225126294d91eb730e3e92cf3d5221da7c34f7985dc8132c1925251469fc354ea52e628db2c418f1a94c6dbcbde907800dede4af5b466191533c11cc21f9e9411d6d1ed0c883eacd1467ce683d849adb26764c322936cde279c9a1730e3dbee128717c2f5a997e41fcd4131499117dadc4c6fd17bbaf7850789153bb539af576dfa936c201a4c3e89bfa52a22042071e8d3672be31172d817ec83886d12a14ab73519733fb1e67c4cbd26f81fe71e7dc67452a59ffb50b99bdbafbaf1ca663969fc78abeaa4ed7343cf2872cbceffec846cfc83b121244c6439d23ea2c371a93395a04e3ba0b5881e98db2de70751633156399167e02f1fe6ffa81f2a6be61d28906332c3484ca72fcd3455f87b0a0e963a7b6d519084dcbc1700f101fbcfc1c9c2042485535b3b4bb0cc214339c93610afeff147cd4dea4ff7c6b78dc467ce279d402d86e053fa9fc4418b78b3a5960a5d1f03f3f700505f2cbadbb05eb26ea895eef1f3288172a778ad24ee102e49c28deeeaf010319237b4a9f24728ed91eb710f52cb1dc9664eedefcc16ce8f62c3299da07d42e46295f718966072eefd0c7fd41929e44ee4836f5ecbb1641725f1302dab419397f8c0c3e8b74d90cabaa1b4c1916d3eeca7372e82681d9b31c8dc7a62996e755b57845095de1b4bf084507a5542b2b8ba97f8bf3fd0a216fa64f40d901800288d2cfd2fe5ab62ea467fc6627a2096d1bf70b3b6cca3041f01b18a681c444189880e3afb67bd3652e11c03cbdfecc119025c78079804c017c2e7cdb9df8553f7f8aa107d14e5c8f894654a0563f099769a8003601af54bdd3094c863b8532b19c68c14f9654d5cfc0926c570c38382e533f47b15f3b97b3e8a68bac235b2f7be7fe350fe249ab78818c027df0d0611a9fe4532c58ea69246e251523f065631963ef8381cbd062665c13c3e80353d47ba8ba86eca1c1f9d1bf4e30fd2150ccd27e03dc04276da108691beef998dd614d5d120d56e54a27c3d8f2bdb4a55ca97b043817ae598b7fc28a760d41236fedcdca22b5e4701dfa477a2df02004450a1bb157996bf8a74a3a5f6116abc3caff65f609ae9bac5eaad3209289453b885a2db48cd1dbe4492ff841b6a8fdaf586efa0a4b046ad05b494108dac72ff7c40747f27b2f8a777069d8d4105026e41b0c2d4b202eae5bcac05d0f6acbb55972e043eef49b2972d0962a445173dd0f92521c8b8b29cdbea60367234af55bb8da82546216da8ea4dfac23bf0de14d8ffe6b5a7458f876f522e220243e80e999451fb6fc2d72c1926b909d0f7d6bd6a549459d80f76f69e946dfd942ceaebb4c0a2f8b3f35d47dc4e0f443b1627a3678b6a96af97487a4de9bb03;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7e7627e6101ef7d9edf2af49f64a91d4e3bc97d88090f8e92ba73721b13774d8844d981ab61100445ca4a6d6efa76214785ef4dc0229b3a1f4fa1ab3dc72b967817d2ee8496da655892d21ba762532ba39fe3b0ad154cdc96c9e9d225f84b8fdc9b908b83ce8d80321ec1909e6460cef83180bf440b7b28048e6f1a19a212276a15b1deb84e14077291d77ac5ec081f512d7ead50460be1c1f2f1ef055b4842a8273d9b0bf421fd3d8604dbef9762bd7cf4d8062e046a060b19a2d1f5bccffbe4ada8930ac4d820798ab43ecbae73a4b6978f70a554a249c3d67e14cfa05a90a1191f5c072718aa2266376e304ef8371ea90ab9c4afd51077ba36114207809467b70dde47d0883405faf847def27b06d5a0ca77aa6d587272cfb1a352c0c74ee36877e1e06aac468b7ff4475af38547285eb9d2758d24a896ef940f4de53c2fe0aebe3c51eca4d1b212dc6ab61644e054c62c0bc07259b977561c1c9c76d77784da987caed584039582218463249437713f24df4e0b3b84d0ce09f9d8284fe36177b5b62d093deadfa5a551a48c8ec7b0a6b598611cb0338433492cca4ca4bb9d65dbf8bad9622d3673c43ef1bb2418936b1e02212f04fb86fe59d0da6f3642e8413ef64c030d7d437c9bb46bd9a4bfdfdc7c632235fffbb3d5d7aa6925bc1d285ddde6ea6dcf5299644f1de266f0fe2009ccd6cf30b8873f59eb22a516e5150612d27a6397fe2faa6b75bbbeaa8b1543f7741b07c66873d9e0044972e71051cf94454f9f132fe6a6ea9f5f2879535745de44bf5c1dca23e588b92056da710c92422ad0482e1b2e55871112dd3cb6b24286ec1075877e3c1fadbd146633ead6706ce63eef30ccd6d9cdaa01c3f50a816aef790fa7f08143c76646ec7e176c5096ea6eb3c627d65aa3ab73d1c886be64e981cfe72b18eafa16eca4ca27a9a8d8de440c09083724aab229f6aa290bdae3bc286ed743596b619f54c1b0652adb026ac2b0de1b493df2feac683d0d1a3570552aa915b9f78ca647c9bba623619a49a71fa4816c547176d2787558d4df9f5edc93d721d769c7e14c4ff40e7cf02aef1cd40a76b634faa3827b347054b5064c7fb956452f4830ed697e7a5be42ca0580b6c5a120c03ed20acc78d96272baac45462dcb510901c3676c33a0e5794dded7e480d24439fdd3e1a718d30419a94e1500a2b79115f9b046939cea0afa931a3e7912d0d647daeb2d71a5e568b52881731d21e0d784a3121eff58867935d1b6f317545006806995a230b94b47f6200c037f482a17879973cf73f0f446bb9c50d8017fd678b3733e490c411fedc63ce393edddb0395b2bb2201c1f6d128fc464528833a4636df2fecde9551a5f84f566458a48853acca2a6edc3f5bf76b7e21cff230d4a5e47d2441b4a73775c4b3185a07522557ce5ed9b686e3bd22b57d533c5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb935a0d836aec749d5492b2971e1d7c36b2d6695ffbbaa3c561a02b04bfc71024e1b4b0a0bd3e98fe04bb12842ca184852468217c711d4807591fcb71d878b1c5afbeb8c6235ed6713d3f71c4ab01ff6fc20a8471a5b56512d4fc6ad06a6372ff524dc217c19df8aff6870c7050da226551a839654dcfe5345ed1eebbdf71839d66c36bc10b1705c05325ec6c384b90a15b4c58a09dc3eeddd09758534d50b328fd5177c87b37a3dcbe958caac4cc9a256869ab8b2d465bace4ca0b88ebe63b6e8f8cd70ce65acb09e8a9c3615e8b1b4a1056fa10a5a72d97e462f885387f0becd06b965fbcd3d91adbdab903439da3a8ec92484ead21b4dfd0f39af6d3b5193b5773fc0bd281ecd6e734f90ef699fb7c2040adacb5809deaeea50e18a21a30cce83bb5d3a4febcc8b7807bc0052fc547b7ec14d80bbe2f5078e8e91f55158574d5efa6ca30bfc54a803a1a5d3f6d36d1596e01281aabbf2d7c56d663a95c3d23feb864f5ca799c2cceb0a5aa0406f4174b76b74f9c2fe91859e1ab7f8887527a2836427afa29fa3cc24e9255e9facadac12aecf87f1f8c5e1296a44b35bc6965636047944872f3cc24e6fb8f1bfa345b47fef9786af7ea7b050220761eb4bd73c0d5221f0c014c480c9cae6e2cc95fcd43b0d45dd75cb766e4f644086a2211524c9fb418c2c701f31e27953664e7096533e34dc1e1caf0b71b7cd5c7ecc55ee393819fe5ad6f716a8064545e461f6c717567148778b5a5350b6c46f3e8935e64dcbb75d67e50c1566f8a8a569da9792eecec01b1e21d396b1f1a8767b8776ad3eea9f5930ac054f10c68a61bad35b53ee1999aebb300ba5c950e3da1046e11845b4d8ef4bc290f708c779ef0988eb857357eee943e71d3c85954719e935a99e290eb036e8e9b3d601c20525c11425b1ef75af67683656bd85add47d987339e4aa7e4a06784d9ef279177a06c5c7f5b7a6db19808f56006c9c401235723fade7c056ddd40e6563774e905919bd4fa6758e28979fb565e71a3a5d1328ae1ccebed98429c653b365a0313754d61d24731c20cac1bdbde21c08418367dc88f565e662d7386c9f67e6a801ff7f87dc7b4433d3576f3408f511090b28f8ec2412d0bda0b275f1f0268bb46fc51a6fb070258c17d20ea41bd9b8ddfdf1f98904d6f0821f876a5e0cd2039e9db6fb74e8c758917e640e1adc112592b175a745f1eb964f99f5e5ec38982ff4d102b3451554dfc728f4ea7f066db9e8febc99710616741193d279096485a416d7ff25c352e7867d9ca9f715c14d68f35d699edc34b572dc82a92abab01f02977844e2f6f972e92a924c282acbc4376b264ae3c72b47991fa449842bfef872780485aa516ef72f9956740dec6c7a1c7fc44eb781acd49c131dd7918885851aecf98a33086908e6c2d1be89258a17b097073586efecadc413;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'he81f7852abb0d124586e7ca926e579ad5112ccc58aca1085ecad252c4f1028fe70e824d0b01e4d55f4ae419e203643cf38546cf4196d801dd40d083ecad77d91b10d2d50f029ffe40eb316e1b4f7699d71129e5be37c12d67ca61c821ac3f90db9beae7dd7813213d444a034ffc8f2fa60f1a9136583ed9984a8201473ceba01b0401b8c82f472c1da284a5bdda5573fce4d7245ee235bfefa913845e7f8229d0191a0ed48a34a19f44310862fcf0f278b7ed7a77825ae42ec6481dcc495099b01789906b40b918601dbeda24f8babc4faf267763979445a9aa4753a569c6960fbdb4f4a9c6aa2e4bab60d30a21e6310c6c2c17d780e8f5b810a745287a48a53885368a2108aca1463b4553ff2fbf2dd2042caa46cc069811aedf058bc587423629f9292fb2fcbc44b92bee16e003b3c6a5015945242f9b526631413dfc7a3f68f30592a850867b206e3bf61c52968f7ecb6aa989816bf053f5725c809b7e115706ee33a0c76dbe29cad7f43af310feaed22442721371bd920a07676b70491e26f9d8222fa418a0cc7b6ffd514fe10ed201a6db28bdc120f947761b9109ecc76697feaeb329a273d9f60933a8d4c25aeb2c2bcb769dca5ec448f64259a77e5553c72e937a225138bf4c2c335fd620577e07924e412322e70a47bbe298d510d82f6a2138ec92e7a221c149664d45955902bd35a2cefc0c0686499c9ee0978fc0cacbd7261e591776c1fa7aa11e4ffbba162fb7d5b2a3b041256eabf54d93cd6e6b408a41448b36fff73143400a952dcbb5b89889f7ccce83c505f0aa1ce4ef35383816e05828eba95840599e2d49cbf63c5a756644e891b5094c0d07c0b113fe775ab2aae74450aed3561caddfab2071a64c6b3c12bb1cf030165abf8209bc2085cede4eace7453ed6fd1b9fe4624d460650dfb6722f5cee984f3a330e47f204a4c7fb2674afc9371420217290ef5959d4e3001320711520e7a7a89bb101f2fdbcb7b13ba4af154a8b5a155bb87ffe7a42488741ffee8ba31e13bcc6a346f25d87fe301ed386c94e9c693edd27dad690aa257421228a2b9c5dad8c0067760b3d808961da9f40f261e0e51958c6e71f754a57f169337d761a6523c77fc8bb30bac8a688ea143a4cdf878a5121f558cebc1c9a123f5b8832e410e6b1310db8712f69d79ebec55c9d442e408ca675be3fc7a923e15dd99a6cc18fa1c6ab260fe0f58a53dc420552df26c74056723b0aad79bec7f4ac55d51266d48d4390085ff31f61e4d07fca0cf9b9dbdaf6ee6ecac7cff74e075125f8a3ae62e084c0d6b12f4cd97b86704c5f4feb3f1afd6e7be9c7cfe32c527c8d994e5335e6f51de17853cea07ad972f0c542e48ae4070e57ad416a9d5509c2d073bc43411bad6b65ac8c1974481d6b617a68bbd3945f7c92605cf2e9155a4525294024a37ffa9ca9ecffa2c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd11baf0777cd7ae571aeec7515c9da1dc837270598104d1c16f9f932091a0e08c0134d87fb8ecea6d71c18a9ce1581e13bc4c9eda805155aa67d111aa87e94cc8f281541f3b88eedd44587f34a9c991a00cc601322d04b74c53bd7784d7daf7cb8d10035f7be75a6f86d0c6a80a79e6f9eca4c96ba6eed8ecff69b1359c22d25c203b5bd15e262a007d5a91b25e8beb5a267be655dd57f67a3e726694e32abca74b1de24f7df7f7258df66121ffd85f8611d45b941cc4271aa0dd3eafda0ddd103ebc215e628d3143ccc1005b74c67a01a566d81e0b7b07a18962484e66fd8b5e0f1a7418663539bfce9a8a0d29f211b4b191e81a01ad95c4f6af7a5b3c33e5e0fb8f7eaef9c286391fae51cfe927972abcaa5e47e18f9b26fdd366d3b1dfcf558043b3f938ee32858c328dd9e130495722c4fe8e7677ca3e0707b6796bdbc2c133979eb3e70b42dfe634436b429366bf8b3f14799524c26fa6f9ff189735212f75e0f990666ebd4ccca362a3a7f3120439c526992336a790dcafc4560e587a78eb54ce36a89ffb2e3631a3eb46371ffdb74e8eba72d38b28954313099ea4e3d4b78c759059ca057f38d1ef0d33ba92ab0cc8098ad6848d66b4bfcb42a95f9bd6f3c90a690b5ce3638871517af48c16c2762909e0c52b03bd68432e269d0d21d54be1c5e9849723eabd963681bfa412b2419c410df7dec4f43466a66f04982928428897f38e38ec9db60eb0b99517939eefffd31cc6da7bbf91288ab7921d0e2d1c5fb63eebf5a9b27565e881725b92503f17c3534e7458dc1fc8814518ff40df4250e85d9988758d18e4e4cec67ab10fa2afc374f30d81d53656a8b175b051ce0f9a373b4b99026203c76c70ff093c8ea1f0759d50efa7aa142c5af4bfe8bf152327bb3e02a21a16269c1ec4df1197203ff6a318358b1d3f3e60e4d388bb8fa181db1680cda864aa9bb6a23c2c5a17d8a9fdd4ae6a79da42740cddd5d0ac56ebffbaa02660eb3bb88bb5f89709d49011fc1f456cfad2c4fa52d596c93104d0bb531a4d78a672c415884585bae70523da6d7e2148505fcac521d991468cf8cda5f5108db89c07230d92d4ae38bd3f71c1e12ff0f3cca6212a72b89277548e9bbc3fe9c496c3fc424c4d565d3504826427c5c7ea5f5ca94f02ce6083d1ff9d637e75c839b1190e43a4059e7220b695b0b55b6a4b8ded4b2951a7393f643ff6f42ad0c77b93d3d2fd1a1f980e0e168765951041bc9222cd8ac4a385b4c23dcf3b680f1ab5574de6fdc8af6b0555940b6de462c801d887de7de0702edf78bffcbc4b7ec53c02e7b053ca3dd885c9d54594a7e5704f945e03108dc1540988acf89259d3c4a41c146885f32a253fbdb3d7502c658d2041cb370e958ab2f06e8e0b74078dfee1cc954664ca4f47f5921a8c9f3041531ed5cbd7c353fb34a7d45018992;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h19b7f2661ffacd3d836af2bb1dd945b2929777b28edd9528054c2e12b062fb3ac84689e63ef2409919ed047ec174475b2bc0db01e2ec9631b76e67e26d8a97205321bd0310883e6937e14363509bdfa78374d303d22e87755759bf8eb60f2a920c2ab8e54480288ebbd4f1e6db7783d7c8c098bfd1a3e90eb0b79d85ca92ff4596f35c7c6292e8ec7b918f2f08d1473fb5fd1ca3610b6de29caf8b18cd463ee59a65e1f95423bdf16f41e9a3b642fdeab2b046c38be451a8ba8bfde377d0c3db7aa8d8e555efba30d5e14cf61ab5272f0eb523f13d92c39cf22200619b3070ddd13279d0b39fba39b0203320597f59ca9a3cc2067f5c8ba6cd2488b9fcdfcf135e56e1e3efd4c9a10f20d7491ad862358df668a8e7af60e64396f8a2e7ad746c2f3e723abbe6e8561066654ea01a6dc7d9c3e92f059dcd0c0c64d7445d5aac86feb20fb22fa64df59f20f467a0e9d6201bcf9b3bbbd08e020d48bd392a4266c5b0a2fd5567e464993f20a085adcc8e46f330ffda01b2dbb911d58e46f26d28db077bb07ef1bdae4f2662ca7898eabe32017794f2f1a794e40f64ffcae87571e1f1d0141db7b5ca318baa969e469efac68deee670dc479ea5075d9155b946c0a802c8885993194bc4e5501538e29b05c6b546279c21b085e7aaaaf575c8e62add0644e5e1fa102fd8a1881259d6eadb3c76ce8965958c58040c673ec7aff241abf201b2d5f4210facabd03e68af5a77ae9e04a495dc2c7fb8319a7f517e7e1b25162dfea7cdbd5e4c546278cb8fd07b1f8c3a9885f578772de179c7b7e66dc5629e4bc1b774828dfbf07c6156b90a080c1afc0a5c59eea5b7e5554d66efa2e45fb33924f77a8ab789ee1b56264e8d6b615f1132b95b998e23aabf6342c2490edca61ec922a3d333705ef57671ca2044ee250dd1dce5f222c731c5b4fe32ea75afe62206747c9c1711c1b2f16c2503c9727542ca21ecad35392bf0efcf6dc0ed796d3a6aae7ddd818839f7df8807eda7e69ce0b7825171503633ad0d7ddebbe24319a5200d5edfaa783884c235de055f45b2be6a65a30fb91dad3a7a650ba5f8ba9ffbb2dcfe4618b89a06abc6bd932bf9336728798a03f3a8355ce052edfdb6ba9029193097d01632578f48847b71f66154174852150fbaebcfeabbf2d5d02aecc1a7b55ce7efb095f132fcd7793824b2bd3836ef58bf6c4fe0b6a9070f769350a4ec3b40cf68e96b2a6b8e39aba06d20b283cb7ec6ec4ef86eeac431fe575ee928b28b9d601bf1bedaf38b4e80e1585ea3cb1d9354029fa6f799e067e15b379acfeed04332063aac3540884935c573fdb62ac0215c3786d28de0dbf031657858532fba2d0a9776abb34f84b261d4f9aca5c8da898df3cd7b022f5ca56554fd96dccc6658b49afc88ad6280385ec6095bd087a6f1567bf7da723e991b44ec621;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h246f94656d7846ef3c86d5c23b4a2f26d1c22545e9804d19a8c7a5817774d4aa42a2f21151d74cad367cca25c0ad7c943d095717d71bf76dcd0567b029bdabe2ffcb5abed7e6adf93025ea1b4f4b6420b34df0c9d7c9eedaa85ba07652307862df7ac63359028ff6de69235e5d7b73df06ce33334775a7eb859367e36b3d2ae881f5361c1e0b72d15eb7ce39e28e7a0331ff4830317b0048dbac227d112c30b9caa0684455cd8ca16af27c32a165210d2b67e140d99ce72c92f0639a69f36729da9bda15db6bdb1f76d05c22694be2e5a25ec995d63390278329411bce6e4eb31c0b8ef1310e71e080af51abf83c5f204e56ec45644b2573b17cc49552d88354050c3f66c9ea3da604875c776eedc966188e7334dd4455dd2f2b70682fc4eb77bf380e594c99582554e11ca4d822570990e2bf9dd028db5fb9d6446cdb16f0a1521800293ba60622776b02ebefd142e6da27e8470a0e37a6590d269a62d226fd30b6aff4f17f463471c609b4b91de57aebb48d87ef49c940faa60e5baad592bbc44f1738fbc455114e32cde00ac1791af388b8cf0bc09424dc9a185113f5d96e9fc1f08328984dd9b02816a86adb5932a6b46fba1d0e833575d27e0f404145831e922294a479024df11f42ab6040c74bb3648e5d461214fccfa92d0da93a93248e5fc29652044924e94952d21225a61756a781c4107bd04fc23ff7e036028c6d442154a5d4743ee3540387588820e2481b2a5e16455079fc6787525fdad447182a366182a33014a1aab35e154a01eccf3c122a475e85df09ea7bbc1af817040d058787a9b9f74c517210acfaf41ac508bf9d23fa34aa5be6f6463a59c1b97645c88b5b0555ef3b56ae84f8e369810b58f1aa74ff6c0ebd8dcb7a9c457969d942cbfdf0713fa96140f2f5d18e0b3399eedde5abcf18d44ef63a1024c79005330472a7e72d15bd7d0104a3680b1d0cb47ca5f2e08b1e3bd02500ce13294f6f3d3c1df99238d7028b6e9f186fb626776f02807e11cb17a777fe01159478fa82575cc54f55f744546e103c2b6f5ccfdc169171c3456a7ee5f116ad8f643b32bad5d55c0e9260c383cf4e44747060bd9343c311af6e1ddc7df841904b79f66cbe071cbfa77773b8fcd3d7b4b7114a3f93b75b2267457dfb2d946a4ffb3fad00b8d3566948f0ae6787cfad4d9e4d93f90782d0fcdf8c2c618b2cb76f08a8dc5ade1ac9a382462afcd103a2bf24f8a1dac22e3421011704f3ad446b4135072910ee76c8f569f1b64a2911b78e4a28a5d923761235c23472dee9f6fed44f8fde7873e8d067c37b538ac80580e209142bd8a7b93da90f732d555a8d80256cd2cdfaa62420c22bdd0dc9a2c2b43a4640195e31a32cb2954ad93987cde1fd065695cb3408d55d63e1899fa72620b293622b1dc7282fa99c59d5360f630cd88e5ab8c00f0d6a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h301a2339c1f8aa381f966a22b84f27d6ec0ce01b9bdc32cbc61d7622c040a73247c49105461f893a540486814124bb4e43d8377b28accc1cdd36f1e564997f546eaf631a8ec238ae98b50ff2c98c5615cf80c16a55c96a531c76fcbb79721c3e80698b60865ed7079b66d65f1fcd6e06f05eb6b14e1dde2e7fe6f8ca61b13be472945b69752bc95f7d5db882034cfe8d483b7ef028949049bdbf1df3ad34983ad0cf54e53f3b7d621c41f6ed765f28f39ff1e371c27876a199e425de9b10b293331535a779f1668a931ab4521ad4e31bc3af2254265536c2a08cd50fc58a140e765e2121de925631d27348cce4955bc70eefce358f1e05fb3417222acab8821e407a47509eb15e694d2e698e0272066bff843af4e153915328c25b9bced812cb398e8cc035f7fe098ffc94701097c317b39511ad8b83a1a02adacd1804ee470bfd6d2924214d1a1b65c073b1d5adcdfab6e81233299239e108986d6c1cd588cb3c01516e1bbae05cbe31761a0c1cfeac1afb30ea2274b5464e4469aa3e00e6725c05cfee7bdc34075bec4baf3f186d4cdbd006077b92fd09d6b7168800c5f464df1dc25bfcfc11810936197304b188f5a8c2a84706ed3efcf5aa97394b4db8cfa0dbecafce2c0df2f6044c5099b94013bdf4ee34a828d11ea0637075f42416067c66594c5037382a52e02fc31e3222948815c4bc1e597bf453001b28a6c1b953feeb3eb338e1a15ff22a0be7be8e112b956ecfb5f727d1c3c670934adcac161d3f42ef316cc2bcdcca6c9ad28c1785a5abb3e3d959084f39b66827377e9a091176fb3c751cbb77021941c4b994e0e4327582f213e8ff76601271fbd62070a0dbac33a5c0c5841ddabbd4e80555b91e788df628bd6baaaa1e41b4b296c6141f1ac6076e0ac70fac94222a7b8522cc2bc8b47b812427c187cb79ea919c240f77f3768cf605107c607468a1354c794b3b629db96776fa3bec0ff7e571bf13a53f3f515c79d774620e971694b579fb7cd9a7692ba4cbf38f01d1431694176c8b3bf2e9b59406b098e7dc5f56e0d10b8265cb1d39a8d3ed882d0809bf844cef37869ac1659c23d952d5074ede24e02150a0c7de91ac455043856ba2ee3b41f3b60f044398fd428f585f23e7eb7cfd51283a5c4f337165aa839368eabb6bcb6fa440b122e1fc1ecd86ee7aacbb5cdc06f676e09464fef924fed7310947e498cf71d5d298021dff21d22b576b8ef478545afbae744f1874576d7dbc53b96d235695a06cc5f662d05e92951d592ef709f1784cda1eddd08c71554ad25b8a41bf75f1f24420f09a76a4c4a0b094e3c2588949fc1a003fdb4858e454c56da320af707e8949f9b5b95330eeeb15f9e47e34683ebcd629a35e483c353f64c8a5bdc9f65a622af66c9f9640569b93be40349c027c62f854722bd330aa5873f31d017525dda4a7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1e64a0c060bc1a3fbf8b0854575ed53ad4996eca92d4940e07fd975e0a2e8e747ea0de0796f1b8ac7019c47e6617984d04651ef531dbe71e3636c37bdcc7ff1a895a3eac31f03c1669c0e3642bee1052a4347f4f8a841127bbd453fe6d630678442e2bee14833f561699b40b42415672c1e364a3f10a23d58b653ea9f8303e46c3626b540d3aefc59373475f24af854048e0b3c7c4520c8990c16de1743b9e05a3d657d165a5fffe154df8a8714703be74cf95d1f16543514ea38a0a425ac43085e3bd1b997b52f888374340e7445f9abaa08f2a05bfd22751e53eecdf931278d2fba086e69c56875dda94a29a1de4693c47bfaa40314fd3fd95ab914ec06ee16ffaa9507773f29c095b122c534f909544e72c36de7a3c94dc650c3a4a3ba945481e053a6759fbd3816554363e185c9e1ec9812ce0af4abab5708b870ad48374861afca62d434b5b29f9c943e80c240d6626316c594901ba32c977c0eb0138d9b720ad8f01e929221bba1195cf6ff0e650a8b0667ce3aa007b17428f06d983b1e6dcc1f6966ea4b063d1a028c768ffd4dbdf5928981f4df40101bd0419c3f1403249b0ea74b6b440fa3a76466453ccfd4806c80c20d95286f3dc2918d5cc2589e80dc92d2ae9d44a2981fbfaa85e41044505167c08380a910af5a159452336b81b3fb942e519da3268c9689279d2539bea01668ae193419ece2aa59e0b81f0bc769d1901f6c92782c82a9b30b8c6e4ff143bb89ff534e827b4db62c871f8d5c1faaa0b67145548d18f0990fbeebdeee8bf6b9607f4e84384dceecb5dbd06dc3de946f64d19d82355207d1b8422e95ef8279308a6472fcb89d4968b1d736a56d307cfa8a59a3067cbdd92a17ab68bdecd2f4662cdb331c4171507e721f7a7b065646b0a0d5d2c3264f899d8c5c05e3185424f81d5b764a887f343a734d4489e190e99505fb27bf70a5c78c314bdb21374deb0e902c792ffa60faef3cacdcadc8c18715aef687657f88aae0e82ca3a6b7c3a87f237b479c41475dab35f1acbf783ce34d752de28919545bcd3b92a4258fbaec369d59dfbce93303aed22cb9cf93ea2552dd1b7126027d7ef796f0cc6f13e7ce2baabc44731ec42b7e73106d7db94feb84adbf625a8d283c5bdfd5d91837c7abe39e837a26ca50bc7d884890ac0086e9addec84615f63b702583477063063774104f3b362f0d7e51169858636efe11d11e88da26d6779977dec12fcf672af9b493a377ee488bc01fcd31ecec34864a00e36e9e3ae4f21257a96b3a033dc4ce99f239d20c6f0e5b36a6b88e98056912a0c0e178963608c4c0993d3092ec4adb24d69c52a9b502d9be71a35b33771b52d7dda0c31b9af5f017fb054dc960a4156d08259101033741c2476b4a1a5b92979923b16cbca6607abed1be4d6af30022ca0d2435c6c4a775b0bbd0d39ae7d25;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h38678bb357a672bfc14c855ccc2b95d7c1d99ad6f6122f77ec2623c02da91f771e86abf1a832516f3a66730c5b7bf6d116581a49b2ec3b7006845fb25585e0ecd49a884cdd15adb92253480e99c384ed39f10b6496e0f9241ec4d732be991be634fed2aea3e835f424243c7e52718d1f710358e37efd1ef40e1223e5f66158b2347f2d0cb1de005ac4e9712f4812a66d4e00cbcb5495464af3e57902d778ad2eea3d13dc73d0e18d17aa8f8acca6d8110d6efc812ea66a6bdbd621f4c279454e415d4d85be63756811813fc154e9f726854e5cef07945ab4e236f3f10b9b9d65b2707437f31384b844126c1ea19993d0eef3f85c81b640f643eed86afcbacb43e3ced577ea8dd549a1f3cf49a769635dd193db787396525bf6bf6858f0bafc7e3c65bbca09d2b648cf5236dd50ba2dc50b0c47a4b002bce436304ee1a39445bbc867a850cd83224d6a804fe052eea9a041135bb24b9ebb0fb2a11c6a59f7501edc82204d3b8f68a03c91f295b9ffd215bc65754944d955fea20b6d8f104df5e2d57611513d41086364ccb95a7f78b56f34d777600386a19d9a1349791dc1fdc990e06b7db74fdb53ec50ec957ad8b86536bc4d6bd8022853cba4046230483df3a003a4fb5b2bd8b4542dc95183977d3e2215ef0bc6729e4b54fd1b51560a4bd90edb4b2a8add825ac9ce64b7df48015b9f4adc580ffbdd5b21a7dfa67904475541ed2b0cb99f644ec2bfe3a58d0e0f068dcff5d85b8a3a003b3c2c4575a43a7951bd8fec0eef301c1f071d4a9f6099e748ce36b9c74cc036b7c5cb92d293bc564a36e8729d9057a5c5c0ce91d1ccef9e5aae996fa0b2242c0da98668822008fab2d791c679fc091050ae6b8dc7e886f3fcc229a7b854fae2df6defd5115d16e7597dace8e82e7327041a46092319cbd5f6279dfb30a57faf60a81d5bf4807e2b497ed4d07d58fee96b1ecbf8ba4fcd745add295499941425e87d9961907d12317f34bbfdbfcb493a66e653a7408a9a7694535130de23835dc24084bcba3483c97f843aa53f266bfd500594901c579a703450e2fe3d36361c8908321f891e14d003b725708ea9bca37a1d9146618cee947ed9f3c10415422e01b5605726013357a97a4d844cb2ba618680104c206dcdf4f7215c26c86a4a0804b0d0a3fc4fddd3ac96d8df30d0774cceab1c3a90c901e4c72663320954db9d4c8fe50429a8848a0dffce3f86110a928e372cde22fde68fbc8e41bfbada2508bf2a61eb3c2269da471f5a52278dc8908853b17c259a0a558d388e963a20797697a34df7588fa214e7c3735a1dc9f41bb9df762b881a6ff4a1df3b3d1d82114d7474193fbcc16424e20deb91d79e280de9232d8f56ea4abc0b62b536d95d95881cbb618b3f710668800f5f14b30adf53d52b72389f4b8359d985b99f4925a722e97e53422daa997e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hab6df6efed8d6862d6b6873ab98955cdfabd614f8e870213eae73b8eddd2410066b6d27c547c0fae0da8d10856f94fc0d85b30d57d8c5d4c96b24259b65b09b2758cae62879fe3bc67a305562b26c9a5ca41f95c42236fc0134ea9d6247b2443d99a2c873a6cf25d11f65b471c61f40083521a7852a997b348cfd9b3ea9cd45f59c064e924a7c847edefb565050e70be589a74bea1642400fd3dfdf7d7339e8efb9c6b9ac0095658d7f0fa2e41e486998942f869baa995a886a1c9fc2129e338030a75bc00f04b9177b9bf30d6000557a69457384285cf50f12d8793c5b9600a7f6ce8ca78d4e60d9fca835dd08dc0d41e377a6fe3b2e20a9cbfc8791ecd6d498045c2eceaf20bcc60bd1f5283d3c122796d24125fb5b149a6ce509922542e2723e4369c106e453e6ca7702bcfe93597c328844d937dd0ad1db44b4a2783cb626fef8dec3545d6dbb701b499512849f0e8da5a32ce5cfa17fefa3fd21d317c70d403006d52d0e48553a5c710f470cf34ee1f98320e7b7875482a31824a9c4a67b53c5ed596b26a1846ee9f029b231bd3c85e315433015e23b91ce4c539b78b496e9f84202c0a8ac9ad3bc556e007da08a1fb612bd339ec363a6d03d20f0485dee6c346323938a2a5294a5c0740638e05dd0999aca1c178a59a2bdbc7f2b6aa93c2ea5128f6096388b70488e03a75b856b817ff626a453f48e6bf921973a539b88fe4fb5ccbafe2752c4d56b33a543380526413f58586231de0bfe5918bb91391025490ac9af7f5f04946ca35c007606b0c63d7e01bebca547bfc58903511d74f1508aeaea64625244a139d2dd5d608da1f1ddc726983cc5dc625e68e84f8392efe36a7f4f73cc72ad48a66b10a930f00fe1748be6663cea5c651ba768b02f3a7a80bb1010ba2f8224325aa6415ac992aff36f002eeb8b8006cb57cf0e57e1cc4b0d396112b55de685b389b33fccc2d618f56081362ce02074f7e318d3150baded430e09a37c9bbde133b7d6756f148476b093c6915f1cb50db8d9716d6ef3dc80bc1a77bf8af825c2d50f4d07ec1c7dc46a8dfad56e72de6d0ef5b1f051b06e4a8d1e18a0e4d31f320ec7c9854e8d7717060cbede63d2f3ab5e9f2ebb736132b1a411ce38d601237298fb2829624aa3fbe7a7acfe8e58e89b934f29af87b62097b4847b94d0396c7142a3ad8e7a81b3e4a49373fd60446050cb1ca2f37e44ef1e29ab8e8fe37936316f477285646d2f7159e3aa99c34d907dc76edd6f3006a37cf5456dd930a5261300a889a54b89d0b809df558f024ba6373f6d7454c584ac749947ad3ac99ae1121da45954c5a0c013217bec6e11ad0959c7a36af18e2ac4153c8c78d10a01cea2f9e540fa3ab5b96a22fa4da335efc477f86a217202b42de364fbf8fe87916b5ab7f48431b782e0a2479faeedb5540f01495bd9b0fcc3bf4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h266c1a07c8e7e8a9b55f3c9e73b58bccf60668b680551ba6e7a32678ef9c18d9f589816ff8bbf8663fdfe07ec553307be6b2d29e92bc6aaf49ae36c67fe85cbaad46b5239094752ff91e069177a663f2955ac21d6ff4c1735178a417d392450983f01ece00a3e6384049ce50611d5999fa4b035d5452130e20bd80ad7a7266ff9fe582ab5d3777fe8104844c2d514b34fc62e85cf6ed5791b592fd9ddba6cf956d3761ba8b08392e9dab58bd799b742d4816b14fbd9657a4eb2ecb5bc7c1e28b7aacfb6238e98977c5378eaa7a06f1a254ee16258f5bf12fb65c62a5d3ade1d389ffe464edf47ed46c00e46072e0c812e4b812d71f5861d4994e1f88b9a2f6050038c669e620dbbdd7b4777385fa9eea0480589fa88189f63f505cd93391fbf24f9c2627abe19b03b3afb4d4e7ca1b4d71d32566fa4f84cafe9206758114b6d7e6aa85121b8e4302aef5b1129aa50d8c7c16b3edf96ff101232b8423ac85aa904ad0ced0543b068baff6dda45069c75a15ad239cda9e9b358d2dc1982c6ae3b45c78ff250e6c70aab2476de018bd5f960cd74c2d27bdec493de453dab1e134cc9d1f5c5c9cb908a3c25403a5c5476906133d7941518f7bcdfa60653aa69d1a7fcbefdf80b90bdd639ac23b97e2d6ea6db901e2f4c392983f9d3ce612b854376eee831c1dbe4137d86a18dc4b7fd6c9571e71511102e4e1a774697457efbd137b388006aa8379f709b2bb8f5f325a31cd91ef8560e029b10ac53ad93d48aa9b17934887bf7a5fd37778886e2d5df30b73f10df44d58792e1279bc8e184ccf7752475bbbf8287c8aa0d4d9ca22465815f62bf93c05f7e62b2ca2230fb67c297f4a943b40e6baaec0251cbd1ce57360bcd4036164cfe8a6cf48c7aa0e9266884e5c62b2fae7e8262692373b869b7c577222a0b182b4b4cdde082deb3f1a5d0e4e5c356a95fa984f24524572004d778276cd09e8126fcaed7f03813663a6ff7d5a863e604f517d8995a9cc1c44a68a14dd0f84dbb2fbfe54236bc5435ae1d63866fe2dbea07b87895d2e2ba0ac7fd53d638e29f98ae59fc2b3593a4b71549718273042b53386bdb583a438f118a764823692e9da66fa695b2f9ce09e6f82377c9cc04f337182b1cab985bf58d5fc51dfbc568875ae8e1aeae03d4fbbd545ba121cb8b3d2cd1d9101ccd9de91be8fa2dc6c69bfbae204618009b31fc0b79c11b22f16d29ce55f1b9a2315f8bc5783c7ac6cb47e451acccecf0615fe489c69a4511daa31d5063c99db3fede74590919f3ca12f6b7b1709ca02b6ab72757d126fe60a7247878f49e3233cf0f464ef8996a7834d1cc67a87eaf47c53ca9657641f6b51925243a68a1484cdf7a521f37f51f183799911bb7fee2c83f84159bb1e9c7274bf767c66b5839cc29268d67d2a04432428602db2904fe9f1661b51c535756f7d10;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha9cd1e9aee59a4fd81019424630f4dea29a49b9f7b02fffae4517b65650ee040ee60e61cc4b576cea29ae7d43bbf7d20a166d5af657f35cf938e0f3095b24536d35610972e860a7fe60c4ebd2dddd3aded4d5e2799700a3e8c4e10230b17d91fe388ac3b254db1cdb4e10f06be440f9325930c7cf37f86e6e277a6f1a9ace63d0c9201ce2ef4f86ef3e6d4ecef175fac75a8af3bbb2f1013d5fcf10a32dd7ac124d4dcf1478c4e8f93e3074bcb9cb02543ef0f862f84d7aed58b33a6fde987dcef41240ee9ae5f96aaaf90c652124f97eb40dafd8ec7457fc3abdda4f9633330ebb77a3aca2f04d65cd2ffd461c4509d395eccb445fa3a6ba628aad03a69c5c713bee14455552f613646626a12a06790abd8fab085a91a6f4ee0848ff9c62f75ff18e5af80610e9fcfc59d4a93f226fed7e1e411b181d42071ebc1d195d2c2bd1a602e0c08dc33a95b8a165a737cd731c2216fd76187dc80ace1574254780a9f021e7bca993f844f3c65498e577bbe972927d56a4ce85e7fd22e04df1fae386f574a2ad1346b95dfecc754d5827e069b1bc64abfbecfd76e8a43de1d0990095446b07317279f293d6653073850d35219bc476cdca329e5848ebad7e56f59e1a88cdf704031d4dea8fd41b0d9db390ef773e53f1aa2416b59b2e02cd5daa450ef089884d9931827b2f0ba119bb87b3496347563feb861c29b22d10d014598386dc1a582b3e1f3ac7403bd61c52706941adede9dad04fde3c25f1799ca94d7c28881ddddc10a20585f530d343dc963643a3cc9725bd14bd65a08016cafa4612a51dbed3b415ebf2fde34b777cb308cd24a01a0a93247cbdae1f81bf01c56f616b0ba016dc0635377ba45720dcc03d602e0ba0c1f008c606e5aad6d4ca557ea036e6a8f0c94d522b62bdeb2083066987ac653fabf57fe0b78e264cb2edb3c74740aad8cfb2e4f62b1faf0e8e5507593e1cadb0fd827802d320c1e0c0f3fd9c0c386dba85ae449c6ccb3134bc5dc8eb3cce98928ad3824ee5481d5fec410166678c02c6ac9d365c615087d33ed03a6c26f0d06a8e56b93559c072880add5ba19b6e34d01436f3c7b50daf7120397bf98779839cc0eb8ec334ef06518529dc9215dee25a8eb9f2b3092e618dcb17082ce39ac19764235b88e744bc10d0abcc1a6c04409a3cd3171a0a54f21fff33132b529b13874f5bc87d09f0a62766ff588f7efb0479d039f735bac192f17b5aaf0fd634b8d28338ab90e4dccde0ae60f0bd19d65dfb5b048c69e32d08428773868e9f084dc9438569aecaa7a1b890cff751ec828fd276c69c9b62d7078812c7963f0509ccc99b4623f71659a755bb007644478c39f6a796c79a5766bf72c22de02c6c4b5082e137a89ede40f65e7e566ec3b3518b2a98d70dd22bb5cfb1c51500a21c7989436d56ab603266082d928425ea15909;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf177fb8e75444a11b046c65c79f18e700ef12e5d7607c31a4afd3f729bbd2cd84cdee6055e337227a833b74ed095865900ecdf5846171c35031e7be8f4a654bbf5566af26da92e31b1d60806156206b36299b669d4df974660e9fec8cc93db4df08ed4d6e18cb93bbb26dcb5622207a7abdbb03667a81fa5e041a8a61204c816c65feb2ff03c9f8e482fc5911ddbf0ab0c39d649e5db7a18fd401673872d0f5b367b92de9e9f2946669f86f3909fe71167de47bcdad8b8aaf3da2eada9b02b401ebdf8da969ece43ce0babec6b5cf320926e605fe5166d3c9492ca99aa17045d97268b640e905d69daa214a20ecba53ec6d82d56f8709f1970e8705036d7962ccc3026bcc00eff1f1a8f90858ef987cc0a8b6c8932cd5d50c472dec67854ae26d6f97cea7da573dde3c54ac036f8a20f4bb4504c9df103e0151b559e7ca9ed6d43cac43f16bdb562700e24249cb8f6f48e508d9ca4bcedd4826b3b82ad708a476c3efc8b2a039058bc7918e0b5bb077c792c12ecb434362888125510b78cbfcfa444fceb13fe85139e87c11bf8bf97a9a6a1c0c9b2fe1170f15f475d891efaaa6ed24f0448108db6eeef856ae7fdb3faf43de0b2320c1816bbe4cac3f9573d66d7ae7bcf1c8f27052a2d3ce2817db4f8d604d69ba22ad5ed3b29fd201244455c7dc7064f981d52ab86525492d20d219c53c2c4924edfb1b29708bd0ba0a858d8b592d9d569427575b5adb52f49fbd5726bfc4af2442c9b58dc2ad140c849529e0feca2b70ea3a5db570d08f4aa58805c7804f80624fa52bf016292313b5a320704ea417d33688a1fa707468134a26ea50f71be41d47050e23479640c70d65383a437f2bc250099c58e942ba8fce671f75047e5b52d2e3c32e9278ede4772a4b8a209f78b4710dc7bdcb463a34a7b7363eaba950ecfdb7ebcb4d6174345beca7db21199140d687df8077e1f1104858ca9fe11aa85b23d78bf3a25e423d93e725d96d51f1c572a6ecdb6706d777f0f4663d9a566f4c1dbc61915204a7046b34eb4820c41aa01df93c85b862cc79e1289e8c675b933f73c236c4f8795348b8b433f9433cc086f14ee71063d27f718121b500468b38b5f6e8c874412e8724638663834452c192a070646efde6c585db1857fd2ccadf900416e498befc2e726dac1d28cd92f41e9cddcaf42c8f7206db88c9223d345149dadeff3fa5b11c901c20711fc056e8af3566195a1283b4a0587e947fde83b1ed56c1d7625210c38330c9091068396e4290f2adbea16817be4079cbc1d66cfb5879d2b15525b50e1749199a2ecad6234eb7fa74efbb028a35e51c64b1c5a5bcb1030bbedcb9cde24636d9b023b7a8dbd21060b6338e6c81a303cad29227b2716bd487f649b7b1d91ff578e57295950327033359aba1297609a7af71ccff45462b74fb478e01461381d23706a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h3b72c62fa418ac75524a45894b72a49b88c072f0fe61d22237328046f874eda798adf1d762b468f0f23a6586e9e72e0cc106e9f982270477cd874b8d2810ee437bcc1eb911da6489b82c7366a9bd270f59786a0db70a59f8ea76dc113996a8090a7a1685c9c31981dfa965677424b09bfd6cb14d601582f5b2839aa8182c8b025ae2a8f753306b3d12b4f1736d3353517220c215620e3e0e7f9b99b8038fb3438044ae96f607de4b6f8c42208a9998996002a6e96ccb33dec3a11e77bff9f541f103229e25cb91aee1b5e263cece23ea77ac92cd0e6c5d692d4ea4a63714f9631cd809a714209588b9d5c2a297b8c558e7bf89720b72f7c0184a3cf1b2f8318d8d27e87c1f9cf279b1c8f22cff82f79a5140f70191a9f927fd9d06a93e7ed6c21402dce3a739b84903d5e8f0f0a08a37a22e65ab1f6170789ec99dd07d4e21707e2e56e70529409a01a1b48a614eee0d98861d243a7d26ce65b8e3c03d87094e4bf76d43e930573a16f96c2530d18d069bb59e0b7fafc90328412d515af518ffc0724f2f9279dc91610d52dd173c2cb3ab5a4f1c005165d1f847bd33c8b9cf57ac0d36dd08ce3f5edfe21eae7274f507bc9c56cecde3eb3ef0d2d6bcac21b533cb937c17ca3bf437ad92a7eedde1821f9fbf6c2b4575f524738ccf4a0896ff987808c5c883b83adae30a957526b5aaf73ac672f3ee30a17f5a0bfea9aead0f0f3761ab9a6f8ed62546eb254417e9f63f147ecf889d420d55106c3c134ca52fe3f219d3a1de2ca3d040bdab2c88b5086a744c995060cf8911d3827a4b8036f0f9c451f9e57f6dfe0230d1973f4ecacef5770b14ba1850b907d66c555a5854a50d342a1e496780c9c29e64763c4b28f68a9a4682b2d8280a3a5be33ae906ca319a94e6425c9659254e84afe7f9d2989b49ed61617df60f77284bff67cbd9c84b0f82119cc75a2b9133930689a48b7d0c16faad7af183c1658794817c30b9541e8964a8c5eee347c1523e96351224ecb8f175f80792c6fbccde9fc65cd3a94c11d0ce3b31472cff911359ca3b94f8a5769804c8f6665300fd77983c939471978d17a4b6dabc6da0face459f19d84eb4cea919e313793dc905b64f548db51af23807df758e5130f0bac57a0f287b406a785840b7e0300233f3dd5a996fa4274a3a5cd90df779afada9d27dd4c474e57a05db0275924b216e38768d91022f593d347f88ca8ef71d54edb5770bb2942c192d8ea21e929c2d0c7eafe9f0d3eccb212506e4a5817ed7f1f624e470715de805a11fc8a2257ec2331f1b4abf537d465f0e07281916026ea619946ea2a4dcb5f130e7b6bb220a1ed311f3b0171754e5d85e666b1796fde5822c18d41639aeec98de8d6b3b0fb1274dedec6527ba4537f8ed4a1100ce3c97f3357a252d3f64e3da773cb050a2c8aa0cf5e8f8ec7b882ef8a75;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd02a3b54578591da3b10a7fbcf016d9b0c3e792318d211d6e32686cda9fc382ebab4935deb84fa3ad670c75835a917207761f515074b7fb4dfcdc5ba9b71825fa6e3a6a1ea26228594f52acf83aeb9ffc22311b63f5bbb57c1e33d597f19d9caca724027f3c1e58c3a343369fe2dc03e5c4d95edf385f3046a5686b621bd3bb2b2e3f0290dbe7d7f268f2a87435a1fee0e51a42732096b500a62b3619d94e7ee547efff05dfc8e31ba03ec0992380610fc591d9ad4d82a342ab3050684b732f0171e56a4c7c526ac5c107a3abe5e3310f7ef8dc5853d91a7fcb0829ad0532d7bd0c5533c3fee5999d5602df94982144e3c61e2e031510f2ad2f6b19dd69c51d19d21fa0da083cd746a6935fa9468466631afd04dbae7187f652999728387ebd351fc3f140cb0265afb580ffd95553e46728f671c24604969ac2d859938a2b73b7d70a82400aa3b05470a149e5dd38650f4c4315d2663d1ee2edc09bd83e5bdb01f8d6180c21a42ffbb9576fefc0a1d9ef2f3ddf8a4a61ba408e9720955f5f601e3adc72bf82d02cb7fc244f7feb6c8cb5b321f3ecacfec6f941ee32e6aaf840a9fed9d37fc6f035c405b9334a98cf91c5ad5d3b33348a6b0e145f41dec307d6aed28e01b1c881eff30f7d46d6e4f43b4d0ffe290810c705e6e39cbebd53cb7a738df095730ed9fd3b93d5b4b76e30599e5bdad935db1ac2654ed66ae29b592c3519d16374c7856615d90fddda148377faccf1e106310c0c28fb7f723959cd03c8d90c923e4d676822fba68317369ad6cecebdcd966581587014430ff1fb304c106bcb1726ad3783c8bb21941b00b7d790e9a343b298deaad1c75489bbea30aaddd723b385d9b2d77ed1d17dc8c50557c3cf58754956bd3ead8bba5ea2781ad270805eb4ebed3c90a69308fdba37977b0725321158b31ed9f7b611d80b23fe28ed398e80ddf8b747d411f997d9617c60c246a4bb62621d568d90a144ac689d3a7760b1bb64cc4ca3df15fdcdcdf89c7c29694ef378f07678c46e8bc13c99ff8c49add830a166f3581c7e6813a6620c9dd9e77908971b6148e220fb9d50ed590d071a99e842de4002027f1dedd0c3e46f55c50d4407a1344a0365aa7a427361a04f30fc9ff417a1459b6d9aeab9eb384f2ada771c687c3180f343fe7d31a2fa6042c2c887fabf017bddc9ad5bc2a33747907032a320a0e87d3bb89c5cdabf7a1d2fd8f7ce6daa4779796a43d0c2b592cb9c79091ffe42d5be2a6dcbfc4f61366f9650128a0e36ab6d6e511387d5e0117d4fc9410cab26f68fd4ed2b6b44bb8f151b54b4c8d5a4ebe4d7c8a387edc4a8d91afcfbf141dfc51543885d5748bd18c26902cf427ee01f3cf40f711465a3569d6c33fa1ae3e5ad1d493f3cbf0a79e83425731a926fc3045e20eeeccf1a0122b568e2c9952c1319cee716d37012177b013;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'haeb6407d547704828c735cd87b8b8b7b94d09ea93f2c67bf096fb193521fc13687936a9eac42c0538b5d32ba76f08c0ddd9566efbfbba490495fd38ba8b354198c2be5cdaa0ac17a5b36e5cb62a654920ba939d1e3ed44a4520b03a6e2cafb6d6e158e9efe464998536ccdda0d5f72cf1797c7d8816fa8ec4f4b1159d0a4e4516e823bdb514527bc337e236ed189f2f55d8e7d76140b3b1ed83eba7051d3d1c8e40e4dd63342a0703dbb86eb7c2170308470f388b1e67f61f24c5228a7b36f1ab1b06e0cf9d90cc09d07c378290c9308da3f0df75d00af87926dfda2782160748195fa5d38e9a674a2903e229ff055b5e138b6bea809b6b7ef24562d3939a9ef740fcecaeacd7b5153205ea21900606921b242236dbab20992bde18091af80bdd60169993c9d4ec8f1139d43a6cd1fbcdd6bf2340168d90c9473208d97eb144074fd72196151515717fe14e4469735b0b593b36ccb216e95cb08d54b5b4b315784feb323e1c973bb25646608ff025ea1990dbbaf750d1c8ffa1ed81345272b4373ebeec751b0fe2e164b386276a2c26d3d710d085682acbf22c29863af051afc3bf10297cedb90b1f0f7d9b7eb7b5c904825132fbedec9919c6e2b08dfde2998bb7c4b95dddd61e8d2ad106af9a9c7cf48d4386ab25dd4d052fc2576ce2af07a24bc83ab674e62cc4149b9277cdc5cc7637a340f838aea94a1f2b12615f031040820518bacdbd8573e02d381dbee8846aa1a15c43917a50e17a05c7add391a6d26c72878009d515f098e8cade87b7dc1f5e51199b9ae32c24a8f4b6083e107a9782cdddccee763c74bfc1a16eb9f1c8609d77bcee4064eb6bdd0561c239e90715f38b1d945ece924047987f44326419b4d44b192251878ece1a16f2c0b2db6c28aa3f28e391ccc08d0eaaa363175d401eb3a4445888104cfdde0c2878205a59af9a14469846d3b8e2e208fe3d1927bf8431f5b00416031aba5fbf18f3906c50221d5847927ffba991a8d3e475e66355f9a6b317d4c611d70295ed8bbf9c2ea2c2f375c5a6b00b8b33dacf88d3dd5a046ad49aad1a48fa1d20158a09cbe5e7fc2caeabab03e95178b91a3d95e0dc2b435e2df6727e84eef71c6183bb1f5adba78f23e8fa514fa28ae7ac7a32508f8753dd341e0e031c9cb6cb5b27104e15ba3ca75696a1326246c966675edb06351bdbeb6c6c109c4962c6aec7a2e093baec7b9be9774c83d233344cdfc7966298f1c2573c448cb9961ccce650c7615f8f9e0b6cc7dada003178f9ef44e49d2e707168c601bb55b6afef0ad05a23225d05954d67057f5417fe8d7ac23cfd6e84af8e201b3291a997b429bf5ad6b295c4c3896a4b310eea24514abefd099de061269623ebb391b646340e22504255261b37b72ff1f3f245535e04d6b709753db8a2921b3d9cccd27245e132d02e7146481e926b4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h54519c9b6625db05fcbedcb7991559bc964f6fbfee5e06b54c4fb28cb713db77a478e2c3075cdfaacbf46c17aaac0356f480bed2cf627c3a80ecd1abf42422627e13081c6b37e15a8f198020a369271df8d82386f74b11d2fd45dc1cc63703cd6299314e5e9ab14f4b91b2f039a86745dd63c2c0ccca22d712e89084cf54d47acf36fe443ac8ff2b8fa1b45afe28bdf6fe31fe0cd138c5465847612cb2005f7ddcbe1d3f667a7a516efd472846a75721e9aa911f5bba37f84da439472b8e039baac586a52b5c283f9462f4011264a9a1481709082cbe45d611928661938db652571774b8d8d6c279547023e7a03bcac967fa2e74cc7792d2f35899bbe0ee5d716eae278d587a3b3b564f96f57d92c40da8e70e031b9f3f6c45b4be8543695480199cdeca0758568a50ce82955393236f4e714c35524dfe371b29961dd2c264442add8b4c8d804da8d71fc060a5312b839f337af86b8a612ab5678379a54a82982bc156f49a52030906a424726d2cad4f632c9eab2256cc8548ac511de8196b4f8c0e35294e7d8c4a469be028d08748e3168f7b9aab9a817f986302570c683480cf5169ba00d5fb9ff77f02f213c5755f47c9aeea0d3547c6003e50faa2ded185f8542af7503bb8af3e36d084e3df14e19ee25fcd0061ee88798bdc769ae70856148b8de2864d940d8ff32853c9ce8183c7312c56c5d506fed799485b23d67a5c0169a2fe4f320dd6e911614570bde0ad71155589b1ab81322d8d1a2ea8866d0945107ef6621199cbacdb5ca7d3e15d35cea6c7b03e5b5e2691050e0116c54522d3edf042cee41dc1be079a4bf3d9d2cae75d5e712df2e1ac1414f16e6a4f8dc4ceeeb2088390e16ac655ee0d31d14c98e738167cf3ac101ba9331f28abae36e911c199f0e51c3d057b88ce3ad443235fbce55f27fe3c9788f91db4d405600395dada0d31f31f2c8160eaf0b1205b4517cb61ba31f8c996b228f6f0ef3b177acedeb23dda236c582102fee9667bcae56d2d6eedcc6af55f513dd216f226960d889a428072fcfa8f8cb4dc9e30fdef4b9d6376d86e5a6808b5a8829f28a57bb00b6093450c771e875cb839463c5ee7b989b78d8e18d7a2e50d423e99fc2a850ee0e96c2c8a052509a1f9fb7dd2ededf217cb95bccc79834aa9d45d77d5a90ea1cb3c8db4853c68e023b566eea00bcb44a369a3998e5f1b5d0b8198a3ef8c3e62cba457c7049f27f3b5d672718b4ac57245ad55d0278c0b5dd9107199f72fcdeb33faedd5b07589de3ec7387a6481bbedb29c0dc5e40427a58bcd3218d527255bc3eb21adc893a8d59cac3bbb2142e16343869540bfa3adf8d043e56196c1f4cef2a8e3967e213975c9d6656462f72b10cf67d85bf53f1c1a2b34f591a0b7ca82390bcf74735255f8a6c5b17098021b23a41668a6f44350e79027cadcfa30ab7417;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1cc122ef62bf9202b8a532404518b81540a75a2dca917da5b453d64563e8f4874d37913cfca50e2f3998d3e70c6ea7d2862aab2015df3c7f018392a64d31634569b51c6ac29a82f52c16de957076ab4bf657e2e31436a8b7916bd206d0a2f6b71f42be4f88231ea6ab5d145164ecf7b93f830e68c6e6a818837dad4d67846b11399fedfa7330f6b7a60514bd3f5f420b2465e564717a6a67690fb854795badb85b1b361f7fbbad4387b96b35c8019a41faa837ff06d10b8368794120a56a7c7a6c8970d87778c1852f012e45422d621b51b0a354276b5c82a0c50e422ea4cc2a63ff62736855f4d92a6ca63460d4d6baad55d4338d805f16f4b049a2b2e50d81228946b6f158df0a691725d718262f9f810bc8c9a1e3f51a41eed6e9f94fb27dc9e04baca53a8e80f6cb93144b89676fd7f194c218ef7022c8984623ce21f6fec4a827857b5b019ca3cd5cb3e8ff8a6dc71836da696fb3a68d8cd91a0d0b64e67bd0d382d2912e9254540821ffcc36b1663c7edc6c41730dc0f39dcbc3976366cb6ee634951d60e3ede9670e26ca6fd1b5cbc0a86eb1ce1d55c8c617d852a5aaffe10bf9f47c11f711233ef88fdbdcb0f87b76aec66d6f42ded804f81f0ca7721b44ebcf78acd8505b1a1d4e4fa067cf81b269273606847c8d57ef257d7962ac8a610c1f20cf4265670cab4e357b6ed4e1f1f5cfe1df005505835ca0f20473de7b80ac2b5d39da92a5e2ee53f1a7a1d078b634752f742bbf3a785d983f7b2a57d9e81c2fc07b30ba6108107eec12fa89ca199ec2550dfea449490d991110930196efd41134c401ef5efd2473cfc0709427945d268f4e8ccf46372386e3a4ed647d996036947fa1631360464845304a4684a9be73125034cd605da2c5748908165969553fe5e652e9dd36e433039bf2365dccdd776d8470ae6afa98710a355b479292ad664d8f01619f8d8f379c421ec04e54c0e4d782bdcd6a34961740ab223ac71299abcc89b6096b9b45f1b901087af0cb42de78acb3c9a63889130b4c304f2e55117b066b286a6e2b1dcba76cedc53f545831e040145214bce72afa8f574d1fefcdb3475ac85136665087e075936806644f28ad41de943b0c25b8b56a06e2356132c7c47f8233ba9c67cd56d1ec481494a025e75d1bf601bea1b720b463bf92d1ce723edefe158bfe7de14d188b1dbfc0a1c63f4eb74f54207c81d01eaa18f92052fd663f77a29b2e9019c479c3b3a84861e87f04b426d318c90846191e9322301f029dd5d522ccaa327fbd648a73f1c98f9f04b3c77e890237921f2766e08f1bbc13fbc506176f1de462f6908819b999071682ea65ac077b1496697c7a738d19e2f3bd3298a78939e6694c4a38e02a5518a5088340b594d0cb7fbf93ad1e6ad466fb98ecf5f081aaa5b1e503c448c746f7f7042726067950636d53d9ef99;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hd74e301b81da3b06d989687d79a7b541791f80f35e2d73b549afdbb26d972c0aa57ef97c4ceb999e55157fac607c117f6913b1c2123ecc65e23e3d1ee0022af4c9b43fcb1b42d58586a84eb698d31d7ba2b3e128a753ed76f1fe3a585f48e9c67429fab83fa302382319e413389b3a10d347056dcaf07192f51f1f488f45c94bb6d80bf78b527bd3b316250071617b5c294004ea649950cfd630ef8b8a51a8a738eef5231cdba635914cc245debf70d81cc83f9180c980ff406b512d7a26682709eebbfccfc1c4ac5d23c60935bc5c701aa49c7eea36547b2ca2b0da586f19769414e42b7527126dcf5a0b685ad6b3025e9d12ad5f2ca6ac13d8e8ec055af9cd0f43a39654e19a08b50a48d047fe2e2046439b238aa9d0aa35bdedc34dd0278adf6a26b931db62b1a0944b029590f42b0cb564bb87e5923b64c757b33828286dc6907f3adc6d36da7743fa80154e5285883319ff9cc9ed5182f5fbae2c54ef1fd1d95089f1dfdeb02112bf71eec2b7bb79fd3c17b5a83427c28be65d3b13df84bd0f2638949cf04947e0fab6fabee90b8940bd4f6f6d213093b8127012a4eba915b4d266f1302a3542c68cc9134f60602550b2ba8a9898e814d49498a012cd1a51f2698a4c8973b380054cc735db8c8ca175146acfcb5e82caf92e18873125823c4f26a554a7bb16c2a7f03b1919d98b016e5801a24744b4b13b93676f107a2460b14665b3bbd2fc88ea060a9dd25e2b3194c69f61eadc2f07b6e5b104991ca7b3a1a5829be0ad0ece99c424d6f3ea8a24f2f31e8c7b839cf2a5033c16fbd3e133329a7db7b78b687afb53111c150dec8e038b23b3fa9af713d909efb38864e9454608aa881f0885a0adfdabbb7cac7e02634dd2aa2687d4a5d9cdd615d9ae1968dc87e06820657961042101fde0ae233ab2c60d8b1dd09463e513fdafe011009bb045a17cdfce69c0ccb06f0ecb3943bc2f985f78468d2d953e057538e601302262bb30061397d7ae68691e0e7dbfbfdd5a2aa367304a4a5e82e6d22ba1bde90091004a2791b2973c8e34502085a1faddeb07dc7abebcff1427e73321a469cf5f94cae7624632a7a202237b081d57bbe4c5bada56f4f938df8d604ae838182a13daa3400dc127bbf7e9aa73ddc9f413c0f2bd4da0461226118972e61c6ea8a429ecc9009e51ab36dc67dc1a74f6a9845e96e01e1d57b75dd81ca7921211438e002a3287db0bc4ba362ebad942d01e3a97a7db824b1bc99d3993b0b1757d7aafc512bbee725d84358ce25f4d65d2c7aa30fb7a5db391dc5e0ba4fd1ffdc0ba188bab4d01552f210d41edd42f30d43c266f92a86b55dd918b31c0be78e36194c3dbde1cb02623e1c80d7e09d30faae4b7fd1c25a57004082935be7792f5ae572853b88cc66404e8c52d6b7a0507a8e6ef0af1f20cd7908cb4b95e1f8322f9a608;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'heeecb33ad7fee15c1d216ec1f22d76af964a35a2aa12599fd0377d7ad6797a4511cb07c82d8d3c62d578ad92b0654eeffc1986fb33547b527f230c042891b8846a7a003bd1331658728288cdfd5ca546b36c538f292f597065dea7b8d87f4f864e688803ea2c0d73686c73f74938863bff631ced6ee3d62980d6047b9d622e43adcb0c17f5614955e53148536b92ee8fe62d16f426d8d63f1610785c1451b5112b1d72a0b7284826bad0aeb42573ff57c8333dea7b96095963e1ad12f72855731e9c44d7143402e2fcf2312267e605a9c33cb2694b2ed8e08df7dceed3765d0f0a375f3638b0bff43937e394fa6b49d51218af08d09c3fd7a3d8b31607544d2a1e64630a13250100c791a256c1eb1464af9b8efdc853726cad2a4fcf088af01e1940ce3790a6365053531039200fc9709e7f5b1939341eca24ba026f2d4aaefcf841e9f05a5cc283c2086722ea7ba14cbad4b844628b7cc0ea8e863e662b3db6abf399a0e00ef4c91401ac9f69fb7116f1d995b35fd94611acb3dfddf783a0505bbcca2d4d22dd32787fc5e56815f9af551ae5bb2bf8540ff7985468ff541b89ce33fcac692d6ac9e34535884cd54ea40a53d24058f48afac5225a894cb09ed9c01d0e2ddc896f934e20cab1843f54620d7214a4d80b72abcb9c994490a5931139bf4ef36c203c23f279136b37355b634585b7241c11b59f7d4201b551c9dcedd8d76f39fa1ce6cecf70409c8ff4b48cb8e91b91bccedea96af87185cd89754a0432397e23d2feebd9daa52c38a19bc19a6d5b5a9d0bd471a3563eee9244fbdad0507fdc5de21117546d7812b9f03c7ee00b96682e3c4126475f3240aa791ff52711d8389f4b486842bede8082fb354e32c1d7b3032c247aa9c4c0f00923333ffba150f8f9fdaa4e0f0f4ac8f0f7354dac2802752de813c9e4b1374c836be5a600d1968ff6d68305e679f0b7974f1da9d9cd9310f6199216212876efc8cb9c5d195ae3b6273661b4f6e02666b549d3e62285fa9ce43fe0807c7d0db0f2436512c8ee6b9954160767c4a0faa959a7b25ebd883a3b2c7fed3807920e27ce0d876986b875802afafcc79b686e733db7d352b1f7dab9b5b69d6218c3e95bc2f6b9db2912ac17550a412f0c85c577e066b6598ad33033316a4ae80b4b5f5a5f07188c7c50eabff937431f9aa8c17bc931d0f8abd3bfff06eb86c91928d61f49c44a320571109382182dd2e0e0cfab8c3f8618c4f5a9a7a24913311c6f2598a1e814edac4e9b77086e32726cb7bafbd6ec0616774c541e89a317f910f87d158aefb83fb1253a96d131bba16a6a012449d8dd3b6790d4dde03db7f37c3eeb7ae0a1317e1cd328b5da7ef416e93722f4c057be21f850c2e0f4cffb3117dcd643f1ffd0c51c3e5f61d41cdc1ddd359ab134054b606dde91c566e677980a4463c79befac9c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h9563b38239023763a8654b55e6fa76b6667ee01a8e6524a20667ba1a69492f3ba5aa8afb834434f80546c869ee32a1af9b3ff563fa6d5aea5181d93ca10c0edea5ef0d12eafefbc0b3c3f791d0c009a12d092327d43a5ee84dc28cd915bcd4fa15ed4ded68e1e5d5a98af601764c55d3b0485f6ac82880c5a66a03000c75a22fd5ccac3bcdc7769692daea6921073c42d66daeee9bff8633fa7c75588fd91d2f553df6c7370858b1779fa0dfbe11083ea1d68e786358f5ff085b84ea7cd8cb07042eb68837b04dadf7643bb3770655d1a6c0d4873068ec6a0de4a48d0a788c3f4019614a4cc143c79432f20ce8ad62152ed3479c9fbeae93af008d9d48dbe8915120b480ebc9d204355b90a45e79f9c3637a4fa65144a4167601b3f7702a2a5c15be18657ccecd014d44723ef097b22e935f304409b90baec30726d57030aa3084096a34b501cc8dc6183f3ae8010b63601bff0e040ee4a5d0837b0cda05cb258e5eb94cf795a93eae05981df7ac08409ac7eabda3373aff5ca0ea4bf07dd66737fa7bde3b9965f30a6bbd9ef2c161b51bc759ec74ccaf07d7287ef85539302a7dcf16d3bf04e338a22fb708608810a3588bf85f95b18febe3c51c9f806d33fad96bf89799aaa2db734e45da92d82d01ab65a7dc1d4af55dbb42122afebb70957c12b70fce6e5a88ca86549944697a8103e57fab64dfa6e45a8af6a9852af737188c22a7d1425bb78043f7696e53b4cf4ba44a0e04cfd46042d40c324dd956055f47189cad2283aee646eca4499d1ffdaeb69cc77dc05feac777c87c03f58c143a510a4cff25274e29ce3219d9e846da5806afc48aee8cdcacf7ddd56bda1db4382650b7677788b34095eac1555d39fb2cf23de8c4d220a8db9e942240345f2998b738b83c9144d118661e183fc9b365a5ec35ca50afeaa38d2ac0b914932859cc0612600b6cad6faff26d5af287ab1d00300f380ea66b35b3120c864b499635c08368a4fa0928107b7cc7b5204d928b37059ad843876c772183df4b07d468e8af3cfbd7f7ca3f5ef12cc6ca185882d095e54bd4ed7fda3ece9c39539cc757605f442f30185f72f53c43c670e35297bef093fb390c2649d1eb707fe5e27bce2f2585d7d4d1f927e15cf31da6801bac9777eb2a50137db99f852f9b3c42071e7fc4318ce15e491fd4ed2307fbbbdefead46b1744095458d34849b83cd62fa7b97f068d65760ac0a2dccbb61be853b08fe2cda9856d1de77b34e916c10e20f357c77621d277f445ca2372d35042ed3048029fee783439146a7c77be8e448065f8c8e0ca35bf7563a2bd93b65b521d9415f9bd440468b97787a6475af2c389b275562656d68cb8994512a6d14ab40d87e44dcd9419dd8fc70e77e92bd5115b503c83054aca29d7324d344389966edbd2493398796a2e473feb67b611fe42a7094d6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h22f5ced19d55a77e1afad52a29e8b95ca4f020bc787ab48f386d5567c0be3c5ab880f2939980089a3d0481344a014e2c630bb5d8671d680df9abb109398f5546a6b5d5448ead162c1c3addce5c0a6c3131e5d09d845007fabf1e16beaaf7461880a13d4605767c8e02fc8fcf1f492db232fd499b6bd8eb1610f242e5a8e6d712d4e5a904f822c233a60c2ced792f96ba11f302c9baf144a5a71a9714bd91910312d097f6afa6a5af9702b51a4e14859b6f9cbc5a910e20525fd2a0534de783bf55972f0f5ccccbbbb051c69dba5b984e389ea4e6bc5ba178eca129a7f3230435239477071b32d250f3a74639cbc912118b009c8c6089eaca3573da4622fb64642591a700063eee818b4948082f6c27b53c10f9465ffcf08510751b3d691da8a0852ab18503aebe97bd3c7b638a97a1aa31021c64a5f9beb78dc89c6cfec8346b85249877d8834d567952a4d746f4297129ffc3f7f17a3a2dbeac776e1bed791baad91fae434a54b2a2eec6fa3a81e95ccb8a65e41556fb956f8f582a06f73e5588d187ee13d35b150934e25861adb4389958facc4beb99278f655cf2a8b5a37364e9cb8069845747e28d8cc771e884872e6ba3b102f255b5ebb1f15e521c28006a7851ee4e036acb3643021d015243bc0437d5efc3e83f2064b8e6afc396c2b4ef0531b6e9d3c90e91061a329b4fde61c31e3e82e510b6a765de3a4641c5f0e645f9b85ff4812af052fb5957566baf976b3c42f990440defa9872978e0059429af1ee905d9bbc90a66fddcdcb94cd261871bae86157f6640bb37427db129550e26c5da85c713339589358af1432f7f2b44644b00bb2fa924602b23a0d787cc4dfc8ce6089bc164c8b2240296a054d99eb2afb0043d9be812f30ea163bc3d58d2a26ed05890407284449c67c80247c8d0632deafa8546911037beaca433f04987902a00629c640784c7c2add4b9ac613c6563b6c426c1735b382d82a3f99caa2dc39d35ae213119ecfd2881e9f5b205f217e0f427c6ee41daf9385cbd0e6f6f21238185aee7b36d9ad181323a5f745c86d358c4bd766b93c5ee8d2bc7c4990ec2f6e9395d4fd49513628f0c52a735a4c48802c964193083db399fc04f2d7e4c400740b6ad3267a49c9957c18a468322d0b5e8ac27b1df37e52a04f39cb534499255928a64bdd9ea668646e2b2eda40e376efe0a44b9bdc0305ce2549b272055fb4f9ad2558eaa20de54c272c6caae14ee45555b1ce05417c98cc1a3c98c16703aba0acae33d42b4a10a06edb8ed0ea4c1817ba84efc9afd66f2b7af2167938f42116e1d235f626a713456bf243f8b8ee53431cae73f9baa9d0cba998cb630c9f1561446e28dca34aee37b5920995258fad9584efc03d32d77946e92b06136aa2cf18f32fd74d5ccd6422927b8a3c3cd505e7033de86a97005ceb6937ee52535d2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h303b520c01b33c501aae033fe90068338f17f5f3f7ed15618537e5ccfcff3a20dbaeb8b7fe12748811a7ba7c2928d0bfa637e28f0a5712093ba30c9d0e5ec2e67ee03c6b36e3622837b0b0c46891b53e7d113d729ae92fa28201aa8cfa71fd8e4712aa0513543ea798481d2e0bcc952c68748228e63c8ca79cb48eb8a38cecd49f8351a66f3b47db36ed086da1fc74c1d8a63acac2d779f3fb137bd12bf256360fe3d416fdb213c56457d4b6bd9f1f521f7550e0340c85ff40e150d079b97f702afbf6c4ab6e41832b063cf6b5997534d1dbe9bb9a63e4f127bbddfad000a09f9c900c52cf13ca47f83c96fd0fd9c4ab4e385387fd1f3635b924d7c87c05ccb004450c58c6c26487cd045336f2d53775e75de844b1f21a413e16f190453e8c8c3e9116f8596da82c64001d9577110e66fba6f80b5f25b3a98e08e5fcd31dab6bba1302cf5d6a55db6136435f7ae7f7c383f0c5365dfdb3867c46caa3becf5557b60a600ff471b96ead3bab2557382086665ee77b48d7953ac93b4455171b2d146bf1b3dd40b580c1c6cfdcfa5697aac3f6de15955f87a1891acd262ed0671ecc12a73653fe00c91ea28282a7696ecb492b06e4117fe75063a491d2367ddb130eac3ab9b886511887bfebfd2c2316bd8e5f7b0f6508ad8700dbf722ee7fc225a7d9534c25081cb6dfff76af41ebd216e40751df0b57265d32c3bd684cbca8e0dd27e08336f7132b4ed02a2097ae363cd22f81f20c2a8abe9d53e4f39a278a37466e7794984d582c0cf243ad5b77d042b4230738f0018c92ba6354ca96c4f6e5da53b5b3531709749902e01ed0bb7e1bd2fb4ddea620a7e85113cdeda1036c06964bc24a0d2d23d46ffbafccfc2d5d5b6ae5737a71c34d5bb4c0049bfdca461599e86666265669ce8597f1cc8a6b968ced9a96f4d69685ee7b329ebf76025654211c7907c11c6ec7af0d0876f635b00e47fcee2599a19cfb358f790c20917b4540db4b723f4cc53dc97bdfbdc79f8294e49bf4930a0ef76899a93b3928c12218ff01820ed3239528f6eba621893971ee327d4a8233f734160ff7bd0c141ffc39203090d1fdee22ede80b1e66c35f6cfab1970db0e4b56604816d9c99a1c0d5381aafa085435917156a6b924fb7467cdd0218ba849a5d1041356f09210c833206b8b8b68ee54d4a03c2e7eaf382c6335efaf5fb937f622cdd4272b3e4e765ec4fb793f1be36e3dda493505f3a2c3f198f376103a7d3384194e06ae446aabfc8cc6e1289b9ec3e6be85294b2c85ca0762028ee986918e06b1a063da16f8539263fc188b8c1ae85e0ca418dbeb6d09cdbc51a869adf0326d6a23b40f9f8bb8dd1f73a451c0602e7cb8a4243df9ce12b56b116f048b1d6b13e7914e77330563abfe473113df673ee85fbc8f8f59de47671036ccb3e831c9bf34e0b79dc1628dcb141b2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5981e930522dce77eeaed7796a2ccf382aaa1d2a301ce5bdcef7e5cc315dffda24e7aefbf24f2b38a3fb809b1bd56d2b798303dc386103d4084ecc02b45dd26c654f7eb5a4c0a81e8a627898f2953bc202bacda15bb8478c00434d32abb928a1e169d2732548f5c8a03d903b63e2b2aa7fd186b2319bc11313c20e0453304d9eaf6407ff02dcf3a0302baf0232a2b42031d7d0f88039b065f6127cad5acb5c7e8db04aeec003ce13f4c876973430660c12e0901489a3b669831f203ea23063a1614e7018d2a1f7092f4280105e8ba03d63e65620c4247d9a107a16d502c2029bc9152fa0dd84f0c3143c6aebbb22b275ec1e70e0a7f7155deb8abb501d78a95f0c7eba7e29f551b47849bc345c3542aca7c3ca0cbfc9af45036fb588606ff1e40f0d55f35e7d75de509acb793d731d65383b1fe41b62d46815713d2507a2d389badfdd21905f730cb1273d60ff394b04da698e028c6f0a9a29d195cc2a44555965f3ea2acd719098ccefee959f85981613a8ef8972f3e6808496be7b4988dcf8f769aeac2fdd939992faf974d980d859d5ff0db665f0b38c860e7fed8a6761d6fae9174208a08a43c81f07c52f6b3be766cb19e159c05cb50a7d5eed21e0d004c3c99f646f339178aead70b923abc0815e74c92d92ccbb61b5b419a0e270b34551194df6ef34827c7ddf507443146b181e03fb2c49014686e25f3ca228460e9fe6da28451203b3b42df25842df454fc722fa2145ea2319d075d1e92789716f87caf7e23d81d53d5b7a1bcc3e705c61e2420e62b00c78c876f9d7a9a19484fa21b92d5a73820f3df00a4e771e16f50ee06d485bcb36a4c58cb3d1cb753af994bd73b08e6a09bc2c5205ebad8ebb908d71a66acbf58fd2d3054bbefce37250158551a23c2b0bead1d239ecbf373b8944efc97224d811575762b8664300a129f59d2b560051e34fca749b63afb122371077ef42143ed838c20147249c364758251ea48c7172389ba20efc3923c870892ab184ac32eda8dfe14a2e14537255000b3c729330e61f2a099c413e88526a2c193f0973f15505e87457097281112c7abcda4fe901ed6a7eb7cd9fdc15625cf17cd7cf6d325fe44293c0db4c041ade4b654000bb0622c7faab2b062206f4f41cec885869c75f5fc5ea3048938f3e01b51f9b431a9e80ff9710ad19abfdaff422f20711b6e02575d54eb4d66787174a3918f893d395a83de43fcbf6a02958ae1de2bb03005c32ed29e9e4ba8da39bdd308c54f9e460cb031bc263c5164b316581dbcd4e3d9f4e8ca35c7ae4b3a7e0bb14a27e677dbe2a4668a504406e72f1ba2ad04e391d364ab6ad4f8eb071bca30715c796ca0bbeaf9481fb2e82425f0385191c6bac0108d8a6c475d1c51797e99dd4df2bc4791c03aced4c19261f91fea11b576f25a0cbaf59b366112651c74a8a4a86ca;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hdff8997e3c1ea8635b206f2e10edc4c8c5540c5945fc1af9f08e1b1f37148506e488ad2873c956369113cfe24688e6174f2bd28ddfdfed5d8c9af0fe7e03e31402238448509d1badc1723d63d59dfb6e007aa3eaac278225fdabc7bcf505507a64b1d2dbbb4a18a34dddd4cef3d08b58e966b9870022381cb1fb729be99a584421310c3f0f0e585d5e586561b27bf7f3d373e33c244cb1c17f8cf996aee2c1b9f81397ccf9c1b017a0a9a50d77ee59b36f0f0a4eb0138abd28c123cd409f8f7b1da186fca4ba805e5ddaba71508197628a92a1cce2cd9dc14d5e6a64f6a991a147c651acb6670ec5c8696d9ca55fe01ca2038be14dc16fd555408dd265719c0874de70da411ac924c2e1703b6fa94959efe1a1e966971237a4bca2fcf7ac740bb92f3541819690111ad6644fee03367f08b8e707068b5eae39f929b7d99c8c96a6366c434022ddff556cf38f8f8c85fd3f439428b5ac5137820be7957bedbc1596e1faf6c37ad31d70694e513f5aa0279972214e39218accc0f77b465b0d9a8579c1f62ecd2c5c93bc5e455d89f3220752e1b75c7c864700add6f2435367e9239717167649938d21f0caa5c6a12d9d0068ad5dbf4be097a43a033a12920d2588d4fb26e6dad5f97fdc4106e619745117ffc3878ace599e809141cc7df8784cda555ebf00f17fe2df5bee769666b9b1af3685587caa4aff21f6b116c0ed2d275cac12713aecba6df3c75142eaaf40418b5391aa59b23fe8499620325b240eac477ee883cef8bad811986b77781435d6317214836c30deb44a01c4727c0b9b90d620655fddc3dd4fb7f49ea9bd24dbb1fc181eea93a0de4a2995fb1663d5f1833ae1681f4aa21ff674a318f18dc3aeb37d2c831faa97eec71a3483d61ec7c20adefbf266a5e54033712dfd40e31dff7085580860e11fcd5eb9c3c2f3e7d816934b2c90bb8df44b3cea77cb007853b1bd32dd905f478882cdbd0e95f2c66f41f781a874f03417ed41e961bf51905de6e86a73f80dfef1c12caf2d0484628f94f1adedbecdbb0780bb953201c17858f613177aa62894c21de4115ebeec9065718691091446aec009a832966e8a90bcef9702b0bf34e5857405ded975a8f39736b0040aac232cecbdcb4d358a4a2eabb662b9d39a90299586f64f3bdaf999d99badd6e88415a0d77d698d75d5b59493ef9d7581a5f1d154771234d23860f803cdc0f142ac13def3ab7b4fea36ea7be96cdebf63b1b4807f68e5f771efb37bb0a4ff5919c4e3c2109227f712f582f227ffca3c71b6d35495fc9a28477e5d7a6975ebc1c64a38f79b2e4d6434ab99b9257dc0e3383c67d168668949dcc7ba312fd227196584146e11d45ddab0dc4887100d2fe26036a457fd5c616f7086a4133fc6070ab1cff28b27d621ead2d3abcf32a525ca496156bb04b1eeb4df76d89b441ace4e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h41ffff0344e979f516db27923d2df23bb7fd961ee294a37c610114ee386938872325910c8e92f4f1ed08164fc44d2873b7a6551224a33192a153e2c62bf64b87e9b72df311532d1992162505e139ffac4ec828774df1b4d42c54da67a3765b8992ab4dd191f020604092333fcd92d53441e4cc34a0b09a7c7c0583610dcc4f1224ad4a39464089de7b55f58f29ffd721417ac121378bad8e40779c9d299a4d0cd92f3c9687607c70dc7a08847b74915ed2f0bc98b8a5a7cdbab66670de5c3e0a3e21591de598197aaf3d2d802cb9486b776e78933fcc95365bcfe69e7127ee11e06ee12c71a215b91502ca52ec5557724270215adfca6b0a2aa9ef97f4115fccd3fa14fccdcbdbd0934ee6b75f9aa1f79e47e5fc0f79942920e060ccaa8c261636a8bc83be3967ff5ea987084e3b4a0a6119e876b74ff0528eb400bf9837a85c280f06f4d79ca87539c29cdd29bf810eb0c376d05318eaf95be5300eff5fb31b5d7f3d2bbcd3d5b5500975995e394d124af24683459f8361e4612102e83d6cb38bddff645608b74f48a75ed9fb72e9f73bd3821cc499de5b3b4da64d0845f33ee9b40743034ec239a80df1d4976b7a7bf879ec8b4fe2a3fe1198b1c560e5b1e2f33e145a9139ba77afe9655847dc9fefe169d01b63eb288315f18ab3fb3b203455dcd4ddbd19fef7318d51056fcc68a2b472c0a88996ac6cc43783b96ce857a2a644891ae8a734d1d120a24073ec4bb7ca4c4ac95eb7dba523285e20c08b5afe27cc82340c6a81213e7a0433b99971930a33df1363c4a1cba52636724b2484fa2b3cce3eaae7a656a737ec252db1d8c0445158ad24e039ec0ae02c7ac3da4778345b2b59604ddf398449c2deb5fac50256f410e079e9dab87e4700fb680b1f893ae64c2397a4b031f16448a0ae67fb5e7cce11258da650d7e919b882cf2c86a5d08e1d5f38d0ddde1849f2c92cae9ff23cfdc32e72212c657f2c7a59489b0363915692691d3929a70e39dacc639931417af33d495beee960e5fa4034930f17f53d557d5636c168ae6050e83d25d8d0844d1813e8982dd7529a4dd066bb03a33c3a56fcf3a4fd9bcdd0261791f07aea44dd66e7a606574abdb71206eea13dcdaf11ff296294f829ac3f86885da477616e12f18c21012453940eae30399e8eacc512fbc412621cc95d0e4fb92c09d7fb6c49bf97dc062365c10f7bd03841665a089bbd08ef4d3191f121c6c7044963fcbeedfe3a5713c5ba7c7f824157119cb3e268314596e8577e41ab51158c21bd25f47f831caf031a17eeb8ec2ea75d42ee9d2ec17512397cac9d156ef37bf96e3495f286e3eb4515342a4482bde2610c7ab1cddd02bb5d3d299dd88188f4b6d1c97ab2971c17e6d793fe1f7035e8b7282821bf93a91a4325151faa265e8a3ee26069a2847394b5340df46bc9af9858cb41e9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h8038a448cb91d5e2398aa91fcac22fd9d40d516a91081b9f6b36a804238b678371eafc6b00de87354ff1599e8675663eb51d35b25416301f1b25b665b1b0bbbf8c26c30aa335d1c4749c04d7500071512f1dd03c24f587e84cc7a9b22595e5de634ecb39e0b982c0c1316f73c71c894cdf2139fc589b8463e86ecb18bb7c8551b8f11bb442ea31b59649613aca90e94b4edd9e72b1124ea461544d278d2b09cf9e05ad30f17bdc238982cf4e29967d9e42e9338fdcd9dc442aa1de6556125b7411e0c6a27fe571c870d46166fd515cbcbc89dd03b9c2b04a6ece8159dc3f30117041bb9193149c25e7b98cc2e820b1f92ba624842625674715aca9511c3a5b30f047f47ba28c50da34bee9157dda8fba86d95c47400f88468b06817c23d3da9d4871d402b2fb688fe1295dfae1394f375ef7fffda54cded975f7d5aa92f72c76aba9ac8b0a2be2a2769e0cf1fd807d564fd5d00324511b5f5ef4a74df8e2d9be57c52c3d8af6e8f97636ef2afe787620b958e6a49ff9358fb9bdd1d64400d1e3d15ddb6d28ff31aa8c558437ad41e407034c5fc2bf8e9f8abe59340157e9aee5c0807a9fc5a11fa8693cd293d8a2910311406a2cd6902f856c21f151ae587f5fced14e4cb84e80215b7c611c1a8c7e2cd3ec1b6000240b4b154da41d55f207fea7395ba706a902dc60a8ee88b6d8b8bcbe2b10810f5580347211c7bf66969eccd1d4cba0a93911369bb539209a4550dc3f29162593c807f90155e05125d3f98064064e2a7e733bc2bd5074e83fb64eae6d1e30a1377c1c3247d6d2ab53764c2628f6a6ae7eaeb600dd9c1ebfbf8b611ac5c95cde6bf8602a2b2c4b065a7f3f02f094ddfe5041dd7f96f21bd5b7cf414e212fff8125b667b30d1efb28eebc6da1aac610f1b440cb69eb084026777dd2db0cf6e48f6e6a0f14381240b90c48400b636470c88eda1e9beb28136cafaf0b6ec2e646b37dfa2b3a3e27117d371777fd3143b71339eec601c40eb6d86f1d41757c60ad682ae369b56568a918e424145681ba08a6e4caa4d5713420a3e95d2a640fa6514b893b5adb7052365844b17825dbefc60ee58893fa72bae081b19e7f006685b69e1dea2526f82eaf269db8f2ab0b54652dd0bbfaa305b718bc05fd47a4d063a6047cf3915163c7f2a8de09a922ed599482758a8161f3000275c957d5c4afeebe3af99783f44d9f29d0e9d4c63da14088aaac9068d7e5cafcd57a2ed05caebe822e529dcf86de9a886dbfda7b8c9be0b39f14f2c6ec15924ae083b728613d15fa526ebe3cff9565fc7318a7811c2d096e071df6f6b8ee8245e8118b400f266d18beee9ac239d8db79c08f859f8cc81c3567cbc7cfb5ec996266cd57b412242cd1116851d4e131f5ece002f0603bcf45f60063b70d8187e5e5ef6330f86b44d26d66e1dbe727fab192040ae86153;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc67d9dd878c661453e93a65a51e1de6d9351f3f99c1df221cf881804550465381b929abd7cacefa1b3aabd63af563c43f07fcd9773c5d0c2187a369410b87d2c47dec395c49049196de720f072f19a2f45b1465da7b75aafad5ce352bb905b6d29294c533a529beb98f80a9bb7379e8985b614b36578e8478e31f3841b573659c9de7d3cec441d945008c1be4e998fa10e74802ec70c980a5790153df665ddf8e7bbe9a8d66ea414cb69664fc3a7f9cad92ed30a6f809d263b60316b87160894453197ec653556700a28ddc087f79bf06dc8f6191ed1aeb0db1e3e0c035ed218c5f3398610aa7209c3bcb4ede027cc2737f9bfe82ced378f802b88b82aa6f78b89ac1bef951728b8fe6cc102ed7835f44cfcc533dbe976339af38ca6dffa29bab5625a9f1549d437afd19b82c1e73b5c3595d30fc2aafda4b5425d2fd343b3ef20c5ce3aeea7fee5f5012e326a8b72aeb5d1e4b3c7e0687b60a0c08c665c69945de693dab1cbcaf1903dee8e8d1242fd87b0f70bcbbdaa11417c3321380c7304f3042563b2e97224fa13a5d7d34422a960a0f98f1ea7a5be8da1e7ca25ceae75e83472538f2bd2df168dd929d1edf8ac48af4a61ac62257da44331e5f7e1f3850e781262903edd345f08ab76190f1603136dd2e8218c086cabeb08dacd6e6e9d21e54ede758ec9efcae1a74de5d9ef8a3e0c2e30d58708c4f96d913d53b171aa5cb0ce09c10823f1ca3a4d671728e955c0cb88ac807bcb4b0fc727968f4b2476c9fcb33dfea1d41145d7a560ee36d3af903b968c7c71770c624708bc4070c730544bcaeb388b96305be2ad966d8347c6d6053e71a5fd9e5a8e4a1ca0129670229d5c5445840b78ed98d8b6eae6dbf110e31fab17e3e57433c943ba43b115c38d7d07f57812e2c22806d90cd954709f633becd5f9a376e886a22aca285c387d68ff1728dbf25ec600eedff12139cda67d784d1530b214a6395df41bea4adbdc3508daa1c1ebf7392d897e4c8a1b83b70d0c26a7cd233c7cf52a484a64eb4148909fa20cfe69a3bfe3fb19fa0508a317c386b99ca663b1dd7f549a8162a9b8cb16915b13a0d53c47b960851bf4246b5c1aa737c97af7896bf5003c0fb098181e80c898ac6dbc4253b729a8bd16d1dded1fd068fefc0efffc66b6a360abf718af06874fcf6b26c194372c86f3c6ef540cf5acc25ebaa5940da2bb3bab7dff2c082db4bec9b7b83b7d4f70669288f4cd9bf53aa9c17bc0a3c1599c7ce272273e6e951e0a0fb55aabeb4dca93c8921f4fd6e7c851edcb8420de84eca3c98f28d679487aeb4752b41639018263e976b65881d41fff659c5ff2745cec2160d11cb9136395b41c07ae71048ecd982e2a3333e24a3e2f9f35d1d98818c9b508ef70c15c96cc2edd916a455eb800d88d31fede75c1799c23f2a6b52422df2ecfceecfd1f7f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h29e005a3be6b9965d78f7073a382b7f7fd4a217c64db4ff3fb067d5f8989501725fade88a467557dd5fdedaba9470d8bcfd35bdc1491ad9afb662496132287b69a63224d0acb3040e581fe812896a6409e4646482d54a932b257f70698edf97b9f827077bb7c2545f3ead02747e6485ddc939f950e472aaa944471c7977132ffbd41bc708d2df2d59a53f7cc5f916bac4bea17fde731aba5e88d4eff23816eb9045dfa12b51c81654100a02a04012ef4ddc0702b896b97475bc2988874976960da1cfbb21b1bc541d8c249a5196c4487640ba0b6237fe084532aa5b84ab942f1f4ce8f0575617de8e895ff183a3fefa5f9096fa6238d0e66361ef501d483264be901b58eaa3daeab8135257692cbed55d0b6c6e008f4da0297aee8f7f9ecee60392d18d06292ed4129810ebd2b4504ac0a97f9dc398cdad3c16adb09b674a534f132e7f306ba24ee11b0afa9656f8edbe5c8085bce8a6d2e220e30280f58b25ef18817f2a9bd81219c27685dbb8e1cd9867ac8448881ecd7033fbfac04dda6f000174c4f785309b49d92f3298a10dbdda470f780acea9a3e83a42263726512178bc0a77d56be3914d4b6aa9702bb8d0d7ec13160e324e06482a271422188d0a85bf87ee03e3b8d0f52870a0bac3a87cda873d5a6cab6db0372de39015c61ad867d27883b63eb9b21e29ce7a49704d4bf70334c6e53714858ec7fa8182b95999b25bb61e2d27c2f10181eacf356c55dda78b4d822e1f9ac1d4159392270056260fcc248c9a9f6364f25778dc880310aa4dcb8dc93f465cb96dfdd99eef7e5015a81d9180bc55506e78fb4b9c8aedd37d583fb52b8f50a23c00709775c81be467ed450c75d919335d6e192aed58307685b688e19f61bd66ff171bcd6cb74843a33de6f753993668b7321ed476430939de2120a7b37da6ce68e39ca583a8d0e5c72ab76f2291236bb2311b812acacfaf8557ede66ad51862304ac0b1b483e1e685f49b627f058ac15ef15a6bd392591fa01da258829c929222888c94a8f8a91120d0e9cd546cde1b10a97a430c9d131004444d40625e8d12d9a5c7f74150e0472e411bc16df9b2be1250d3d5e377111d99757b2e59e39f0631f27047d96d5540ed109880c721ec73e12e69c5236a248fe3b7f7a452cc7c906fc48c04505bde3a065f01b9745092e84d528b8930a776d829c2929f4435d8a1a442d17050ca67180184f08106ce783999ee48e74d4e95e05a63e08197d457e489d171c4665910fb29cba78f53f41efed0a3d84435b5ed5f355a7e50e3c9ecf6d148d83c98948bb1c5d9248010d7e01c43ec15385f80df22004178535dcb53e7fb1545b4d16cb02c4e76173f2119087e810f740e2b7f29c3aa90216bc447c003bc2f3ed954ccaa61669546c0581cf0b4e9748c8e1f4048f0317eb469ab890fe2230e2e7a475f542f934;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hcbcc6174a573f67a3ffad1976b2622312ceb93e62dd9b9542247ee0889348a4b68983ec9c802b35fb405879d2cd66ba2e0ffc9ebba7a4eb38d80bfb23d8917dec994ae7c86a67076ed35c3e930663d5dedd0855add1801c3697b64778a65de7e3db89a186a4138c316f4e9c9c986cd14af8ef7711010df92adf1262cf9851dffe9208c474b1900269c55613b10980ea92a13bb10e2b54e3f477a489fbc6fa7377edc76964e735a3d278f6d50757c899c6eb9bcca9a9a75b95999581f981a0e953216544c3e308340b23341747e96ac68c1c274cfd8fd06ca77f5c881fc38a772a170765dff2c7160641e7c8f5e7bb6de0789e54526c16e9e7d76bce28cddfe7f4678345c1aba0d72f10c18326e736364761531af4619d80555625221f9f8f06d7d350ae64c4810b8efef2e8d86034cbea297a365de54a3923287ff53f2407aaa904978cc931118c41313e7742d246bcb4f46f81603d45a635d775b717e28b0fbe2b6f4f243cb88266a63cbac63c6605ce92e3ef02ef4686d73f116dfc935feca1c407676f94382376a7cce3c1e459a6ef9d03f79155ebbf2c7873ed7e0477daddb9800a4a71b51556dc98e2f46c9ef35127da6bd38b4b0002bf52d76d4cf099c233c8d5aca6fc6040cacce3ccf6cb64f153634dae668c7f50d4b516df9ffacdb14e1c8479aac5a6f9438629224951a1c2525ee6e1ff7e31a80ee2c027e7ebc18878240264881ff7ae556ede9c90f9f98c88754dfad552689fa5a279f1602aba7f207cf60baa01154eb721607ae59d78522a0c78f7320d48615e51be7c928790176c20fc33392103d696efab1a0cbe50c3d0c185f869df98392b91aa332a39a704e154e50ea7368f1268435b09560a8e96900f32ba71437374dee7373a4225cccdca1051891de738cf979c0946a6027b397d9a87acc425c2f219ba21b685514e74f3c85cba032eb85b2aa571c869dadace0d2c428d5393e92808e074c3d67b049870d01c0b3452c7f57d38fb63218ab42b2bbd81c0022a15223ce282d33a4f298b97360bda914b332dc6a20e3a3c48985da9005a305edfa27d7790d3f805f03ec8045b8a7659d2f0b64dc359bbb799e2337dd65a68e9b96496c8f29bb70e98a9b79a9d3949eb16145b22c947d366f9710bc9372dad61494c56b086ddeb446dd42aaa09b3ac547a42745ee5702de17c4bf7424087687221f966ebcb64285b059820b74a8b2dd6a663f574bd34f9eaf2e274aa0cec8ee89db35aeae29e977d4e38174126280982811974adee73a65a4da55f7068a539ab6ae8f1944dd780b865b0d0527dffb76c2a718ce212c287daf30a4db6cfe364149b98704809a2aa613d386a731c25b4bec7c43014d672c7dcf4d16a0e7422193f5d2ff5fffad386eb279a77e8f6b47976f3ba80407086612e79a3102cea7f7d2a0eaf4f4742879314e0289;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h63d14c9fd1c0ef59bc28c7d223b374c3534da241cc005120f4e4e79f93c3dcb398ebb45a243ed2ba1b11d709475e1ea6525ffd680474589bbf09442f61b89d5966cb8e7383bc735b02be35b0e0659fd7248a023c79fa137dfc85a313ba33fb287eeea39b06c8ad18a00f6bbc2e84da3e6ae5f6cd580ba6efd5eedba8dfaf051aa106d9e6a76937275f7b199307bdc7faef912a248addeee321b4ba33f7b1c1599f72a2811aa82dbb073b321b937a0d978d2a8e881bc45955cff92f2acb4437a408458f37ccbb4e3878d6f712a7cf96a731859854414bfbb3e1b7c131b464a8997cefbe05266c18839587aa2b21b357c99d391c49d3b6f9db10bda3555ba07c05ab90db71c35db2fd2f2f28fa7acb37ae2e8af748c885276c22a234327f7ba12f0d5bf754ab2f0716f2d10bc496cc059cdd9a71eff2c056b39186e6ac57c103fda722a66704e696b80956d2513b80ce0417b16aa7f92781c073acf4c386010b922533f7fc2223736a798f534f5d94a60a1eff7011e93a43c7fad3ad2b8676eef1d13e1f706c16252764c4429c9dee4b997bbfea10b01832ce046f7f9ac0f6ecd39e76a8b19d12fd1e6623f2c37236359484ab1f67946fcd5380483f7411702ee377d9776e7d5de3cd9d041229edf2447aa7b932734b2b426fdad4309a0f878cdef1f741da1d0a479286ad9ee93422ec9e6ab690d144056e5011a2edfb020bdcf2869934b3b1f21d837e2f991cdbdb997c9f6ae2b4cc1bb58020973ce0ce05d07b3d266dbc117063c05801430b54fe87df7bf7f29c40e224f422f60132ed7ca7b49602ca504b1bbd7d5fb18800b85bd248a8be925ec31fa23f10cdc59190d805df31240c1f8d872aa298a9dcae2f0f318beb437be72eb1faf24027d5ad1a0fadcd2096146443ac93eaabc14395b3b279c93573e7a48db43a387e17fa21fb24dbf6c6e28852cefcb725f24f6483e9e22a44e930cef9df7a42f3665eec491ea6302d3da7602013ffe25afeb0108ee38a5dcc87e6e934285e20ff6b0485953e6657e38c1a97836ba44f1bfe653c20dbdaa5075760ae4cfed520204780671aefcc9d87818dcff37b66dee49d16163ef57a65294a3d7dc142a6a6e9328cc9fcf6c3d98892be60e522f6608bd6d4bd2403a8c7a5dedc4be92126b590af9a376c607f53f431997fe64d2412eb0a49a944c82b127d4a58e263f32568c650c950a082f35c32f1a25bea43269b1b7bd315b5e9ee3c581c5e1c56294ac645ed06bc29b0bee392c59efcc27662d6ff9224e1a4adcfcf4747ee4feea0a69c1442185d265ed0602634b9c8db0fa44aa743abaebd16738aab76a4b94707e1fdb316299dc2f4f994a54150469386fe6f6dc17905d822c7c57bc07acbe97911bf64fc1b0d8e6cd75c2c236a6da3e23aed002c97490fd0627ac9d5635048080fc6cc99ce45196cd0f5d9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hcbf7beff15583313f29a0da971698e71b4a4c419ad19d048a6e5c77a1dd0e7fdc45a27b5a908c3df5233ee5ba7023395955a3e0b168be8d7f56202487a590608ce280e151ef1dfd7b00b7616c7e24c7f9aa1d2f26355cbcd9673b810295abe2dec96a21b4050f83eba6a5020c4887e6a9705d700e7ba884fc1046baa77f3c886635c50e1d2a937034993f193e9b56db48b1c370433bcbc592a7133e358bd8314b4f3ccaac21181b36805d9db71d66b1043b9eb757ae4a1c68d75be04c1566f940b4a0434f6957f262aa59f1c1dae9f70360933c4a852e51c89133d7811a0da4d907ee8b67cfe26de282688cdbeb4d542606fd74c6b15786fa5323e2e5fbf721c89d8dcd55db46e46cd84b929b89c87fb7e67041087ba00fa8ef8514871ae34eae4c60ec906680d3cc6dedf0d18cfe6a7350420ee76429a10921d71523135dc51dd1776cc4f5128b06dd997377da1c01bd1784f3471ae73f4dac987fb031b44ffa10b243f37d73a55d9d21b2ac125660054dd097912e10faef56d014b77fb4cabe50d1ad2f05a6b84f14d8c50db1eca8a41736eb45700b44d18a4473601ff8f944f18fb50aa0ed0531b2945b41a9ed51ad5baa651d76e10915bc67c98861b157e364f281c6717c880ea6437e82885eb6a409da6812168cc87a7dcfbd95eeb86588ca1f7dcce8b5250b2970efdad6f910b77b72e6f94540da9a29510f41cb34438e56fe35c4753a57a89d3fe433240771ac020809ce2152a14eb18259846ff7ae99e3ee20c990ac3f810a5fee85216aaf6e9be43b93da0d8a403af507ef1041730d6fcafb05056ede84c77ee24990ac4c5204a5d10afe0b731810b4e646d3c71d42ac3b365646197e54b4709ab6e5335f6bf9ad00ed4a34e6accff2a09c3a5e67b175c3f5449c44424c3951c25686f80a2dd9c41c18b9464e6e1f6e1388380280edf01d32ed125ce5a560250e8e4a6b2454dc274f4ab2b0225fb60b22662dc279756e987073c31de46bbf98964bcf75e9484dab44dce944a4aaf26427a4aca601c8b85bb266b3804bb23bf13ffd2ea97c150bd980036742d0b457e4dab749374df6e6525910cbae9c5c43480c99ee960c4a136c633107041201734c6ad1a6f966ffdd5d6bf432c1553e449c99e5ff42a76bf435bdc3c32a4d08757140b72184236d2821f39216def771422900655501b8067d730c6ae59b8fe924bab039f12cf0590af4fb4a2582ff1939769b6844f724b8d7ada29be14aa43ca604a26094cad59aff39b7b9627eeef71f9a7109e9eddf39255149c1716a35dd1f2a1dd71d1df82db28ce8f6046d1186ea6a62bcf92b6f9ee6056da295d10d23f825b835c2f0334c72d4f397fab106fe9356dc9689d1942b38f0b9dde62a8c6de55de38b600aebec77ba59879a5d481336be3176f9ca47ef7706c7bba982ecfdc1bd9fe7c6a8f25;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf0dc845c0cb99d7a4acf9110896f74dac3bd9b56367f303d99de8fd82b849e014dc61d6b5968f3e3f440bcf0f0dcd2d3ebdf2e472b46ccc7470c0732b5f71e3ae35a6e689bb8b727458b70805d2db64e880c287d9424a09e4e993fbe0741f73720ffbb9855412dc51730ba0dc76d512adb10c7cce22f2e65371ddd66aed59cc781856592da83ea734c948677675a093d708c7aca07eea21a591058b41c8f1dfb7a430c1062c51941ca3621161881f8b66ecda1a467568158f38cc632bec39f2c4002440cd77448fb261150482fb71fa46919be7f3745a273c34dcc7c87d7fb895823bc482894390e5f4798f7f552176f8e6e78bd6cff1cef4edae372463c6e758c4e885201b2eb4df2e878843e626eb529ff043f96eeaf999a6f8ced711004e8f967493f846c2753840befeda2f888b67d69abe76da7d3761bd64c0e541e8fe9e5548bedc9c15e5b574b053af8a41cbb293add1258f3612e0902494fb618f8c602bec5220c551e901e8e870ada5f99c099e6902cd372db3b76144fc0e0eb734dbd32d8130a47bbefb86567c8d320dcce058fb96b2bf2e7a121ba2b87141766583076333a6e17d32575dcf1cbc1005725fee6e44caec755017516ae77513c517d6292f33bb104c20b868f814fac1e116b03a15993afa024ca8921b8376c2815214a40490f39b7b7404bf37efe82466ac4bf5a29c24dfb318989154722e8c6c0b56b3dc11ed6478396a984a2c11e082a5965ebff4b12f37958606f046fc36c60cb229e0a43bf92b1de1a68dd004296e271e6923aa0e6f0583ec7fb5c19802d3104a8bd274d2620bace9be556f004e2f1ae62286198525bea6201084191f6d292a8c21528ea0a7a76787c64eefce52950909315aa6a295ec788eac74f227fbf4e492f9f2320db5d99bc2741e0dc051ffae3c1c3a25fd43f705a334d196278e961e973e57526c18afbc726014e5c90c25012f84c8649b341b9975436f1707c05b30e5bd0383b79d75e4bc042756679d42a6d670213f4dae627652b634b0998006224fa11e4ae153c8f7179578568ba36b6c0f363be75a07ab25372b2326a9b2eefcd64a31d1d0abf5f509a90ae5de68a56e47bbadcb7afb2e9364e425f4d50786d719457bd746f0d2e35e1eff6b9ef976822807758a1ef05133da58b544588dcc0c08a42b46d51042d32e5a92ba4ed034b0376cb285e3e0129026fa581080ae43a5d90a34af6292a12d090906e66daefcb70009316a099541a40e04ac605c28306524e607b5310f403262264d0003c0af19d0b3bd3f783e8e9579af96139f8f7cc2f99d6c0a483dab93d85fefd6f9609c0c4c548ef687cdcdfd1fcdc865945b433b6771cf759bb04083c4ebf54e861f4bca8ab3df55aa4c821058759180c441312617ae29993cca5b1d5734bc435bdf04dbdadab1cf88ebc50dfcf59ac20e4151382;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h5768a1d4f602d175ab69aec9578259e3813519a51a5eb5f7c7f6ac9edd354853cdbe7aad1af1d56127b2928effff4984f058ee13ca691dfdc4ab202b69a443eeadce6d7e5a72b93d99f085340ac1e80e9b38662beeed933e5ef11bfae60e7165c0b20397b5f4a1e6ca559159fdcfadaba6921623eedb5070db8c81796c9045e226bc39aba77e253ac9e55f8c34dbd5f8dbb46ddc7b15dac570c519371dd03a4e2d53934a59a9adcadbd4e4cd4aff5a8937674e03273b7519c5fe364c7d949f9c46937a3033900606d64de70a7b60d3a9a295466d577e00fc1beaaeb1663a78bff8d875d1239d5970d1da41b012ced0daecdfd91236e914d9a8f1f6cd97ac38592cc24d2fb232fba4a91b72cc7488e585051770090e6a9ad1cbeedd5e51a04b471864826f33b36740faed6ced85764372d81d6c94df805553f9ca054b92bd1fe1b782a92d307e6629163e3b70423b572e842180610f3cf4018e4cf2f6d8ad910419da42fb4a8f670615753a8218349dfa1eb9489ac56e3d11a97b5e3af1737c53b2a3d2d29cbd0d026be9d8bf2a5b29cac79b51fafc56f045a5ddd5dc8834b9655600d200b84570d85796b081f8e5be00fe79d0998e2e60cbee2f374ca7f8385051789dca1267b74fe1790544e7e17f9daa7c213850f5bc001a4b3b51e15f82ff2b9312701ff9f4d81e264e4ed77fbd4f24259b4323e9dfc7cc46d82c425363529977eb2f95e2b5d4a7912e7d7b2802c7a16d65d93791cb7456a29184b5ab4ff39184c9c68f8548b75d07b7736e3facd065d7f319789db3ff7f53b0f549470bf6e7e335dd885ccc0247d7ae24f992adca5c9b51c19cf4c3ee24908d5ff2e29ec1754b681e2473691365afefca030597676de51b737040b2cf7fc0a179455bd92ace36ebd8c6fa4c4ee90666270a35306e1fe26bbc9c2e3e3be58a9cc6b5ca04e92b3b397a2075837ff916607ef4e3e0cbfa1610eebaf101f62a950a374ffff4509320e63349eb468c9f593ad71546c223975ee3022179966871654e008156537052dc02c1720fe5fddf0b09bef659355701515bfa1b58a1389f27f4686adda5b41df353b93ac3aba42b7c6384b172a52fc0d14afd0b103b388ec5ecb9f9f01e9f4997f5663842d4a64e3401590ca61534425bcf501cf5f787906810bb01aa9a563dcb81d0ede401cca5c27a46d2f04b5eb9c43594ea7494d8b7526dbdc4cd85d021a3d981a837d05da3e2ed43ca0f93fbe7c76c91830377c88f60397ae0e40e1d0e3395f8cc0984fc9b8dcd505c85a35e1b459fb3ac23b702955d7e07c4acb976b77f4cf13a81a174b4a71f4f879eaa0017576cbbe6c98e937aac2c313cf5b5e1bcdb510a871f0f77107c1aa8a4c2ddc7c71e9abc9786fc5b437729bd9f4ace52538124c44bc39879e413f0e2a9223916896b4f608ac42fb0ffaa40a137c7fa0a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hce612cea8950d5ce5c75585551481d5ff2c8206442ddfb8d330dfd177c511c9c6a9d7942b2a86d701f2ceb33d8a50af43b5eb76d06ee01574a1b2ca7fc811ccaf1d232be60a214d4aa9b3095e3cf48d38eec00bfafd77ef48c79fa33c7ddc02468169c8e2e1a858e15ba42acd54c8f40c24698493bb44da3aecb59141920179529c975c02e013961ca38c02bc6f0d6e91c9133c4f42078946d934fc390ec0b133cb6550f025c62339552f0404e193edf50959dccb81972eb79c539c4eab503ea226241e305124894228e1fd5f977891e116d88e8b66c9b44398cdb365cbbe7938c99121007f842937723b42d726d0f1d6369a8c64e87bc0b65de7f1cbb55a210b6dfef74647cd0875736efd39e0bbd656b1a9934ae056e95784f78323ba2afd9b4452f01928e235fba5d6cb752ac7a258953d042afb1c8e4848625667295cc4555646bd1bb55772a0f391fbcb342bfdb71e5f9d3ca83cbc8fc80737f09802e4d5a2fa3db860e0ceea44abaab8996390c69e35836088eaf48566d380a968b2c71f8f34617ae1d2e794881faa78a138f548fff60be9b9bf147fc9702cb2bac378e72e8c75960f74c42a921a7557156598faa0900112985e68823fffff53326c0a2157f7059237897761a314fea44572b6bef17b07ee07485ffa5f8eeaade9844d0725375433e5fce653bf491504ef720f95ea70b7f0cab10a6ca3d0a0171fedebc61e76317a7ecdb43e4c08bcbd268b4059f8b45642336820c7929986690486f390bc6a804040725edf511ef3958f95c8a0a44ed7d41db9838c148bc812905387e42e470e9736180d623c2ccacec2de674a214727277cd36a0daaa78bbb636ff7935ee265a6bd487c6a5785c08077f8ce17efb416a5750b7b198fe857975a4a039437ed336225e24ca12d0e119071775e4ff286cf6458728cf108040ee9890ffb23da8002079f071627f227d7d2ce8d8dd240631a663561809953ea704d9906e426c3269e57d7fa2c7da4737e5b1367583da0b626cf3b1b566a7bcf0825287c9fcce07a00c242d82b93704874f26699be70d9d965354d2a338f82394ef4fd221cac6a8490ed95ae95be372cc9132ab2e44c9825bd85a1a78722d2cf010f22903c7979de1d49d8e2a86df80f86f9c7c05ccfac8f9adbeba936c143bbf8af0ca127cd76409bcf1982731ace0dfbe749f2d53b59202c3c0958f5c552c7ce47f559f7d1a3ab45d14d4fcb0e69d251146780cb98908561fb4f25cd1d4040c88c88dcedbacbc12bc1923818a2cad1513f6ee53695e3ba2fe6cf035232674f4135e2ea736c82f033c8efc481949045dda614f57a11a6f89601a86ca441cdb92a1a44cf5f35f99b760dfa53cc9a4f3d3730503895495b9e405795bcc068382eaf9818c6231cf3ba14375f6eb169b9ec43ccb45a65b46e2d4a686d3d37a4d424319094c9fe9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h734f6f1a0b4d07da134731907b628d2ae3e54714ad2624d755e3f9f02bc55a41bd2873c75dd1deda70205fcc9df33d1b909d74557852cef2745b4c1247969910aaab20d734eaddc40916232a99c8b1d18b94e17268634d38fafa4f77f08717aa80b69ad58ec06bc8526b520af9245d13aa8e7af330db1d5ad4b9bb161b931f867a8cd3ec3af73147a760592c08ae6dc08505e0b7ff97201bb4faff014f662ef8d90032e74da33a578ce25137ae1e19c9601ba23769b3e99a65f4ccd249b1fea25a497d69c0519647668922dc09795c2abb001ed7389f9ce7af5fc499928cd2f4e98c2f38f3335f4987545c3ea916f71531ba1bb1b71dd7402d1f4f0265b1b3814f3d915c47e815dd5f719ad3a2eb27e44ed5c7b66e60d0427744bc6cdfc972a4e0a534f95b39c0d9df7d326be5ff852733449a5b3fe12dcf61785b66199584f3baee4cfc894c5d43f2d80bc53f130de03f1cab087fcd83acbc8049194581008ff721b07f7312e6543ae099ecad428bce4a0f24ffa5e3b378915dbfe7affb47c12c48ca6cc2ec41222317a60d5746ab8d6c18d8469fd58dfbef7ecf8642ab00ad2ba743dab685aa008ecad49add4f100a5c7a46157e78a7d7c5513bf3ae480b537bae294fa415080cfe2035a4a2717e1218b16b3380a0a2f37563cb803a43eb044f16281f42accd945984c202651498d62651e50216e766477b46760301d3ee387c44315d40a55dff92e059efaab9971d3e88e8c3b320573b2bf0a0f13ab6ba831c460beaa9bd2aa6ab59df893ea7cb7521f6a0c49b730700c7f4075d54eef4c8df8339d5c3dceee6fcd31b588ec94d18adba62745e91daa1339b83f8c054f7264a5c69ceceefd4067f39e020e5f905b406006d6fbb0485e5e14b83441cdf727258c5ec88b8989583a7d176fb0f083149e947be3b56f3410788815c38e3bf1195b4bcc660218c97d5b8775652be3fba325af5cf73b0b95c9c43dfd041831a41a4b1ff6369963ce9da4f11a3370eee360bc4f5662ea92ae78c212bc8d197edb0663aac3a256bc575cf8d476bcfe3fec8879ab84c67666a111a56376631c5feb4b973872c21a9e220bbae0b17e763417d42d866a21d5a22f2ef7a0d298cd7f195532b4aef03b0879d978196a96ed050bd595421eb70af239ee5b03e1585bab8c142e181e146af8f53151165a28f8819c9d57218c324fa26c0405e6008d06bad3183031e63efa739529f54f1be9a0841f24b57e335edbca8c1c20a1413c39528e290339d846a951f3a30b76ee0f6cc9844bc6b64b2a4a4c92ee437fa1e3ba2ac3bd70037b23fc134cdb0d2cfe25e440ac2de35f041b7be3cf253bcb1d966f95ae073ea3cf1da0dea25abd9216f94bde511c76414465ebc1013fa65ef7bca4aebfad85ccdbe8b12e52a3640b492e52755b8c56193f7644f9d503ba4d61b14716577c7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1c5b1e924943ce01b93414171f4176c3b6a140528408bf6424f2e7ecd18c6b494fadd1a75d88cf7a706095ac251b79cfb1d94054fb17ac6dfaa656d521ef3e2ca7279b997ac06c8cae69cee062a4566921eca668234c016f6642600de7c64501617ba672994607a7bd9cd40a311de4ede11c3c21152ae8e3728b327847f3cf4a6949fab4d280f5fbc7ad2f90b5d7d38afe301c838f06d116b659e264fc3b1352050f76a725281065be9cfee660a86055c95094408de811eddef3b6deeaafa576308f453e1cc145f9afff37898fd3982940d597dbf861fb4ca42ad4eb84410df6495ba191029aa552078158fb3ed29cb4c616cdb2a8bf0f572c3e233a8e80dc8018764387325ec7d0c60100ac083e3cc51b44bb6b61572d87ea78635e95d84af70568d710c2e3170070ff3de0b839557e45bc6d99036088d154488a97e3ba192769deae46983c6181fdb3cead50e893a8d9ce02b2a09c95169fbf4f0a3b5c358ea9fe5dee8ceef706acbdd2161128e55d61ecd6c514b55c8efaf06ccfdfe13590d1f6d793f16dcf47a073fab82b563334e4dfe0e197f83b6bdf67be33408c4d6e1c01a1489c853327cafe4c616438769091095af8beac0ee69016f4582052ad23638f9b6fd4a4bec09a5c4024a9623b4736560d842c4e4ca9a627729eb8a35200ac585bc4ffac557bf9955d0756b6afbf50d7069fd698efddd896f96b2415e3a19a5822250579e5405eab57d310df8ab39c31cb8ce8a63380d01e69773ba6c4748644fed88a20449d41e074dacc6c4354ff4a7680e7537cb81854db741e0ed4cc2a88c8694b585c3c07d69bfe43060831e50a8b5adc29f4abb9be7bd3ab6f9291d4c9970afee2f445649e7480ad7ea2bbcc48475c832415c17309b6ef37e4e0a7b71641efb30e20622e7d696974046c4c53491f48b11b7ba4ec7fc70efffc015c03ba47dc6ffbd53f86bf915e8330570b08a627fb764887272605cc07ad9e5e0dd84d168be2b56a4d8539978265186af1334ca82dcdbae9c5eed3bb9ed9ab09dbcdda5638b6f16312548e86c1f9ba7a0ddd327e323e98ef4ac6d6ab897e9acd4ba19ec291b9bcc213b9fdf125710ffa4ec62beb28009ab423e50165b0b657229df3f6630fda58d0d2908d0350d5d862e24102f9818f47627718e9dfb22f9d9a860faaf130827143dc9daabbdeb5a5d28b4be349e188bb5fc6b00e263f835327795ec4c08e5b8f7d3f6276fa708c8604186ee94a6d983342e16e0dfa6e2edcd2f872dfa1a991b7e2c81614f33131142ebc4ed3a1a93f456b7e02b05ff57f98808108d4b429151e6b282d56082b215239203379c22c2b71e753ebc5ab53953ad51547e685c794cb50a55243992c6a5c954846a5de52b3d16d66778cb714aa1ed1c8e8f7a375b0a4c57298751f6792fd1afae0f3d3dc6f6d78aaf4799d8e8b315895;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h1bd60ee40fc5199fbb190598bb4291493084e6add1b35015bce5839713122da59e880cffb567a5156ead72f614e14e5abb113b2f51286aa8d1dee1e97e0b9091bb119a336bf884fe54edde862669f849a72d339418a1ab07b15eefae30a264316f8fac8c5f77620e81d03d5347bd15829d0627ad92281991b3123767903ea0421730da7871835e23d195a0efaa561ea9fda54fb882f321e9aa34a25d011c6d1bea0334f6a6ae0e64709f7f5cc3a03ee559d315dfbc309f2ceb36f3310524898b635734746de6cdb2ca0257711438fdae7b92a6a2ecf25cc2ff97984c0d922d6efb8eb65a17dc83180d921a76fc1fd6c952121805e694bfbd02d367cc7a2e97fe6d0a44a907f532d9cf6d78e5772e0d17256095c049f7fa98efc43acde21eeee145c2d752b5e1b18a9a3cda5cf258e08f42466bec017ccb04ff53c7bc2938b8ea65e7f406b4f297768df397f16885a25c3939e60ed4dfbea3469f742947972a5a86e6e6181112b84a5c30e7e5f311ea5df13f74682bb1d18976fab88b74efe00946b6461eedd379fba61b9aca1e7b42163d58d76d9a3fafe5dead95819cad07c270e1878aed0b1f962bf76ef63a7fff02f0d26a59980e6ed0289a72fa6950e89023e5b64c3ea3d119c489c7c710cea94d79e784e7fbdfdf31da49cb0752f47cb7d6ac3af918eb6ac61cbf9d2f9b42aaea43e2b47c168020b766e133f177efd8425062dd52a676fbd9e146729cdac138cf23a15363c033b4aff31bfd1813c14b9bc2896d8377e41a36b58ebf6841435c88100f42d9e28739bb779ed7aa6340f1f06f287cde229928e94f1416d22b2aaf69be51a7ba014f63366b709daa9b8cfcfcb511a084dcae3424d0c37e39cd8808ddc8e115c42ab2612cd2c07a7f829b9adf904d817edb11813636a656795b0123551e92b8789740d433d6df4b274ec010fc8700c0a97c0fa58ca1c231bdcd7e0f533c9f91c3313e4d4db42269eb811fc22d9ff408d3268d6174288e28e82d94956aaaab79062c4f3269bfccfdd93fb7c2fa44710b824adc09d43e70d8413658670a07175b302be3fff4a795bf0cb41cc34ac7a21ae3dca4241bb8192e4fa61a93072b177be012db6afd7f380ec724b06c8c0c477979e0d4d41495daca0755887ac98c04339c876b0c46aec853d1faf2841f5137aac6fd81f3820163af5318130b8d50fbb0fc2404e335c521f9c0d8a0797ce14043825dadb482a895f80bb56a2427756fd726f3f745a7833fb6601b81fc5b0b3ef457dbe76170f32e00c30e4fb2afaa0ebc7ed48acb1547bb09ecf009f303123fb9a97ebc39c66505e36f859c5f97925a73b64901ecd7429432aa6f200d7c5e1deeddd418e49148fb9baf448f69abfe2a742a90b709b60940f5a5ed18f2724e09208f63d39c5da5599ff66ff618e2a82bfed6d46a7baa04781fced7f0a534;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb403c6664fbf8a2266dc38c47cb677b3d613994ab0d06a322aea26f8b960d0983809bdf47954f02f30a18c9e4eb56a2c530dbca66f73dbd844625d516e4f6a15748be87dedc0f8e02574339e948e624592f7efbc6aefb0009780cb11476e438ad182a86d4824eb0e5710d1a88febf912e4564a73c24b5e0ef9a13f9e59b67c2a1dbe02cea1d5545539f529df4baf07373fb469fff994af88a1bd334a4846c75120a1c8e5520ccd76bb44f79fdeff41085238f9ae1e2822c37faa43a6b2124c6a7f778ee453d619705ba82f9a22674e6a82ec381b30f1e8de59133d8428324bdb492a095585bb2a02ec922c5921295a481b75ea5ec2e570ccf0d989a1bcb3de4fefb6ef7de28a5a94d9ba248aa2e19da1e8d9f6dfec0e697070fa6653395546656a0fc9241dbe14bef23739f7c79337aad8baa44c2a2c6671b9d5cd6cc5374bf02ad8f378e4fc81818b4eeaa3baf201b90ee91a64be12baa3e33fb779730b5ffc3ff9b8e705b17adab8bbe52bdb1636ed1351d4c76faba8af75c30c513c71cdd17f2f9da6f1c775206701e0e1f3794c9ff47b08cb795cab6bbb5a6f854a0992f5fcc30517134f059ddad95214cc73fe18733b2448300d03d8b5a76a83076493f146530e2f7f920e2fb9a30e069257340e89d5ade93d07b7ed8a40e80dabce6ab3237c96e88a4fafe665886736c961627ae9be91ade41e4d43de05f0c115be49500bf806b58ec9c66b1abe473055b60ed194aaad422b84549fec88b2bf19904cc4807b805ced695735103e5e0517d7d18207ae795a122436700417c49b43cf96fb103b3f1362ee418de87929ec5290a6ad6dc1da08614a929c6c97fe974b8e4b6698765aab7e26f1fccb069548904e855cc6d1e1b255db88d13ec443500bcbb10cb45cd363be217004c78a56a2c1e838aa2cd1729450790e8a5e4cf68c27dfd860d71983c6eb7d40dee25dc3a099b1273aa05b8327a836fb11d6b9d5f2285f4f7505cf384cf2519dc8ecbcad54dfd355e9ad55bb44df9edbccb484a59b0394b996c193325f8db4eaadd77956fd0b04cad8ec297e56c89571039df59ad708dfbd628b15884df38a5845a2a6612bf7db0bf2498d85cefc94db802a94feba71ac14de0a88f3edf23e2caa0cc33bf3518acec2d427dace503f06e7ed2c7250f02fbb3dcfbe4f0b84de96f2993233cb72033c854d1e04e4cc1ad5c2252d61db636ed1971a7a1b8241b1bed4ee2fa9a912c5d3df4df137fdb572d8930f29c71bbdf5f663a3eb4376e5b73f37c228f97a33d3533da58e38898e003da8457f0c4e3dd46b465c15bbd34b8653ecb5d7f7fd5cc2eb9bda801091cefdd0540af577d5e0fd811224e1200ddd48f7db86dcf1e4c3a1944ac2e71047b975c8cc215194e223a9e12de4a9daa4a3ebf500807ca40eace42ee9a22a767c37c37cdb1d741718c5dc8112;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf9f0d4171331be9c34517e9aafb8c8f01b31ae429a90e9415ea5558904897f6aa8106c6f3b1cacd9e3a12d9b4b2254e7de3c5eb88db2ed0c41c2c2e213ab2e215ed88a6b3fcad9593d0fa4d4355e05a3d1f86f4c8cf0da0aab9a38fa06df85894897f17483ea5b0628643bbcb174a27f542399bf04e1fd2c4fc0a233460b2622544826205c4863002ecaa7f07592da01849c6c93410cff677167871e6a5a34735c0433eb3dd3e4ca4f253c3a9045efe701c1a8d0aee03e6a6447ff84c4b79335d3eb2e0330bc9d60954747475de679521d2e8252c08f522000a129d7d9130db45920b70bc5d6fcd682312853414a54aaefb16743bf9f85367ddfcb616b5a3876667e28c2c2fcefd2441571a60284ff4dbda8269baf99c69cc4b0d1b161e9c00ab42821ff98efdfce77f640d1dea5060d7ba097cd49f8b6fa57bb85fcfe16c8c4a6b1a7e92d4322c73be35d705f13cd28a2ae23ba0f8a9e9dcce5a9505b71d7364774e6f26775212994a26bb641945883cb7b0c0d47ced7ebc13c4c02b2a3deef627ec0d56be3cda04b76c8a35c3fff217ef5150b3cff48780d58ad4af678b9f1741175bdc9823e40e6cc84f23a20ecfc13eea1e39cfe0131c00759bbc0a493c00ee587f9aa16e1f3b2ed3e691af15707793b216ecf2a302a7e5f64826a720712a7414471bc009c3bd141a01d36dc22134760a515cf883d25375b133d768a8d2ee85ae97b13b0a6eb51fb8ed0ec919f61e01e4e70e10f6acdd7a9ac8bebd476fced6c92ac4ad402463735185053c37a7edf54c37618d6d0f3e0ccba4e143d95d24e0129a7024364d7cc9173bee6fe5403ae473ce788701ef7bc4c11e97567a20516f54c20f812fb12aa8ef6c2c42958f9cbe8b4a4900a8c21b635f0ba5e79a35e561c2c043c3df2a05ace0890038edbd84e271fca0aff9faf701e27daece975a52140489565c7b7632e907ff60ac1d475dd6e2f0fd374003dc4baa639825f5cb79d93af692c61a01f18644eff7a85d10dce66ab712db3685e84ecb7570fd206fc06b9ea6594e2591dec9f94d462d77bd5551560b34d490e18d077e37ae6ce185b866118b37ce3b664279d40c83e07405089179c5b6f26f7714926a7d083778e6ebe8a2b7b8ec316392515ce69fe029770ab514a043f01560e5a5964cf5d362994b887696a7bf9afe2df84bdc3c2711cd295de9580994673fc0f4fa48ddf684d4d7eee1dcca993e67a31895f1ae720cc2ed6ad73b939c4c8f2f66572a6b3b9413e2de1e49f552cb2d72fc020b7ffd1c491a83ab0892c3df9382f5150f98a33c7875a38a33d1168a1596dd48f30176bc76c4f2a8fb06ff73b2c5f72b28183b32feeb2c9e11e8795cec0981cfd22b2979854bea817b6e92ab57923c5bb5c01904f53f9bb6f70dcbc2b2afea851f2d56f5ce835f6f3af47e25dc74fda3e5b9463be7f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hb6fcae99de9774894617d831e7a47f3170da6928dd8fe522d1a4acd235a1b3a36146552f883c861c90589bf937142f897449367fd27ce1d229abea020c99a256bc337da867d72a4bb12cc7d0671fd1dbee4dd8b64820eda48183722a036473283d394b17c39a2a13478804e7a888e7b60f3a440666949f0d41fd7b727fd1a47bbbee3e1368b72c9db72f6213c227fab3bfd5ed3ded543e793bc9d4b79c887190e3000b7eaf133d3f5fbdd0c2d79859d1620bd82a3a6cb3d22e015c7ca629aab7ef3449b1162910a4f6a457b41fc93f93e896ed516e867f6b22895d28fecc96e05141d017e2b485d9dfe122bd39a2db9b5e3a98865d2ea50cf345dcfc04a0cd0f1ebbd9b11c85b5eab74fb275bcd12f841cbda182e2b1b51cdf4aea7221735d60d7feb78f3a08a98434a7468e175aea176830ec27b98eb0cc8f9f2da0e6144206db66e869ce2022525b3a4f7770180d3627966eef63feab25f903e462fbc3d95bbee4dc04dabbfc3df5925162820c99e267ba9b64484a3797e6e6d24029fed565ce768b7a253658336714e0c734dadd024dbc030240ff343f220b87a8f6a468500940c109ba2f809992d65fa6ea541853789216e8ef3ff4e3942400092e228b9f60ff54c1ac5f30022ddfa78edde89ea01795e4543f95664588613d43eecaa48c12429f6ddbcb3f8d7d9ac63d20819b48c2b6c8e1963485f85a2f226c736b5f92f84e871b8d5c67af400ec95f4b1412d321138dea6a952249bdf4aa76d49c6d6d48955d96cf44c0ad62a3a02314cd630d0daf8dffb2a27ed40ed71d04f2cf5288018c78e365ca43cc67196f6a1c63a0b47fa379635e56687d8ed3de6c0aea1912d9f2f509c9e8d15bb2de1b816652c5b05cf0c259a1a0edf0005a77a49a09f5ebd135bb0e66515db3eeb019bcbb85d70a2f94f294db057130edc53be688a279c147488b75897bc2db36044e621927cafce30bcf2b272ee61519aa0b7343394a4c52c3266608afc157c97c8c4a9fb2149b66f72b02ec9b07edee5b86141ce091837a52c728adcd188e4a2e5894261a248b370682799d7ddeb12e62c337084667d76f8f82ab7abd7e638c2cd8d37c8c155770402bc5e1129bab8ef0541b96c23d9e03c07bae792ec18622fccf6f15c6faf50e7d521d07455be01a704762f62a277a5f7bb834a722f87f6833841a23eb1cb6c06e229755f28e72a4f142e898ed65e1b76d40a504673cb303b07ce9cd5eb0f091f0d91fc913976613792405332e6f27fc9444a9e12413c64b8050b44a4a2636a0d6f1e942c85617010766b7a72e2f0533a7dce1b59d3b5d89774754bb3bfac7b8d61fc507fe3518205adad9d1f6f12f7a4c06c80d951daaae255e3f032d3f4d57e3bfb5364ded5199f6a78a08134f3da343a9cdc7490f0e2c1524cd610f48f1c5e7bac6e7f8acb2f1eb7bd734d4010;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'ha158474fb634795db60f4cd3fadf480d30397a70574f42877f5bcb3943583275885c6cc6ab0afc00fa175271ffafa8b7226eeb2bed6a89adee425074791709d8db6137210b024eaa1de622d98d8e9786899bfc1ea29ab81d79ca821315653d63b709764cc919360797c4d090aceb88d680b53e43c583ba33ba0e98cd67420c34339aff25187d2a8d73ce8a58da3996ca0ee57adf00110f8675e1db245357e382686ab3975257d4f011ed77ab45914e4d49b42b9ad9615abb6df9fb3847430005ea8cf598dfe1ab1e2589d507236bbeb88f450f7840741d0676894c817304b3439940e29f52db93c9fc529087cf8631135d133ce4e52e6dc07ddcac0c59d4cc6fbc77896668d2e2cb084b9009487e746bf8d793f55a5ebe91cfe9358aa05b8ff8ba98ee68f8d162f93c076ac8c87d3f214dc17f1b0de0038fe636622dbd90a7dadcf548bf7f143a81047c1823860f29eeb69f88e1c25c10a2d557e168177ad5ebe520aec0d477f7ca0cce665e6d8d4e1ea113923b78e114d4f9bf7708c8c58b949be55a6262d3b29d4564d70a870603850ba85a29173c993e46faec42d4768ef20d38df662cb3d3f50d8bae514e6c27d1b33b11b69d7ef92cad25fdd34f57254ef15165c98348f9c74db472a477589eef9a5993bf7cf5f8397e53803f975dc8fb45cb92c694dbabe8198259068c091083d1fe5241c7b8ab6f6ca9d9a53fcd4ceff1ba932c659b4f4264439e39c57f3e47086b2fcf938f59e680a1f64c08cba54a7fef37cc9eefa4e9411817e07c78d17961dfc99b2ff3dc45d75d6ff1313a45c95350442684e066352c410c8ffd42a57b1be218f3e8944b3e8e481d303c394e38d0c4bedad68a8229d7b64f363ba9e1a2c955f664f3d8cc2cb6db348834e7f35fe6de3b1d4d0a10da92f2e0319e7bb90879020b63dd027535333d7b32d0ad8b38d184f3de2c0b5184023f5143a6b84f69b2daa89247ded099ad08efed18850862a8df93360a83fba4f8ed4d18f09c6396ac58dc32588a5c62e08d4c84611734384a9fa5375674677aff97a21a1a8f5dfbc82f823963e7828b13632c78fc15e1027263c1abf944e48634a016091876d5a65a8cf36420f0e78fd8da378dcae636518cf7aef54cbe44897dfff187cd4595b04be3d68e83a98c6a7890ba27850f16cacba1315002f0e3e3d64e44ba4b706586e313271fd46612eb7e1e2961d8de2ca30869dabf9f662421054617321fb7a60943260810181a32dfc985aa67ae32bbdb33e6189759c2547ba18d07f576393e9ebee7bb6c96e150a7a69818898a4ac2e72d8042400a836f6d6fcdb841e2d5b90575eb51eee1e71de36feef249908deeaceaa1422a59c07653276d5bb2a3a0526ed2a48a795ed786c80398f9f3f1569970571d4fcede67dc58a3a2da692dcca52eb7a701244ee4ac9105fc5ca46d4f1dd2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hf1cd3807bd3b575e09ffc70fa8b5a2a7cf3c262a771267c7f01a0b1d9317791617c68b0b542417c76870cd4723866ef7b89ea765e77929a56c413b58792823fe275845c7145da1ee935cdb984ea192f1e58a78576a59a8345199a4c7e1d16b6ce5dddae159b8a614ccd8d88343248c7a0bd98b497154cd0c3834843ddd125a2bec34f776245a3606bfcfdb07e438933f57c23f683c55c7b0960234106b7296bb0d0785ba82f84e540b917cfbe253389d4de01b780d850f0184424b07665a700c245ba607b026cf4fca1340f744d93b370bac42d5fc62da9de10ad42c8b962c5ead03a0b7cf1ead14ab03833da387547393fc1c4a04058976bb22dd2889d5445146cb6c0ffe6d265ea29c43676435c28aaf596e7677c130ca69615f8fdd89a06e2ec5feafb61d7d3ee7a9dfc4ae99b0a0d48005db4ed87f6308613a3af7cb00349329baf4c3947822b121f1357be79b9b6caaf652679de8183ec1588974eb61c10d4bc10d5f7ee5bf12063e5a7f38bcdd415f94e619ac21ddbca6a8b0c8c13e5e129125bb8be139882cdf85a3c06476b91915d127277f2935ca3b808a7141e000e3f73fa4ee20f745cfaeb14b55746aac730abb6b1b6b644f5b7e847df21bcf26b35b6850a277f9b107661972e7c011fb6e4871512565fc614b6000ff04999a84c01e5fba4f0a8016c16d8539bec00c80c7a75027d1b1bdfaa585365535a9e3dc58776fe32d8126cd34399671d8934efca1436ce4c08678be736fd9a94bf1e1f358094d0261fa3338688a03b338b8dfb106fc0f29c789f6520e8b8f39169a3425a21572835e749c4467bcf930bbc3de763187c4afc088ce99f42e6117b8856f37edc7e928e4a7cb4058dc9f426c636e1b2354f26f6e9069ba7415ed2272effce9f0ce0a90b12d0ca9dda5c624aa0554cd0ff0d911a547557037c4f69e315dcbb16976f55ce637192d00ccf4ca764b26e250cd520c90c2ea843f2100fc209acb3f5de7e59729b28c5c34403cbeb21bb8da52a02f08c19ac66ff2eaa5f19d840089d7e70943c51fdd0a8a711eb4e9579d1a119b8f82dd29caa87b5764b88bb98002fe3caa7841ecccfed39df40c8aac068028d0842628d1cf113e874e9dee34519ce49d151357ea47a4eae1f59af1daee2c044e17d4e26a04025c4661a4bf5deebfe2f31a3535bf108256c7824cc1c8991480709287749e088227be6d374638eaddbea50f17790d78c0aef0aed0d75fe0193c045ce1a5d1dae1557be0cd8eee608924733ebb75decde35da792ee097e0ed729519374f18e5c6cce4f053f53e50065c5de0715a89d655d64cbc30d3e500bd8b3e76929a9f777294d76a5e98ceba59ce19e7e18deb595517ef97ad7afd03cb772d2b23401d0c6cdce8eb4856b12f2247daa953e904bd41f20e812438f2415ff772deb76aeb5aecd91daf988c851f8b5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hfb5feb032293fb05d6ca405197d5529ea00746ba8911c4fedad2ef58cafff5da79cd3e47ec51922c2ea4a2796e82a74e3b1f44a5f3ca047b6f643a131130e3297a7921d7b680fe5d8b925276799421f44cfb827c7d572617af53757368e184b9a4abcf057f53a1af97560b53a8453ac9fccac68a4fd4ff1b6088d641840ad7bb713c80c02d110fbb235b8cbd4ac74a196e5e40bbc4942537790baa1ddd75685709a39a2da57cc649fbafea64bf337dbceeca0d5696d534858c69ab8dd8136c9ad644c2059bc2a551bc700d28731634e5ac2fb07f7f730d464753c658d2448be244f55cecaf2d841ff565d7a06d1645f2e4759519c6348df2a64c43c58e117d0962b12f5ca20727add9e1911a8f33e1feb4550920842763cbc77021daa3c2bf5ad974e5be454c33205dac21e69b925e076cc4f9364cf2b6ed45a0b2b0374e6c5bcd6367feb26b3cbc130cbb2d3fd38c2ac8763325e5e0f04713aa9aaead6335292cb665bb6c57b35abc5fcf34a9f1005b295f808b635954127608512f9c821d5c84fafabc28ed2c1bb0f57a46afe4fdab8e115552ac61cf549ea7679610018c3428793918c92f820bd6cd5b1abab6ee965baf6a28813c141e730d310aac11b424ce5fd7aa66de136ceb7cf7acdb07e864e99bc3f0164b476f9205d89c1de5c106a0d700b6eccdc070192cd0857bed7c45f28bb625ec0d9b09a3aee6af907fe888a43d79d8c17c0fd5d122e126bc8e5918076ffcf108a501c61cee68baf17e26973f50f3d3206c7a79186c0a2ed1fba8be02af353da72c2697424b1ef284e5da3d90587621ac00c9453a5fc289c6539f2f79867a9a32d38d90152227f158d74bb5d060790c1053a3d8eca96cb52cf453d4a1facf681bcc407a57e7d78aadd6a1825f0cd0942274819ce58d77226a63690a1e2703d007f97f298d62c123b1e9cab448451090ff62a01ae5e1a8674be4e573386af39a7be38ed9a58919149d341b1abb4e776b262ecc0242bfbd2937c97915323595b4a12a4580960921697b0f90b3aac3955a8c06a59b29cae0f1aa3f7794e231af3fe34c7e9256614c4cb220cca30fb9b4dff4884a3b057b83a960a1b25922bbcf389e3b87d496c929971e98ae302ac324ca829baeb29650347aa95116636c99a4b824a563f790d5e5f62a63ecccd83317d2144c2852d5e210cf5ab042e7b461cb779f44ba8fc5ee89eaf058431017c767410ee40c9b3586f67d245b7a148a8c85be263c1af6db81b36b5a030e55463e960060ebb0958366b8421879949df0ac69f29d9dbaface517978da76246e46c6e95f314fa3c461b7ab3e8cd179b62f4ab50f5f5f95037fc352447d482e95f8f7d00e64ab34a5717eb9762f30e9e1a3ff2e02e863cc188f43d4afde1224b87da81a1c9385b3875a5e81ed19f1ddfb3c85c99f0e92b38c51cf89b4e8c5e1aa;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'hc338ad2ef28316ec2a613e6de6e6b92237fdf8913998f85968e673e9e5edab8dd2cbb866930f8f32b61bc204e30526823f05dfe16315fb107b9a972dc9c70c68783831544ff986fed3dc64ecf6aa9976e5b50df7863c74aa82231d2577c52cf4b46d6503a816ca371b05d55eca4e81b91ffdd1fe478cc1ce405ee8cc5f0d13e06d9d3415fac95e1d97aa135070d783455ae6def9bd748d97baedd74cbd51538b3821010c79955ccc94088a6b0985e7843300393779f615ab2680eca8c6f366d5a587657c606023138eef8319f44fc289182225174a8dd08dd82dab4b60b0d26173e071676c53daf2dd2d5480ed521533f6b49ed7aaef6f777f9742d2473a9bee402a0b724ec754ca752896e3feaeeb4e2976f11a6e2435d41f0340ab351e97813c5d5595042bba56acafa372c84744b5794551a08121ecc2561e4074ae9c14f435aea92e35a174770675a7d6fd283aeb33beb46177da5a30f36c9e962c2be757c32451e282c8939b0d69be1640eae216bcf3ac8cd81bc79a6b3785d9d35ef411d8f57e5a803a016fbd54669d02610617dc9b25df5cbbc37348f3ccecb2af861cd042410fb27e8759bcb6c443b14ae115b6563dcc2588a615de0df8423fde9b68476ec7f6d125dcd7124abdfaa1afe60e3ec8dcbc727181eed52ca8d00ddd2fa824ce2d9e806fb86ac49014b6ece1a104678f7b3a509f3bcdf84c23fe8eb2d3644891bff542cab0ba0cb59f28f8f411c75f7f6ed70a75405d01c94815874b339bbda6fb95b810e42c69ac2ad848d9a3047689e92d5aec6dae4680e3069155d89093067302d5b22dffdaa1222e8a0c08c274b8b02936fa86d57952e5a454b023783798329f84701ff88ad5c6c27a4dabde6c9c8c54d6a58813c7ce052cfa9dcfa3c4e9c942c0dd9de03127b28ddf544bee477e3fab59f72b33d2e22a725e98196386df06deeabcf8d0cf74f4f0bb81015ccd2cbde558a0e7d45d7a3fcf60f1a2fe155e57a4eabad49bb14dc260ca739c458745b70f2a279a9d6866b2977795fda0ea76cbb0d00a30fe67fe7b85ee78896ebe8f0696cbe1ca1916e4d9c2b2a7e2a28c1a8b700f500c397675ad909c13726e3dfdbe00195dfd1769967c6d4947d72d49a645fdc44f1c44c15c96c403c6fbb775b6cf3273fb9cb1e696f49e76575fdcf6baa3c1c5e0951dc7dcf47ac5495ee059e3fad7973627afaad0a0713df80ef954104b1bc6308a33187dec59b276ebe2f74a4305f57a80b5d8db1a0de21973caf9d2e2e484dfe3ad9144d00ca8a7d68adce47ca4c77b41b2a9a229303ce08e893fc9fd5879c3962c45bba63994daca37a6e6a29bc3057a129222951c188a3fa14e54a73862691980f062162fe7bfb7fec1a3b2bbc24fba5313e9b41033c932b73057e94f2ec4be70f3c182af294eb68d84caaa7055945ebd69cf919058c38412;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h80c11a7beac1588393d453ba029b1b92824253129a6fb0cd83d24dd656d8997e377746583df3cde6a250005b8841f41a00041c4ce02869786fe64386252df3a2d17b790ec7a938425bee254fe514edf246710b7f78ef747b192dab55b2bb3c6eb6d7a2412371a48bec173a0b1b5eecd4f5aa68b0b5f73ca718c8b0fb72b61ce32a6fb9891e4918399bbc6f03f5f1cf985058e8edbd3d5e363d2c5802ef38be82e7448a8870301f539f5bec7f68329a53922a0fa79ce6f72f377816b00d66751b329daaf1d4b54c08bf9943c7ea40ac97ddbcfb4bdb0990a7fdb8aa3f9306a7d6cb864bd50d1bfd91504800f4dc19b3622aaa18599c888e4e362f39bc61e1b35efae3e852e256225e1423e6a32be23da74b6ac9a9a6d5e2294b2b6b34c7b9d39ba27fc1935fe168a83eb6342b32d2755e8cc074bc09cc209b035e8687673ca5ddb0419fd21cc7f40820cda6b0dbf29643e3fa2f3bd657f62a068e8544a754bb31d3dc93918db2771080a7b2182b40c4a1c5e27b0c6163e30fb14251ba42d4ed81a01d23417103adcd806de83fcf572dae59a8e2a84d9503f1f4d2a81a1d7a76f55a6a85ec203e26a36c3a2afc9366750b6326022b377fdf4b71cc947e264d930b07e80704e1a8bfce798fea8e26044c40cfd24c2e2856aec535c7709214a2c8ad8e37c006837e9bcc64b35a6cd42c54299f572acab8e696df77600d37d1185f095f66aa7bb6b035b0bcc1a1a396b1ff617ad2c22af2a0accb226cf09b13b3e45d3ca8ca0dd1067f793eda5b717111ec083ea6525b508242cbfccd451d35b5fe651ca3ee54258358263bfc74fc7c61f26d4c58c4fe72415d0eb51a621a816f5cef1c2f712b8ca2a4d58ec1eb6d0b7d025584e69260864e34f5d1c586cd48d484b600875d4c561c8e80c2c81cd74fd622efadf4b41bb1f62541affc242d8eeb8837937b8cfeb3ad6c08004d248cb18f6fb3cd2355a5f8e586414a757dc45cf1987ff90aa3dbda82000d961b14d0eab0feb0d6269484391b639a79fae67dfd5a78ea51151437b27474c2edb6159f0670169c9d89cc00111c2fff5d6675eee064358a02ddba73e9030d02f40fd6f5eca3836243ee68b07772333a0b8d753a6d5db92198ffcc8dc7b6f89a97c511a1361a22aec8ab57c967272deb0ecf0db7779f691bb094d30c0406562304c34357df43c89f77bc46ff248834c51d1ab38bbed45203007aa8b4edde539a4edd18e0800c5264176cb3e62995607266bf4b4ec3e0665f0b59b6666a406cd024872ccffdd4fe1f1af277629a61030e6b19deacb8cb4c1d7f2046ae505d4a6e0dd216f7597834ace9d623a1a4cfdf0310c046bbe89f7e421e60d9444875d6bd3534e66ee91da7923652a757c70ee1fc7c7f7603352abda5a9877316a53146c61ef6a16848ec45f817bcde38a38dc1c035026dc95c53b636;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h996164754dd415bdfac9514e5a01e2bdfafe1d093ce478572c536047402bda55567e4ab8b64ac3849f713a6a9e47f003b98508d3d4b79b4cdd6571a1ef3fc7b1744534d48e53e34f2d6794a071d3c6d10d6bfa9f8158a0598a795953d73bd7474755250d68ee90adadbb3b63d5857d297989346eb0c1cb0d76a3b46ef6405d7c0c5b25b0f3939df7c2b6a3b9a3d8e8ecf2028273b8963897e1699e024a2cdc4738cd42505ebc79e1ee65f0968537da10b925055e90d68992b5058471d5d7e6654f9f72d6250031313eea65e732de7316426e9d539e1fa61b51cfcf9f6eaea5796e839bef80646692eba344491d0e183c784f51535120006b01844b8beb525608758e87ee4445296587599ee54774f0d84601b1751786609b558c2c107eef5fb2f395a57333fa2884e8ae0a9fdac3f051f7dae85ef3ac660280334d457dde51f02fa9f56fbf81711dc2af5c0bc57dfb80f7fcd33a8f9b41bb215e7a13832516bf3aac230e9f3c7d39dd375cba73377b40961358ee244ee35e7e31a17d6e3aa7ad9e75abc3e11026d105d6e0f96fa04530079cf86287b66e8a46cc4fb3d7344712150da36174284e6d28c45e0bdee28244e374b3603a6f8b6664908be6d1b48564055b65dfd30f46e20f619a0d25381782c81d18d751e9308e38e7d4a32fff31b1ac358a9f5f16b3a64964ed2bfb04835e719a3bff0d73898c44ae1f69a0cba01e738ca027d21a4772150f257b195ed5fdce3ee9b01ffe6fc1f1139439cd414bddb7369ab1b148b45aa6ab07f456ed055c67fe66508324b8b1218f396bd1c358c26885e89f73007c1b90d886fdc8eb2c667e7c3309f1fa5ba854cdd01b95c8f8fb7025df8a268d8bdde87ff8f27f80b0e833efd7ccc6b165c08cc64ed04d3b642563aa7b3bcd31dce870b3f5d62628a461cbd8ac8ae3bcbc520775265751fcaa4d479086e47d90338ea40315be398629b996404cfdf49829cde91c513b2b4ce6e111dd8321856aa71918b72a0ea6305db627d2f5893273c19066e4a194f0085564533c4f1757c576a9f9295f0b09b1f1a7a6573ffc924eccace71509cbcbcda034922b1d5af0f076c2ea3188e1cc9469018e99f81b5fc4c12347b185f11ee65a11bc66c07926946a625b50e52185393e50707fb1c264b43a63a547bae0fcc35e728da5bc74adc2f0022f7f23ceb9c5a6da4fd60f00db73d377342a0d9f8efe0e21f1f901c90f3b0e35bcdc60c964b6d6e113b978f78ec3a563e755be564d016886cee48956a9c104ff6cca16ba98efc40e2e07439ea6c9ce073f8b82048c6cdab15486a493eb67d2553c6d2d512bce0ed82d768a94b4fe96700738b4fbb41f4652443a3ffdb9eb080a70aa8736020e3a84eeae4e579fb5c35ac9cb8fb5b94190e9827afed47d29bf22f84d062fc2e6e63d43b22fe57d09938d966531fc6d9d0038;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h2db8c75e211aac446fae2b961602f9d5fd435e3248820f354d16506630272691a7e62079fe1cabefdce0146de6f23e325a7a2012775ad2e2d141a1aab1b6d20a5010606416c5a723251ff9b90473ccec0e223ec4fa102825319f559cd01eb389f320ebe09376f360c5f47080f4754f577cfff720386b53bed1a18475dd3458903895626d6fea224cd8631b3e862f1c2eefa4a30a4dc79d1449bfa962d1678bd99154c7d33ae796e370d8a3db2ef24f7ab32fdbeb09060e1be0ff339dec0f99d695719938a1824a1a1a39161bd9f8525302583fd19b407e7560f000c11623c2a1516762e0388d6e8784bf59e757e9b4dd43faaf5e495cadd9d2f12937f10f2b4e261d98292da74e2871eed2bd9f7606ebab4c9cd9e35851313fd081ae644a71711fee92c563a49534f94903ce926fe67024b01534489aa78cd60e357d1ca9e4a68c4d39a39840586b5366af8d7f0ecc9fb8b2cf331c7b7be20e4574b0acd5b8cf9c7fe238b5345ddb157b7283f308f1c12ed7fa67f7d0d2694ce569a218ed0ab19e73726f239fe121966dcd4461caa266936088c9df6a91917cd2005504b3c788aa8d3907694c48f418617117069ae906b4dbadc4f8e85158374dfe4f8de0f7b3e82fba58ef6ffd6b1ae1fa206b8115033f1c5ea5826aee6c8bdbcd4021c65dd3a58505b8ba70460c6beca8aeec7b54352fe8c9b24ad5b4a314fe6aee2739695d89c273eea88ac030079008c663b881f1498a46592c6b5dfe72e79294d59b2209b96cb20f82b77fde5cb7c35ade20f867e4dbcb4594d8fe48b21bc9d107748ba0f3be5d3687a407ee20cd39a042f8a778184e4975f83ab56bbb9f480925d163483801c397f144fcb0b2262f71a6ef42810213796f801972986a6f69a84dfba995128acbfe892cee7707171574695c36a871706438a00bb74b3c6a925c2ed31687b71c322058d039fc45e6bef6a5da2383f298450a56daa21e88756e798a046faac95b723dacc5d29fe029f12e714aa80a15ba11829193118a759d94c28e0833da9928878eb5c2937da6d439eda5c991ef5adf97a8c3c0cb06ad3c9964f39c4adae29c6d23a7dfd7df8a3fe8f59b4831cd193de1325aa0430dbb05d55a17609c0e69a3f424c19e30f069f81b32c89f5bf0729a5e2731b2c2a7667089e66823e3df7c9a6e72a9cdfd12e35a216b0ac8499d2b261a50ef022ac90a2a919e02e069ebc87f9607b0a88aec4afa238ebbc95413910609281d4e3d3c9cf55a0ef4261ce97b21b6d50b1f19a3a367d271da4d94dc92593554afc5e471059e38f9ec55cfda401b38f48398478047ddc4b915a42cc6b4284424cdda48c64bcee792380866c5446194a90f8c1e6b3b1dd3d7eb54af0c3b4a85e849fd2b8d4455d242eef757c209c6f9ff3a655f8e89570b26c709925c57a0a062c6b96385340be5c5fdf84ab;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h30cc8d83eae848fc48d48672aea3711f08aac0f7a866824714ba8217a70d9621cc53758a6640c656f2bbfdd5942dcd18f079d5d427d2a6cdcb84311207996b209dc8b36d060480f0120e3c059343ae28040b1d9053394b73afa047722f589f1090cc414b6ea59ebacb297c681e26f4d369a6e8ceee75ecdd985bee2fee15dfd272d16ac69d27c8089044499760103043ea256e16d2b9caeba48cd79596372e4935de7529eaa6510c9f51a2383a3f0b7d3037c1ed392a64d30874ef9602eb1f81c810723da09e5e482b280f221ec873701e8278ed1196546046fbe3b0f4f40278eb8431e0608dbc42c35f81cf4666afc341a01d9cd525d46bd769d1bb414a1f766ca20b4fd16c4276f12a375d2bc019745cde8f662b9fc7ced55169f1987fc5ad0e8723d96639b1ddd8fa5936762008a1c966de062ecbd0360adfa85401abb539ddf402e2805413d0e215ba9b231fe1a5088fda1adbdc3bba5dd095449e44844c0ae5b6dc2904b654d0793879d814ea4deb146f3eda322a0f3c2df1574f62c0225105988a92472253da9ae4aefdd83726eee2066417f2fe7b0a5e23517b7e51386362f45da79ee8c3d654925255127d058a8cfdd84e54369bf714e2886a568b3e860464d47b8d919e7a68c0e853feeb873c6fc6eea08dc291fa1d228f4b9ff421a2b9d800192e39e895069f405475e6f48269533c9367a8fd98d03dbeb2952bd4cc7510be53224dfa07bed3c4129a5432e323474ff42ec8a64374dd249ff16c61c709c929b14f11fafdeb4c69c249d9c1bcc0183d1dffa72d4878ac5945b5b2c26bfe2bd8d49396a8aa601be1ad2e0eccbed8a1ffee6418a8a4f3fd899983161b17ec439c480b111dd51f4faf854a0e2a63363fa732ab182e87bbfc8ee6f0dea609c18df57cdac081dd7aa45f101f3912c45db6a1c8c63ea92e6ec452f63668b40268018df0609861f0b216d0497f4d95268706bd9900bf2880f543e4a10c884b56c4a1020daae86bacd399f497b25f9740c065381cc17cd8c81125fda84b34363cf03cf43860408c0987faf3effb1261dac31913e915c3820f13717cda3178ae8a300f25a32f24ab8fee1fed2b0248f211f5b9f55a55b47b776fcce1564c130f8a852ea694a939c642ebe1597e4c01b155c773c93a2fb54027f2c0f46cc53a2c703ab5c991f153492e8c13d2d4a46572f921459cae7d2bf3c0ad4bd29742613347491327aaa4a5d9ef3271633df08b90c8e59cd67cefd45b7c54e4005541faa713f1001a9d1bbf0e47b33c0bfde9f43d386fd0f5f0a945e049212fb2c032b6c886d110405e15aeda933d3a45e29ad1421562c61a308741fd07fc88eca69d7fd5e116b445f1def1c202f03df6ae709ba2d006779856c8e0223a9eeb3d333481ecd732f66d11c769bed9a8e27350ec48dc169b69cb73baef4a2718fc222528b7e9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h76c43a6e833c1c2bcf55ced1dc072b5d1f46682e0779dfbbf625923a80e91ae23fb7a2637d9752425e6e405041d6bae659a000dff23c03503a95e16194740daaa1531ad05bc8569a5f6eae768de689cff21eeb8b3a3808230171564b7d326b8b181525b43f52e2e805dd33c8e89f3ffe78828de4cb2ac4d0e7c897bde8b7f038c03525512204a85c966248d60cc9a86baf1599cc2f25a5e71b7c0db691587122c6ad030b6915d3a8cca09e3ac8ab4276a25702e1655abb0637bc39200df6ab0a043c855d99637eb09b284b461035cfc3dd39317549bd9585fddfa2a8ea409889f13e43172c50cfa41b2bf50dd715a4b3fe379e83ab030aa24cbcb0ca76ed53b702012572d0b09b885a8e939c7c0ffb8cce1349364d7db91b97fab00b84e0dfbad30dac49b2dff5882be33793664e2704d2eaa8c1c2dcf44e8a3c7532f5fb5810accea18df1c63cebbde1160d882b05eaac8d585cca7ce44992f5cc0d1dab6bf043d326883d1f1dc88521ac7b40461e0816daecdac3a0fac6ca660db99fd08bcda58156482322f00f1432cbd3dddb87dc3d6a64c4cabc94590c875b80027737439b19c80f5bc729009d49044e95bff0c238fbf6eb3e9fc2f411790f969bbb17c011b68e20c893e926bbf1de4ab538ea4ae752f1f61528228bea9b3d98e7bb107514b6c67fd7b38b61876d9886a0ee2d76505c3cf0276b618a044c9a15dcaf8f69ee2fabd7b8f308472f31505698903a07f32e1be186b2c2e35aaaf088aa9d7e53fec6247949a0363a8908539a4ea1bc33f041b39526f4edd4a1000049ebbefc3e5fb74f8eccd26d4357b295fede59ab2135a49937e545ecf39765cac0159438d10784c7bbd4c171a78d1144c2af9d772c6fb3937ca04f5de9da2d233aadc5fd0a3897b69e7e7ba07a55bdf5946cd1d86fdd753f063993641dfa3455dad83defb4cecded02559c9df38dcff8d879f24f2a6fe60bd2cf8225cd82256da15ddcd596a23858b89c6b9c43705a373cc26d1adc6e2775ef34215c7397126f29620caa58c547dd49746ac0f27c392a01d8b674cfad00bd98a4623deca107f6ca4be645a06bb779a7f6bf1fa90c66c97ebd0e5b1ac8baf476a3a85dab670dcdf313bdd7068088e9730c7a2c538b7c6c7c7881eca184da66418bd174305430c3e6eaf2a3c2ba666bf9c1edbd986f6033a5c5509c9b1dc289c65c668807bcb57af532f353ea7e8a2a0a14ec4299d0537bce94e25cbb468eca50ee9fae715945dbebea41188943832e222371aa93656e6237f649b9ff133ffebe392c6fa027789b896b48f691eb0ead02569b5aa3fe6ea448bcf0124c7c105cd76f3c2a2980c1b48580d3a5876fc830ff3fb7ce992ba8674f569a631b10f8ac680c7298bc79230d7b9552b1487e78bdfa40e8caa5ef99ba091300e30fbfb20f682f83612d3b58f9e491ff9bc9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h701fb614e494dfe6e4ffb6f039362b2528cb4b123af84ba58fe87ee01e568a614f6788d2df2b9b8dda4a6b82876705903214a21f33b7545728e8937d68d7e00d9e3b2be6541e15bc7eb47b4d966f706d93a716c2d0c8f65431c5f3c34ee80c7882f60a48b9c9ed69e3290b01558d45e52510845ade8860400c1171fbe6457fb3ead9d65217d7a20387ddd61fcd5f9c611b62cce426cd579792c9da3f865ece9dd4401f037bad862b28226d0b7083390cc5daefb47d59b295d1704d648c9b287bec15fca38f1eea88148d306b1bd386db8ec357bca73774cafe8de7d87a295deddc9ff29d443a23734f8213b1ba4bbdc34eccd380c451d37f63ff078fac579c0f0c5fafa48410bab8b5bbcf63b194019ba20b362b45a9ad7edbba05b31cfa611e0c75beb25387b30121f1a41a5c12dcb08234c34181fb50c0df2662945be89103b36e393de28fb37819e47a9a88102e33de5de131b370954ef4636fd9752fb2763058172672c9fc90112c830b2e128c251cd313a79bdf1d832f6d29b8e2f70845ccccee604f44d3da026c8fe7fc344523f5077e6e5bb8d8145f8c46cd2f601a0dde4b46869db12d0ebd245cca51ca99f809d79b39be0eb333bd27de81d6f7fb906b2c9e0ee0b9d24db77af49a09fd6f5aaa4dcb4ef3064a216cdb6c60007c112edd1f761192a8c8ce14cd4b74a2fd076b8413b74b8334233171476e8b3ff41352a7d634c4d0c4719b3370d0fb000a35bd82ff5384314575aa29d3646bd5786f23c8290fde9eab3103035bd6d33396e826e861d6f79ed48d9e67b3a412935d70a3d23201a1fe2a2e35941b6ffc30c14222643cc8905c93e79fdf22ecd97bbd3f8949556aca391b9eea8aff6b88a6c7a9bc95d7a83f762c02eaf2c04bffb1df497924df0a5030f10befb366a3d54541fd25d3fec1b735b68184888fa1ac0864bfe481cc2d41c0394fa0f09006aee0d5f92935c0b809daeb3a16d95de9fb547f7cb3c95a960d91d143e7132e341c6e86af74e41f993566b0fe5c002c26f1e4a1b99b078d3f22669a549ee27029d4eaf7dff2312675ad99a38b9123d3db79bc8f05e1fed0e876c73510fd47b4db6b2e47faf7e76ea2efa3ff0ede70ae7e5e372e95b7a9ca4b23fbcfdaa93008d72e14f513a9c6f9e8aa4d68ba3e5e09263b4daf3af2639b80b16cb461dfa8937fe7c4089f88f7c116591b6b5c628f4390be1d5d5576565b0b29376e6ebf28dd03ddef8c949d7781144b94db9c08f6794b7854dd5ca69974e9d347bb39d3696395c715e329252035f0280f8b59717fa6b822be32d4524aba240c43a96e4c3ef63bf31567478b19b8f16402db4a0c67e5392efaf6127fb38e0919885dcfad53823e8bc523f232c09b8891b47d634e25a250c6377f8aa43f68592044ba369fae1d1f0f56780cfde565c0fedee6e4fc4acc73c916155e0f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h7bb0adee4e6f7ee2951aa6ecf3d3d4028f4d90c96c6716a56343a99774bf2dc166d249a1b2c73a68ccb1dbee25669a5e63ab61f8089386592141d6ee0297fcf0159737ba12017c395864f5775a201ab7b6b83f66bce54ed70bf437e5e4fd021afdc435698ad2d49e15fb44a4a9db8c814a9806cb8a9a67f8cfa3ca45fc207a837028382a93dc042bc4c250378f432c84d121c69ceff084c641613c1a2a4b6baa904ad25de125b4a4934d66290ff64b52d0c052d88518f4378f5dd92cd092f1c40b26f925a6a9d6bb05276d68462bb2b682b85924f942c2eba03326b639fb26e21a46033b6568f8e309d2ba4a5ddeed26cb356ebfb6bd9522b0352b6b565c8d85f7255a2b5ef61c9c92643799c01f553cdbb35220b06a9b0564e1da6c02f2d61fc99fa02a44a8c8c2f92dc7d442f723d5056cc30867287a890806a9d8c88587806e49ea9c57e379fc5bef5195ef496096bf4e48139176ff4bf173150ff05578e80c258d2ce42f5f73221a643e87a40455bce3ddc7b22c9c16bd34279452c61bb43c77d631a023dca63e2349cc2f369450e71cc7ab6c9e45fc95b3fe273136ed6545c43bf3add978537d44040f1793e4799fd1fdd5464d181a3f9301e0665934e1743ec9ca87e4b81e7ace848670edbda3c3f99f1524e54b700711f9eeedfb9f2a64037a3831e91aef9bf2aba41275224aa60a3485008573063630cdb573b20d6a9d3345f7c58bac353dcbb2fce4721b2aeb9703baa1f029c709b294c00e66a26b30e00e592d3d84e51d83972ac556b7b46dd5308f0341faf745e0c5950477789e9680b889fa95c638ddabab6d9a152dad2d66ffdb72c43db1c113dce035f8967cd934dc61affa9b99cf141603cc5b7517a1a296698baeccb54d909f3d58d02ea5bf4a07603702e8d86a0807ace88ed79486a6fa077612a878abd401faee921dfa7c2a06a06712697335f6f05a45426e539fe3b5f49e12b135b35c1c7224c689db982cb2344dddf317f23bdeb03c1024ad2d213ebdf1c54846dc4b3c0203c774353eb414c2be9cb9ccf83e939e602fcbb6cca70af531e243068f1b5823f0178d51bf441113e88844dadf6b230ca05c969f10faacb5c9d0f860b156057a80fd9b0b678211023f0413c1638fd8078b3d97b49336d3145786e218e82cfbb5ea00ba5ac56063eca32bc12ff66ef710cb5030a9f5c0c3cb3f782c7fceee447dcd07c1c5b281ad3ec4347d461796a46f1c66475b29d878a4391c4ab5004e4791af2d6ca7d86bb1dbaac78bb3a7c7868b43818b05108038dadf1bd897ff5733215851353c65842298f56959b4cab31c3e14b3d5373126da5d00190bbd8c16517a89f3d4be6a2d43b82349961dc15e01b7307ffff2519016f92dfe49345a8027c67a7aac55bb90654dc395c5b7c0a2da576d39ccc9457c2e606abb696570bcb84acd6efe46;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 8192'h4790bcc6735cabc1e34fc04a05dd5963ec9bfcba22bac98792d5e896e2eb214f02f2c2710154f650e81cacdc67bc60ae1560bed89eeea138ecc7393ff11550c649db0411f5f45a97e63872363b5966d91ebf257e50d3fd0aaa2579259bfa60a17c6817d291a9ae2deedb8367a0337eae95773c7009931d3acfe13361b11561ea87ea30e43ed5f132aa258b0511c2039ad53949e5adc9a0a792e7223e5924e5cea74194dd6360fb312201c459e4cc365fbf2c94a485a2c7d1f19dc1927c663f3f6e4e365f0b3e7d5b3c30550dcb205c0f2a40f06ef8b975e1dd9dcbdc3f7b0b28f8825173d9c52adbe6d7cb6228d0770e9080d9feabb19cff259b5d4799139d616bd2f85493db1dd7b3dcdcccf518159d11afb9bc9ca69a822aa2a37868a1f80e98bc5cc79330e29e1c3eefb3024342a36d7869096e789acc194b7ef37872d3ef7c90b36ffbb4eebaf7ee96cfd8c6599aae89dfe0391cf6ae79d7a0cc931e6268624d388b48c280c71f941d293e41bfa153fac6fd280cdeb4bad87c136aeeb660c697b3d1a056641a99d15a99b09c04e4756b8e6500385cabcd03b2ead35bba6c1dd934e5f9f9deacad4468e2b6aec246e6b24bbf46e69ee53a51f1f9c472cb296ba074fbf318df1fa69e7900bce32829a3f5153dd90c9135fdefccb930dfe6b7e4c1941b6c7d0a223d3a8499e207ddee29d2250a6afffd1a70d035697ffefd5105ec572af87402fc5ce097cf7a0ef3f98d6ac25cd3c8f76e3fe44b98ff41e386d6983fe6189827c25b8c3c495f8f76911ae9cbef1a27d099f220f09fb4a6fb5896b8291dfd09ffd0ba4a4bb3e58f3ee7612e6b8770bdf9011b4585b5c6a6ce635fb3ae69498745f4706b99a1def1bd7f59246056fbf3709ca670799c4d17a37b63b15637ad04144bb3b49b1fca0f6a5cedaf482d7bf011086362e93e79e0a7238cf07c5d40daac66fe4a5053ddd34d52aeb8342cceb6cc4d77188ca92ba640b19bac8a36b91d2a835329696793de3e06fcd08caff6841b14a0e1bbb06e7d310ab2b54022b82a712a44af5a4726a74a39f53dab7d69b18fcd8b45cdfc1b4dc15266b8d816eeecd981db55a242a43a058b152f0cbe4d82a00a9dd6c347923eabad994c4bc90f258928f7d39dbdf8beff3a07906c3a875e4866f04261841d18f1ce783e6ffb98a34169827ac060f9f171bb0feed00ac484c6a98bb63b80cda85b8ca7cc3b894e9a9a25f24b5aa2ebb4079622a9d8bffcc0ad1a50aff3033275bced70e4e48fea1c5abe47059b7c0162b0a25c63cd42a7b34c47a43e3f6c4029b3499b4c4f33f3702c2e716b1726f0e95b765c5a3abc60b0c908139a97c3a6cb3f62dcf02dc67628c0a702b52b64cbe00683743f368fa77cde09d37ace765263528e2996bbd46bf9c4d48d436ba300503c3c4b1eaa679652b5bf7588ca5806f9493a;
        #1
        $finish();
    end
endmodule
