module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [8:0] src8;
    reg [9:0] src9;
    reg [10:0] src10;
    reg [11:0] src11;
    reg [12:0] src12;
    reg [13:0] src13;
    reg [14:0] src14;
    reg [15:0] src15;
    reg [16:0] src16;
    reg [17:0] src17;
    reg [18:0] src18;
    reg [19:0] src19;
    reg [20:0] src20;
    reg [21:0] src21;
    reg [22:0] src22;
    reg [23:0] src23;
    reg [24:0] src24;
    reg [25:0] src25;
    reg [26:0] src26;
    reg [27:0] src27;
    reg [28:0] src28;
    reg [29:0] src29;
    reg [28:0] src30;
    reg [27:0] src31;
    reg [26:0] src32;
    reg [25:0] src33;
    reg [24:0] src34;
    reg [23:0] src35;
    reg [22:0] src36;
    reg [21:0] src37;
    reg [20:0] src38;
    reg [19:0] src39;
    reg [18:0] src40;
    reg [17:0] src41;
    reg [16:0] src42;
    reg [15:0] src43;
    reg [14:0] src44;
    reg [13:0] src45;
    reg [12:0] src46;
    reg [11:0] src47;
    reg [10:0] src48;
    reg [9:0] src49;
    reg [8:0] src50;
    reg [7:0] src51;
    reg [6:0] src52;
    reg [5:0] src53;
    reg [4:0] src54;
    reg [3:0] src55;
    reg [2:0] src56;
    reg [1:0] src57;
    reg [0:0] src58;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [59:0] srcsum;
    wire [59:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3])<<55) + ((src56[0] + src56[1] + src56[2])<<56) + ((src57[0] + src57[1])<<57) + ((src58[0])<<58);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1050854e8f0bd6080ef901dc8be5babba880bb47916f2d90594432b7d76facfcb86d34e4c6c4bddb1ed6de7d35a0dc435000ae6fc9489362eb73b34648d0fd0694138e06f6435762e442726143470e4592905a9ed35cafef45725601dc5e5cee995a72b940ca46a3b14fa1b47f9e68443;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24c3f86366fdfed2f1842b7c054a053e49640c3b7f7aa6733be09cd2d8c8f895733adcb91e10ca40be7af93c1a146f5c49b1a3e593a8ce76752efdae84e461d1fb1b1041e103f45bdc5756044255c6a8706dc9198e24b9a433d350eb1858ac60860b0945c0250f393f6d083d8dd8d3612;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5fb05616d522f1324d28cffe95a43df6a3d96e6d3a789b056bc4f2ffe38b7a5583fb9b5fd1042afaa452cedb4c6602c24fdbf27154c7aaf9bbe938a70af3bebb5afa0add553e089afa469a21d9cc46d49aa6f09bd29aade9fc1610935928469f9be2fdbf212be7e8ef3ea46771d8e9bab;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h521b462d401c2bd7667e890342a09061a2b6363da49aed43a56b64a4ab7a005b54c0f1ec5157e81264ca65bd9b724cd754dc660bb8903949179b53e59407f8f18a6e036705a219108664036206c3c6af1af209e32f90d7777d7d296b8d0a43d565117a8c3f78771a8128fa004c5135ae4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h310a70f3a9d1d76b4a54bfd2a109bf56f80b4a016e69fb571cee5834acbc0f4fb40665bf54ac82cbe8da0f2eea4da697101cf46682de1b8b884e101bd522ed00fb8a189f453c3682a7969b41215a3142c895acd6dafe26ae38fa77f922ebe9f91931ed63ab9b0060f601dfbc984ad32e6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32866b2c70b4d3d5c7e667dd900589a21198b3a9076b3283ebe98304b4fc85b18304fa01859e2825c00d6078444cc88fab705c14ced92f569fbeeadad678eacf59f403a7b76672ff3d882f4e5beee26c1911ddc5ed570210d22229138a5d014dbdf54f92ba44ce51a25d27be1e7621af0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h317f6e2ea4e436e07d194120c320282fc7236859ee9106c19fc1237ff4278493cc94342a62d4695d05553472a6b8020438f619799b12965b3a4b06610ad844e839575bf4895e9da33005ce42636c00bbb03ca10697653fd3b111c8826511f68f30d9de31ba37a99d95ffe6bd5e04d0ae1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha51357c8df8cac8670d7a11dcbb0dc796772d42ddc41daffc2c950f55fdce0e01be0a6f6afb583529805166b4c7b2a8c9ea4a4c031796cc5e9b97cfe3b40f57be8779146f6ae1cbc33614a08ce7b517336d1cb225a4e64568865e029ad2d570714c4e0e82f6002ddd001da7616588f0d6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha48ab7d26f63c3ed77f81e4c5d9482b2365d999867c85f4385195d459e7a46c56a1eca21af8ca2be056fa50cb2f7a0904fd2466e2b85637b676e1a064ac2009dba54ed3deacb83f9a67d4f6c4f5dd9bbdfb6623e8ab1b3f54ff66151ca9af2a3ff77153b4972bc466ac9d864ba5bdb558;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f63317271c337a10e1f9cff22b32f6b5e8dede445b54bd521512225cb437bb4d20eecaf681df33ada9635ac432a7f3fecf07bada0ea39c0c12d2e4d7dd83d8e3b1561d2e0f06795bb5caf67c812734c59a648c4c658b1459ad19573a3fa76b9c58049abd8af859e6e407cc7324015991;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h371065cb7626e63744432c6a5c964168bb73b1a2c1b70ff44af3f20bf983fde2d03d5d25bb4e28fbc0f823eae88cc7da9e3d035bbd1396e9790ca65e8318e3b3084a18d9907d5e81d69577c82ff6728b733777ea40fbf8a2f62d2f429133274a419d84c58fe4421f170121ababaca7476;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he588137d68502586bde617638cbe22413f025210b39d9f68026910cc57d74310cdbd20a4ef2281ae3364d6cab8adcb0a3e940d0b1772180f072a1a04f94d86f18c2ef6a228c4cc86edb059c434820bd69956059dd0c0e45869ff4c7584010c588fa446885f9026871b3c078c38689a9cb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h673070bfae22824050d7090e9709a8a7ae8016c07bb81f941883a0c4a696597e6d0e76119f04c202623590d7a42858dd81dff607d9ec3d02f29a2b4160ebd4cbd3d4ec602e00b6573396a405b23ed37973d940bd887061ea8bcd716875d73152ff6e7077f478a9da522baa9cf84b3178c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he4cf253febbb7f9ab6e84c8daad5397ace7f54e21f0c4fc312405e9b4ef506188bf411952e65986231d232c8bffe6e13a82ec472c4e4af46afadba679ae102816760bebc42df3e90b424ef94b4fd33cf51859d883872694c328b136631029079818f1f816a82fbd239bda0c86631f0d85;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4291e04222a4582faa5c05c69fd523a34fcab01bd73783b9c6bd2bc26482576a870ddbb5e566a0d37d9908c7147a04dd465041d3ce2495ef761d020983e38bb724f9dfb1206a1382ed1d04bf54bf1839af66448a45f575c9a6f3196623a01517145eb319ce7d7b09003057eef39ad0893;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44673eb5c65eb90f30aa657a117f7ab45decfa929e0944dd59b9885b388a9a4c7fdd600dfa886d2ad832c9100908d78b8984bffee97643a4d00ee000e0232faf60cb824c3421587def331e5849fa8fd36c10981afb78e94df3d547c6478e7fe308327d9cce4317d5144005cfe42fc4b5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5311901b8ca912dcac590bfc445a4e2a51072e6cf17be4ae9b580e9a3fbd49328161db303d28a35b2b3f374ebe3a185a19da643956641c06df8336d8a002e7131be6e4328f504bd829957a47d823ec49c0008dd6cd717f45f9b6585bf7c1b1a5be141326b1ab9c6ace78e1d8716d88f84;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h723693eecef7509fd0d3e9c1ead253f67c01f78824cb9fe56de5ee5182e137c18e3151b5f7577f0d3bf9fc9e1f4d8e76ddfc98138290338fc62b6ecb575e10747836211c9109024f21e33b3d132da97069329ced279ebcf02ac75e41e1fd6596e6c3a6f883a2eadbd68aad21779dce034;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98c8d5b6358798dbca773886d90b591fd5f17a3f767374add78d6d608e488432fee65d8f1386d43823c591bcaaacdbdb49b9a73f12f4408bf1e03feea0d67fb4cc1ecf812ac573ce830446b528167737eedf03409982676c8c56e6f588c38ef375a2b004ff027c549b0d9e7f118cb61cf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf2682904f55cf56a0f717136ca4a60ac1aa961aa6e081b3aec0754b5fb41d7bb0aa2bc235548780a1cdb924bee66341bbdd45f129d2cfdda417815fab120123dbd603d0ee741146c8fe0c477128e030d7fe7adf1d4d343f97715b5333de2bdc41c32ce552464f7749d3549d03a376962;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9aec0697ae3359a8709f9426758b585d27bf1a4a928d25b978963eaea60b19b21ad7b23c2ad2d9c91a31420c4bad3d92d3d753d0a29e1d98a3324d458f86be2c99a12a6e1cb6f3b968653ffdcacf60346e147be3adc34406de1860a0b19688bf75f6bf41e2de0d79ce139da3016a2cfc7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hede10fec023fd6adf9a652ba698f572ba58f24399bb9ed6210a4663b3e60f29697ce35bfc57298521e31fd1d9ec2acb43c76ece27d279d7d073775a506c9f0becabb0b962d05bca2ce576a2dc8fb83e9145cf744a9b631de7e0b763ce2d262c0e28251377491c5267beab645bdf1034ef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h556744e3680dffd0011a524e10959d72f868a49aaa8a1ac6fbc921c61d59d84e884a089dea5ad0cb81e009f17f631c19ff31a9f18924259ce9d66428c5f401aac9a642d01e1f531298fe3a2ed604c6143c45a406645898cc7e2b738975bfb2206087d427e39aa923fcbd239ab1bfd1127;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb75d8f5d1285dcf825c28e1dc4360d5441d066a764888f004b4b8f8a12104c00a41cff8a184bd5591b9fd29c123a3299163c2dabcf4fbcc44c21b31fcefe30a1f8784cc29028f554a70a9a24e087820221a37a0c9b561213a15746c1f6186d0bcc81bebf72e89c6943950855d66e99e3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b6fcc0f8d647e2dac388be01b5a86036e7a5bfe4e1b28e6097c763d31997080d995fda31249c4e9bbf3c2075c3c33d059fea72a456c25cee7855e24bc2149660c6fee4100cfefe2d2cfcf99882430a87ee2ba09e6d5177250ed7b0f143b53a0ccdda4f3061ad11510ed9684422b7e2a0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha176563c2f4b264e2108d3b128e2de4fe6d70dcb6ccc0ef057f36c9385e8b2a730c9abd6e5c91a209e0d10ca06cc36b626c6e8400961d880690cc05d25ed2dbaf8ab0d807b2061374f2bb324b8680ae2a371a94cf44bd9cda8d53edc879ad91e0ad128fa38383bb258b841d7a6dccb0f6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he25da74e073a4faed80bd3aeb720d1c5ef81d140ae1db941b36733d79d58bb666aff4a53da26fa572cafc9d0324972e879f2639e5584228a70b4cd2ca1a08540f1c17aa57676fb8e8b199534162ec7245fea783c03dceb6feb368c7da7bb514b4434492b0e82dff0bd73332877a681b41;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f9fd35d761bebc9e10ae68c1e9279f1e23debb13e07616e504605d357f1734cd902967bbaa5f70409659db4c2c9573e1206a86d8d694cfa6a4b587d29939942aa2813dfdef300eeb208a2eb221018eaf3d7e24d2c48124631219154b12ffc3a753671e0dbfa51aafdaad8ecb24108632;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h867b36af076ff971ecd15e57d37a4102260cc9a7edec03f4928252b3e72234c022b3ba33bc8ed9921481be272b78fd2e5b98cd4cb7d2bcc04b7e1cf7819f13da7928e86dd5a4512b699d140b560ad67d8907f4275dede0de7f4ab9a0bc75066168ef7b94c59e64c7787a498678e69fd11;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf86b2a2abefbe0e5d36151beb33db770d8adfbeaf437ab491961e50646b777c2fb4c02797f059fec82192bd6cc32b7bd9eb0831eadf1c9628c78fc2942101f0e7b34738d33d015c135dfd5cdd0d92f8400805db1f8d9ecceaca065ffbcf25b21c16f27e1d0adf54d5638817d91e90eb45;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c053e9985bdafd1993e1f51de0aa2c699b8e7e888eb0046c5d49ad3e3404c2f2279527eac4b80961bdc3e1b1ac110b8b97423d61848a0d654828cf9c617578a8c0dda1d54932c6e708a5baa10f190c18d8bb69de5c5218612dabaf4409f87a1548f95a855df33b964407cf78d57487ea;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha64572635cfce0c5aea1c91f75ed332c098feb9bc2e5f90389ee985818b8f7e623a26c84901cfc80f15f459aace5a6758f96aef34d928d4f5873bf0e2c4e968f527fe451230eab90dbc564c02d933832ed5310490c50ff2e40f3b5ccda45713ce61011ed87259917f7c6e057895b4e629;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2bb9d2049a2295d96289eae4c0f99617bff8484fa00bbf1232789f0815a46076c4ed11ae97b7e2ef58385ff59cac5710846629b8e73e998bdab9a63363afd108e4ee407246698a97273009809c2ea289e4035ef8a36edb5be3c505f8fc252856691dd722d0f914c2fd9a3be06febef9d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84d2baac77c3b9368872b1b4f44436490f3cbfaa0ba72dab47b0244df4ba8f6136f761850d822e37b6da5100f738be8f056d30259b67d01f2926c56f37efe6817837c65b94a1a9467c961d06ab0481abefed139511b803e9ffe7c3b7f240008da5842fd6e0ba116e73d93d14deff349ce;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heed2d41552a2b544e38f5fd266d51f878dae4976f443fb0edf3d4c65fa094984b4995fe711488782b1bd764f5e6520315861fff833306498bfbbc1f2b8ab4d95e413094556f1165650348888d67ab356d2406cf8ba98bcae3a6f89b25a1de2f62637d09101c4c7af58f702ab73ce0809d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h913407fd638060a6ee03d98411b983ede30ef8c318917b993492d78e465c06015c06b03105ee4412d126019ac865c47967f86c3f137d93c8ce67765c01a5b0f3578e2eec22935631de9604932c65d59dfcd7c66b886a71fa22a3c6c3f7ce5c4bbdd1e23d9328da87b924a91ad311e96f6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb8dd4d1ad3092ecf540cb98cbad3537f06c5c6d0045412c1443634eafbbc1e7e5944ea821e732c68b5c29559a5ba545e07a77bac4d37d432defae8f5afb0ada0c95c70e8f6f55a8f5a75edff5e7d085399467eea24bf82e4e89e2cad4eb71e848e93adcbd48c369a1f2d883ee92c8be29;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h19775f37f1ade095900d9c32cd4489347d16b7b7a3102a080b7557dca3e2aeb05de38572e6aa608713e712d25af0940ef390e829906cd6ff9689761b3f05cd97639010c28ba382ca2d4a79fe09431c17e36d2c884e2009cfd11c5143556158e596024dc67eb6a1547d070bb765c123dc0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf0a4b01f4b5cf8b5f8e5978ea9d332225b0c39841feef36d1f1e1d2c47635dbff522a8030b5e1beae4f17fbafc776c3ada894f2629e5c44b502a8e2fe368b5924b70501edf2821142f99c9cf52b9da0040a29a33ef98583fbca30b70f8c8ee92ae33a221eb5f8e87394e7c4035316d7e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c3eb0254864c7b25456ff0a5db96453215c436c971abbbc290c29c804f99fd7b9fdff15b28201ab2faade63970fa44149842b052e75a56a65dd406a61a29f347f2e05b5e6247354d35a2039172442620556478b9713eee6c4d6d721bfb382cfc9e456d89585b6fd6a1a1b1095dae5bf4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e960b8bef447f1327670dffe507016bb540cba31688e3eee1f2ddbdd69f876d74b7c6f1d6d4a85ce0308049f61c133d3478726128558c024987482dcfb6ff2a80b0df9070aff5b6d3d49729cfc5bcc2bc54556d94d2429f6448052a45c26647021a1758206725cf03dc37afff35972a2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32a69e114c25cb470abe58caef926458d5fa3077fb8d520326e6ec95ebfb32e485f8cc0f4ccc195da42cd96204e3897d11911aa9b46c9b45b5b70a9e648cc0c3a6541664051ff0900abff0b6546279f592a9f3146f7f7bb0993e3dc56f50849acb4b6ce6447d16ccf60f9ea60f0a41869;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc71e69c729d761a0f4b067bef508a6819ad45ff36d6623be208e60d996952adc7a18bed0debd30141ef8537ede5591ff605bf22e23d1c5be983253fab69183b838a349cdb7f948e0c99bd912b4e0e8d3be2474e606a6f429c6685f17e8eef61ff4ae9e381519b0baab85a26555d503994;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9d0f835111047115dbe5ee1bf45153467d32dd4dddb9af10193a49422bc030ba1c46e72b51d43cbb292958afd06b5636f5b82b2cc3cba3a487c019cb6569a901ea1bcee190e3cdfc22fcb61c7c582ac2b87b375dc91ea491e801177960df7166ed933c833e4afa1a752ee02e1764ec8a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha15b3c4563f3e55eba2542983eab8309218723bb6610d3b3d18f387a62f9887b072632009fccdbf23274b7fa7863d68c106b84681694e349f1928e7aa145e6c8c3d77ba9c3391a65aa25ea43a965ba43c963794c655326e14dad42ed0b92375c54e15be7c3ba90d2b35a72ad6eda343a7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b93fa3e72f269193e44f942a7ca5aff6f78ee7328e556c3f210c2ade2764104b198bb7b7ed0473debe30db0d99a3c788cb6b04216d12580231fe843380159830fb4f57609c14e87e1811d7f75f4b6c2f133bc83b68d2462b277be0b2ad42654be13443e8cc15bf8e7edb2f9bf4bae0c7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd54cdef116b9284c56fd9458c6fea7b4d5a04ae5ace5a07ad47e43f1bf80b092d397feb31effa2f5f7c475a45ccf6efd242961fe6695d76c610e43d09b9636f387b845c69eb5cc16682362274fa4e3f3a78b3f04b1eddfe53ffc4fa9be17485004a74824636e82b4a4f22574289022cf3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3d15467dfc2ec7daccd91cc2c2c26b2ebb07bba961e53e598f5021ea545400fae6d3effd265c62c45a0de073dcc5871dfd556774ca8aefc3ef41d10e6ea88d9abd26aa9603a8dfcd6e86568c832a6d5df9bb62c013ba9c5080c0073d919b4cb4c83f6a520796f2afec329be1fea81406;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb304085893ac8c8cfabe536301a84e02019dcf4e22d5d0ec3de63ddc7d105d568c453ad5e97dc621f42b9755b816d5af94e7328bbcce2843653775b1a22273e68c32a523ee80d60ed79b92699937eed99539cba3e4c07e3bfee6fea1bb1ccb92a2efd1b4cb80e56bbb3e3e36cb4657ec;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4659516f79ba80fc3d1c9de4e69bf24702078ffe7285922fc8a793a33d42584e3b1ca68f3f1593241e52559f514e3fb10ea7b3eb9c8497993999851908d4fe5f16be3862416cacfe2e1707abb3df69b41af842ce7441f01d722d5854cfb3070376ba86ad42d2f72c9ab9d752a368a9b2f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h67e00809873c7f425d1db05519bc33f16ff99d3ee47dffe8159c71260595e66158858b60e21e77418e7c786eaef0ecc3f3abf36c9c08e32b3569eaed93fef7387fa4800ce533909f9c9586785f856c9bf327a6a96ed4c61861747a3d3fc901f9edf70758dc2562184eae6c8f8e69ed024;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1bf92e0d00a50fe6e89bf0e603bae286757f3fd5104d162e6c7bb52fc1467fedb06f8b5f33fd15e14f3d9b0287bece7c88ac06e2b2f9e93e4c54240163dac5967fae3cdf4d0f1bd2b22c5acd0e8760edf54c3cc4bd05fab66ceb10e9e3c305ee8b0882c1f8d7f16e16f33be0e2ea11844;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf531d75ec0631d9e6488f253e0f97b354c98b07d84909b746554f17dfebfee21a96f715b387d4dc93189feef78691b3019c22a791f89d38b1d176777a4e4a73a1e93ac10b282d879de4c372891b600e38c4eb605de508c89eb6edbe881cdf676c98fc0f3cbb58c64483857a154eff50f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h63fd24792ff0e0366639ac1c3c0a30164074da29ba5d64ae32ae68a18527f8116c4ffb7170d0a375dc0ecf5d3756a49555f187c57aff0864fb3a7ca661cbf323aee65ee91268f5c3a6fe622d9a03c7f754843dc59c030c44b97fff6af5af41e67c073c604f84efccf43ed8a21eb6d053;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34c37532400fb508dd10459e22554f06249828271d704590fc7a86ab2dea2851ea33d223652098610a04194a75e0ff1c8ad4d7b11e0cf8e9b9edd1a07bcd56b0bb93c8cce983286b2850c2e031294e0bad649e14d459fb6b5c7aa4fbc25760b5a7534f1c8d0208041545847fd544a1f37;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd934dde3066deb93c568aed855582fdb607c176f1c1734d2243bc8528a9ba0824aa8a1ecd6c9b4c58a8c2b076525dba23968801b12aa94fb903147b250bccdd2d917b998b1e7097a4f00d2c4e49557ad88c1044c562169c40f1cbeb05dee32c5522102fb43a2c3acc57d0f4716b396c4a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a90eb12625bd1f797491884f1eda634a1e63198944769c5e41bdcf2378e3caabfb15d7d27d60543044e29c5c9177e406ce3f4335a89b48f66a6d0e75369996f3b63f1a505e78cd1af887e1b547c57ce91cbd9d76013f94f255492f14b6b9ced612fcf59056e2a26c175e274725e88b1c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcdc327d8a811784e814efbec2cb7e8c62b02e8f855e862ece03c05912fc4afc9930b62470e6b712a5b5c4d5ec427112149b4efca400bf26dccb83597d0fad9513dc8c0b0d092fb687ce2a1d1e54a31e1854228a23b6d585306e0acc8a7599d6b2af79410b2512ba900b69731df9f18a51;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6146c72b3369a141850ad21a3a2896fbe035febcfab27f73deb49a49256f628a58e5935ddb2984210c0e5d513dee8439a864444ab08c5d61803b1e8e9447b43b12dc5f10bafbc9c5721f0fad1e72950b11a03882fcab5a802ea79a971f1d343738ea777b3c8550f2b4215c5d44b4f611c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc46f4a71e49063fc35317f0c9e8ce8fcba067266bd1ec3f47af78e8f6a3fc1e6d8e9dab385908508966f52eaf67f2167738f7eeb7ae9d5e08bf21933888d64de2a226e16dad32bce2793eb38e41cff677b13dc54c0e6c44f63733baeab2d44286469fae73e7317ceeddb6c41f7852be02;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab20553199dd47f0517794adf37306bf111fbfddf8d454c131fad67c10622daca9d00ad78f0d6d7eba96fad6fb4a58f1d1ab0ecd43472ee5524ff84be832436a9854754428832e79077e2b4985543c114c0c2c8a666e0ec11653236171f77903dce390b10bb5c7bbbe1fcdf8841a7dfd2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f71c9b32e84c98815c8ff2caa5d9bc0973f29c44d22ebf47350f929187cfd94f6c265471e61248a91c857640455063b3f979e9e97d9068e728a3cf2b20cfcd7b006fbff2248aece66faea01e7ea8e6831ac8de1374fef8c7f5fb0fcc72ebe94a1d5c984786b7acb7fa099258ee3dbd9e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd6559368cc09ebbfdf738288a13727489818eed62d45b62f8ee7af3e8cb0504b691c981090091442fdee6d8563594541ab4d91d6fa8cb212d5480423afe401d22de2d439a8a54812ae140d5bd419ebd52e53cbc6a1fa85986520339f612642fea61dcb04f7937a6e85d243e58c94cc4a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc9817d4500dad5597dca18b636b58acb8bfbbdf142eaee9cafb44dd1c4be4d156c3746ae2fccc5c41cacd83ba7aa0fd93c4d1b5597d30159c2c33c225fea31b064bdba5292cd147c03cc1d5383cb5ae3598376602f9e27febac2d751f1a221fc2dcc1775d192206ab09e9fe32cf73059c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ef5855797039c49c7da85c88b91815ae312a8270976ee0b93b04d55c88586b0ce1d80069e079e980e8d277bf24821e79bdd7ecee51b3c802c18920fa42e36431e218644cf982b9043c66276906f900fa4c53326452b8fdca47ea3b41cb0ed21e1a62a4258df44cd976bf4bb81a2b1132;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f7d19d7886986514d006b312135af0a415beaf0285c67408a7c434b5bd7706edc5b95003595d6b4da88bbd77b5efba0e7ff4b39749f6bdfa0b0982018dbc4baed1c09667217223424461e4c4b83ac2ec58c9fcabfbe8531090537cd6aa6af604456c4f087e29687d3f2dedcddeeba01a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8610fa33d84f2538cdaaea1a6284fb22ea4a1559b46fd3dc14358aed8d92d7669cc337953e09e575f12a8b3fcbeefa7f5149d778b727a18754e8440a83f4755c36055d6cbc13f14b6eacad6dd50c006499367f6439f7cd80418ba9a8db8b60979ffb0abc8f1d03604715eb611f17d67a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb8de0b045d2a74454f46b94f75809677c6bdee72dfbe51a82c6e7c3e236ffcacb6ba2ea0f9b72cecfa55b36639b58157c077b9645e83d4143df0e3478fef407c97e7492265c9ac723b5992e14354d5438cb5b44e8aa65c75dad17249be75422f3e1dc1c0de93446f9cef39afab64b1710;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47bb2e62cdba8668524ea30791cb38adadd5a6d401cc772f0fddcad0d0b642d28fb72c83d186a756246b42b278f5b3646f690fcf18224a5c9c5ca712c859b63bf06571f78640dceccb2afe74ca8d26773c8fbcd1bae180053f38305b488106c432237d2473b02fa770b9d652cc08e94bc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25b911fed259ee7ce9694627f53287945e42d645a3c7a8bbc50dfb2b42e9eae0ab52b26aeab0543c3c4918b0fa486a73964bec44e55cfe7b8fdada9c6f78e532ead87cc38a4260c8b810c40199bd9ceac723e9249d9ac8108d40cf19912f266f936fac25fbf918ff6b56d81a44890f160;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17ecc103bf451bc7d1a0180f655db537c6b0eb2bf4c32484c77f276df7ae5a68afce30b380263f6486c6291eedd821624d046b8c4006bcd93d4bbf96064bd6daeffef0b9640c459893b3d4592db75bdae1cfe810a6471fd38f7e4d0c9d37ec041d215cfeee2150f6c0de05f04a18ca48b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h577cf222bb62729b0171e85615c25f5a52b89e1c11a8611b49b07dbed1219e4ec3235abf9992cfaecfff2e5f0a3c464b0f754c4cdae95bcb20edfd629a49266449454171388425422eb93bc2cbdcbbf51fdb30f0fb4f4e7f4fa14ffd4d46659e747d88386f139b3db93e031e46e951b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd00b7e4cf75d390f0652c0495981966436cdfd4ac15bdcc173ccd2b0343736d73fdf7cc15e159c17fb8d956fe4f7f2d86bf9450260254e981c033f375764f81770e169ca3668bf957c77bba249a33ac84433ac903aad2e5b07366dfaad948bd2c3fd2ae6ee02a0cfb74f477c953a972bf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38ce6f0560e035ed5d2447b84adfefd81445a96adb97deac3e7c23c999b7b99f53522e477505eb8a6d7e3ab93c706c1a17e3162e72176aa6a26d07e3f778d541fd8ff708980538dc81f469219de8850e5cdc278ef96c17a1bb1d4ae834b7dadf535becd953f2e08de5df4c1f48ee00147;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb5428faac2c1db7b37d1e37786d72f5825709036fd9616172537d285e80d73f5385403d27768f82c545843ca7b12517119d03e4329fd270fb72f7116ae26ed81087839423a61eab53f73ee01025eefe90acaf7d5d3cdb5d3355d1ed1ba1f98df0e7e4a3d63d1711310720dc5cfa945df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12ae795013b9b326e31839d9fbb77985a281e217b851566be8930d33318d87432f62b72b18e057f4e4cc55603b9f316a8f97e00ef0dad9dde4943c3d71c7ac172f36507ca8f6fbfb97a231ec4374c39ad51fa6a7859b5b4d0d34cfd2ca63e29e2214684ac6ab60958fb7ac1c7f15f004f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf17b0556f4cacbcfdc8a855c9248c7bc4d78525f8791a037be66d8935e2a41a4435c8aacc0bc9c7154dc4ba105bedbebac3c5ca87ab2d938278607cb27e39b7fc249edaedece3107c1ad4a8cf4b974096b4654fdf2c57d48ac00ea739cd3d972335c3691b728194d0b23ad473e2169920;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca4110918f05f8e2e5774556294b7bdf5238ef7fb038a662a0092ce3bfd98b75bfec063163194d51d0f6417446f91484f64c587bb4175b4ba86a06399091c5e51a091b343e12aca3fdb0d3ae8fc8d237e1be934e36d8949a9a8dea1313673e7d566fb16361e9fe9f90c0ebd526d888255;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc790b5cc9687484504630393e643aa894b099e690174339f6dcf30c5e77d80f2b92b6b30c9a2b5b15b9aedca366edc7bc6824534e55bf0cbe32ad1a3adb8f9654b04261f6309dc8192f83df20fa25ce8b0c95a2700eac678a1cfce1748f0318dcdbee4dd71ea6a2073d8ad950a2640dc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49239415508b6d9b1e45815f4c3684f84668a2cc3e494af7245c94f7afed3444dfc492d3001464fe4ca47637b91df25ab5ad7068fb3c42e353847e5f220892ed00049d9dd259add558e35ebaa29c120b387900095b557c2abf7abe69e8ec189935dee273a7f4772b96d087ba9868b001d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c71c89f9d882e3c34108190a10e2e0ed79b130cfd73ff170a29340ffa9f9b62f6a1c6338724735a6dd8249239a855288afd8bc84e8d46ba582c9a03a2a8684589d24d2dbc354c8fe4be12158ef4a0ff8b568aa37389353f909bb2ea9be189734626008c5d26b75e6baf2a0cf5ae832c6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h597a21b3a2d57b4eb1851b2b5ad2ef438b07cff52f6cf8fe57890f59a3907767393092bfa59e817b7bf5912e53536f00c9fe6be0a2f7d6a897fe1c8e9e510084c691cc4363afc2f1e98789e2b389fe923949302614c17f59362f9392931d08d061676e2743899ea40e5f7a07c82e7086b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37ff25beec787fd21a56cd42592ee9e7a103582d3e0650ab531ce217cb05920d645d9559ea691a35666358af53ac84961b7045ed8a803476964e98d33a56dadf27a9313f7caedc4c6473846d068943ccc2470679df1ca3508176f79e59cf2db20b5837a267a5b73835b316585b31513bb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h82cca2654a5f97d206168057d865b2534864343ef4de293cf549d4eb6ec1e75b5841ee1c1034cd46812644eafb873a3baa7567ac045fca0c69fcb30adda974bdb3b56ff27c76a40f7ca0b026e41ceb6327bad3777e6f9732cebd396f7188070c132ec0d60b9016be7084c497c34a90fe7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h77bdf357159a8acf20c4e7edd8c1e2c4bf37f618bae3bec2cd768ffd7a49e476e164bab6e68fe5c9308aa549e87ca3cce57db4d68e5321690dfbbf9570b82ab40bc53e6e1dfcdfaa14fa39191a58bb4670a577f9bed48b1528549ccc2ceb6fc53d48781e287acd0ab0da6c1de5ac390f9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab0f5c52d9bdbcf775524553c8f69b95891f1926ffc5588ff7c856d1619a583f30bad18eaba569495542a6d51fa72ec1b01197d21c9eed87b8d666ef5d5d84d32b2ddbcc808153f1ec31de10d094e5c5201c66db2d549a001e85a1fe69de385e73ec38f2ae50fffc45db2b0e5681e2e95;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e1beb68aedfa3bac88273f59c62bd5668a1851dd7e6f3048081ae74925f386d870f187efcc9845941c0fc435d324a7f95c5b910ebb9477ddfebb70339914fa6cc66f7f2ea49651dbf27c8ce45ee4638b987bf0b661fa7f2f72d52306808203be1330478ea6bc4f915525a75ec62e5e13;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5c08c27973ee0e46bddf0a4ae7a6ce2ba9e218bc88d6766ab416092ad5beee9382b1871482f6be5cd45033f515772e6ae09be9d5069f166c80d865eb17fe99311ba026d9ce282c9acc48fd63efbc7773b98a1169ccee631f9c4b3d765c5d9bd339fa519011562ff021bf397a98aafa28;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa46b868dade0b721f7def84328887e4835228c7a738dd396a41fb3c9d289a5c0d860fcab962152f19e37540bfec102de810ad0e306812e42d6783113a2d6c89974b213b247855f6d2e2a9f4c82aa67c120c7976f91450b76a7239a8e1425c39030ee132c68f7d1c9e9ff6a1fbc776e0b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h834bc0ecf3a9389965b09bcb0390c0e9eb7000b6c761d0d6c4e4c86d35f9c5817f5b553a862eccbd1840bda63d9e1226c708ef306ac8280e7d74a34ea7cfe457e86f577f192e4e02fcbced5b564b5d426d2248eb9f727b6cf8aba319fac7502ae276ff582323907ae90c20e92a4894354;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd3a30d42804079345bb95a4fc88da7f298908378c56df7296657fd8108c13b150b35090e7b9b78caca9761f3044f01b2e63096c3e4f602b3b97d19a58ae48be30266655492383a1a799f5a44b9602cb7af3c2432bced2ebd8be20b9a28ef0c83a312953cdc6cffc9e6e8f00dc2bfa8699;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfb8026fe74f2e63b07cad5e787a0a166a46fb451c1890b843afdd9bde1fba415d99895dbb0e876162171e488f2731a11702157172c848b2c1c55ccfce4f91a301950d8a8a7e5f8a56bb30109d58bc4a09a1acc5438c4e3229be763140edf98eef835ee6407a33d0362951eb720a2f1d3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h67068468da45152da55356b76c1d49b4f8bd615052a5461ed4bb45c79b39f2a0c20cc431a5d1051b8f9e88aefdf963e06e6ea0df56235ced9f8af44d6c202cffc1e59c37b79d40397d4ecc61cdb7fd8bf1430b174e29fd037516f8255593346ece16341fe733691008369defc80613420;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfea0648bb4d0cfe5652a8ea79fe36b713e186ccf768c20748678ab150b5f48983e57336a94b5a77c17af244f31940efe8b20b1066b7be4bab768d0a32851ef207212c0a972ec084f4888370ecbc9b27332be034f8c098c3f22e5c436c0b0ed42d661e9de7ea01952eaa8007223b18c938;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4227836b5f1f855755f619322532db0ab55993a319e21552bff0e3fb85e1ad5085c0126126a1efec6591d8a1d0c8e5b381fca0b9ddc283bbe8829ee9ff56f8e8b5906cff4a9e5ee142fd83cbec4ae81df6ec0757cd5ff5f49f279345faa63b99e8c14f1d0277cd5f54fdf6ccfad26b60;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6834feffc196575ab4260f455c597c0d7eb5bfa5d1266b26e1ea50d1be2cba8f30cf266c6a2d57689734fa324d6739ea44c21ef7b7909591ad272d37f942157319fe5f023aab993fc5ba8cc6f86d9091171b883495cb769003150e9ab4f5bb4b42c952dbb12acfc86666b0394ea6f5e2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff7f12efcaabaf6854b11c16ab9cd4f855cd7468debb845296138dce529ca58abb708ec81aeee56b6c3518fcd67ad72ba2ce163517f72a49bdebf2d5322e59f929d6e015bad4b45ddd05645218af55f5b76fc45055a9a27bbd67b3210e91bcba7d98e3808649698768f096833c8c4f8c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha1bad271dc05ef1c4176c635afa947d8d8c15d075f5d10a22eda3c254a900112b4ab301e24466c9a51d32d0eaeab332ba5f8422bbe208f0afb95f82388a82319fff3ecd7b3eea7e26c603b2794d91e9b4e14e8107539ea221299f531116a15af1a0fd561cddc00e799b2a7413e6e2d574;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9fe2365bdc3b1e8727ec18a758b37bd44bb8c75031c10faf91cb99b30f00b100602009c86522f5fe7646dc7822342dc822527872d77b9f3b01b5ccd5e8f2fb86604c5f3a0de36d906afad0d982e45a3c13badfe1805a8c970700f57bc79f30444313663e7f331d2c8e4f56b56492b4e22;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8a22ca29e4990a853ddfc65e9ccbc05d97a687fc1d034497093dc12aa30837bf5b9905aa2b34f0a0fbc71373a7d5abb5742682b18dc5a70a2e9e3bca344e675d5d98ea1b255003b09261b52f4331cfa00d8ad89bdb8d77787b972e8e7539a947f60b3b2aa92162ef9c0c615dbf953864;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7954be770c06d4a596c996fea3606212e350e73c447791a18aacfc786fb2a4ce72cc67263dcc7bbd4f767ebb62f05fd7c53a7c6446edc9c382f86cf06a9b99db8611e255bb4389ef01c19a66eddd88174932a75ac5bcdc5a81b1af1b3535a0eabdc38af36b11bf15f01c9f727baa057e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c09d3576d72a24e93d313c8d035127198429c8689f59c0ffae2f4e5de4358de458bf78b97ada049f48adfceacbfd1e687fe4d1d1a6ad3f75ca0fdd175b3493a534efd78add3f2b997bd3eafbb4d333933bde12171613859566842c67528e3ed396dc7eaace045189cffdc8428bb609ca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6b839da97bf3cbe169eae87180565878fc7c3ee319a8d6ec7227e29022f5990f9b51ae8fb84a4f57d1fb0e671ee9f190a32700962aae9a98e0dd8270c56f598fe0a2824efd37412a9112b88684b2e98b7d8398450b6342df62dbf88dce027d1ea34e38137f20a4ead099ee082c38607b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h515b18299184b6f43ac68f07a1bd19b15e6e1fed6632f73bd99f334794940bc87239aebd13400d5ff0988b0e6374aeb863887dca3739fcaa9c855f48ab33bb9079ed0fee1e8048f11beca638d6ea7cd8f778f7cfed11f83bb79ca4c7a86bc1b9abdbc64a84c56a5b7a2899709bf511e45;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he21daa23d8897aa92b1031e1a01e9031cd56e466e64fd8c780ebdc151f5cefe1897368127e4e7ad5eb5e83745d49c69c284923c892c97d77448b4ce94d94e1cc326922e894e508fc065ad930adbd901dc36c59753f0247a061d458036eb667988a4e4a17ce4c1c92980de764b337b9580;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8033dce3d79f5c1dbd7789f1cce55b2239df6189dcea7023ad2a3a6de42b8409d5a7fadbdc5e6df20ce4d53300697fa619aa8234855cabea51200aed64817ebd96055d95713f3e97c32379b3317e7eb4a1e9809a44b5aa8030facb7ca107e82a27e35be2a7caed03efff90195377b5f70;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3bdcc67e560d7703c18a912663a3457ad0d4d4b868a213746c8cf4e18b6011071a02c382aa8e45f49962def81c0d932412af7e072b460095c19dc891964f792e3df8fa314d3188f5cd2e7d3812b304b6ce084ea1d33a0224833a6482acfc77c162eab9d422a63237396dbce0da0d9d6f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc603cf36cab06eb9c245534e103e09d580d2212829b3decc37e95f378624e287affede7c23318dcdd1b917ab82863eef1bedc0b6836bb5c93a3f79bbf9468080cd4de35469cd0c16b6e601484e3810f8d64a7b7c322cd37a5fa454d37977d69d9306b6b7992461b53a99222607f4bb9ad;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h430e416e2782143f030452aa03c098219b6ee08471d726467b4f6b1ecd4d1c9a190eb95c47158bca05d110ed54ff92e5e7073fd117d294e16026292c97fc2edf848427852c1baab584d26c8ec12c02ff8750c2341c123806ca8f1de8f60a8290d70b08804d8d7445095cb648bcc615fe3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68fad5f91f935eaf3de35620f10777478b9ca3d507285f8ab0c8f8e8721da371b985dce4aebd2d297730d09a8f08f56fc5b1b8ebe0b782a698c1247cbe5160b9b56d53a2e577989b73b1182473bb19d8361b37b522c7ccc8ca115df1ec636e77844b4eef496afafbaf2d520a95f654eaa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h551422dc84b0b843070b9e72a0863f44942f642fa5c6bdb1a74283fe7205877f43757488f62b95e32b735cf2d085123283394b8872aa29185c957967a05fcb219d8b8bbdac1487462871b77e0764d6029b932f0f721ba62f8f3c3d25a65684b9ddf6044841d4bbeb8c479737854c8b189;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc196863d952f20af77651ba692325876ac73adf095dad6566e695ecfe17f0e99d3a8c5ce1a7b31dc251705355eb7e79ccbb65915b86fdf2f24ac561d300573548df40e5097de81b9fcdd8527025e172fbbb23a17f0997f9b6f564e2456f02c6eaa8b2026689354c827a5f16409970de4f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49fb3b928da26bba34c7f0286f947ed6c997522e0e5071a9720f4a06554e13894947943b28c745ef8f54a44df4bb2a0fa8155c505bafa0a9d170e0a3f6c4cdfbecee661ecbbd14ab9383b8daddc70aef564f79e8c6670d219259998744d5b2617258e9377325ee8548280a050eab91f34;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4113400c6bd3dca18a202ae159f219e772b34b8e16018543c37d89dcd053083abbea51f0d80364b7c128182332fab330c54e089c607cee2a4c72e74086c9bf33a1ac9f6a349861705ece8836cb06e110c3cc2f5a5381c47bd9ecfc43bf60e5715c9eab8c64bb3a417bf22b438530ffde6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a2811ad3440006345e48b6d9b9123bf5c34b7e74dd25bf2a112d68bae3d196be82af50e7d01d1fb70a9b0b4192cce29f1fac9d71406db87478e8091d523d2a99198652abacdcccc4d1e6ddce527f5e1b2479262fad7e58b5bce369a6e66f8cde78e5ac1ba6a4991e9ec33467d8375e78;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8957e2aa937da60db654dfccbe0555e06472ad7f85b1e1f1c00cfb9215f8ac41817ef179aec1d2e0b6d752c48157c35697b90ae96e33ab6fe49350ea1daf35a3c30354895883f2b6a66cb639c9a36bf73fc8b864ac68a32dd0e1247594b5086e2522b9c22435d0a3452f84f6f61e786e8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2d6b401d152310adc4bfa1b8f90e83b31eeb141e91263e00c660eae30c8de406e34bd8c96cfbd935db04c969e858aa81fe8412d9cc64f943550e77e3be9a8dd2b994cf6997247031fc8db65b87d09cb172f304182d5a8db8b45698c86fe60d4b03ba0f22603ef266c3b87789ee2205a2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28a96d3b22f5ccb5444394519a645d4af9532aea51fe3702f4c53cee836787dc7c9a9040ba7d9c34a2455c3627cc7f3b2e817bdba34e9d7cbb5576e810ae7062fc37d3654d12698609e107c727f16a5cef60f32da5f4c757e25c43bff95a1d9ca6600ca800331519a10404887997fb227;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb34fc6fb64424ab6408beffa3247a7b68f5fce0261d8b951651fe5e2d6a9330558b09f0afa9d8203bf6665f554ba4e5f4597531d226a1d6e950859a37b6a3b54c5740ef3d223ed07296f66d21b468918dc424147fe1660890d27431fb3bafb587b74977f28ce5d389fe75fbda16905435;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc7bc4db45c0943ba5b794cfedcd85de260f0a016926353fc40919042f3e5d5888617b6b2ee8abfdd50211797160c6e7b5fcb9606a1fa471370246596c4355c45348213a7cc88daf6b563a27aa589fb35167c236edacab162540f5d114628900c451cc37d6687720e3aa9d4c529a7837c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9be984ea3c635c3504a8dc218859a510ca6846ef8cb9ffe23b6caedb1ef7d7aeb5762a2aad0c97ea9241c20e9eb5136dc4a3cfdfb13f8d5ec5028cb6b853071476a80cec60c77b44b7ce39866bf98179d129e717d1148d213b18c07246f6a1e1e214bc92e5f618c376fb5972fc339ca1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hacdec5d233c53104ab25e40b59edab85c26e2be30e71435d3b99db1b65ebb3fd9bdc0f8c0e8d6428031efaa40b72583dbc7b8d01c76e0a659ffa48c0640101f8e1f9aa0fc43510a68054164509320a69431779c88d1fe1dbdce57405a253da10b2629906c2617899c9c0ec706c5922034;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce4c5819574c29a8fdfcacb6387e4c7e8c630e051e13569f2edabe7ad7f1b0e3f6d07f3c03dd7e0ddff13d2cf5c2930d3f577d42b9b94d500f4c2df40948110d15e59b1669e32e0c921b6e4527ed36ec7eabf84db1fd607fd25a8855e3b77748a39106ee430ddbac7f7a2618df5c9c6d9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45f4cab1854d741142f118851672090b0e3d55fabeca1d4d236d6036cb705244cbf0e0d3c1ddd713ce5c134027168453b4312997083ca7cc0712360cbbd8ed574f3eb92faf7a17988f024c1205e09d70489e3353d28bca9f8474ec247df6472b73cf2d8ceb25ebc46a89ee82b93e7482a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7db23b77a089580445c96f14d5c5de815c592632726e1c84f068c4e83202f661be0e65de468263c3941347ba420a96d6b1351137f3fdf18a1df84eaaa7a47ab88054bbf0525e97391d6a3c0cbb857b1892c7c9ccd29cd3aa43cb6f55c75231980180ac9e716ac13963c33a2854b81e5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1c8e94b1f4e294273846458ec9043fed0cf7357c52bce7e7c31a3b9e6ae2f6462006257679e014bd0290a742c8412e3592bd6d1ffc699c88b5d0d243961521bdf080073ed7345d2f68aadd97f0c5d28c580203306a11e92d63e1be603da4ce7bd42bd49c4c19ba808225391856a3c9f7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca9203dff3a43655f7d5d3b7b420fb6bfc24ece32414694efc11afecb93eca8c8e46937460b78f35a8ef843474788edfdf05099b6ee570a46f20646cebd1569d3d7c5aab4ed374b59ea513732590705745659acd51563fd4e8820701f1f73b9ee901269dd93ae06fa3bb6f7cdde23624;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a9aa5d08b2176f07cc110b57d3de6b2bc876e22794893e03e3d817ef9893c7fcae7635352618901969b220bc074d96edd446cd0a10fb7372762e43fbcec3edbbb4bf2c764bf151ec722c60ee01d2877eb1bea1e8503ba9988666ab15a762bacf514f322504dbb4a513a07f2297dc2b19;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd39759788e729f9f9878a837d94fcaa8d1632e5576b4d16446b88df1b733afddb43b09b6853157f2053cca7c72407751f9f5886e3748c38275c62c75c6d2619e1251835e7c4e8c98a916bff0b674e6cc5561391be84e0e1050ec2899f9e9aea7e81815ed9554b36e458cb7e6eba9ed6d8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf26a2ac8b42034cec39a4670ff33409449ef2084ef4696275c4dd883435bd9a8bb1b6a5e6f4c99c58babbb0c44d5e8c75c1f94e19c79f2898506a36d27fbe45a8492f4b5c49cffc586cc7cb2a134c8004828c1f1bf9903a901d4a200a3a7446bc65a4435d6601449dbc8f3e2b558cabc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71edc21f6d4a1e7feb18940a50ed4784c11869a16c827575c180504dec3476fbbdf65dcd4d60ef6024853c72c1731a421120764490003ec4d7f9da44583a08ea60fc850e56d332b53e63f05d88a115a5ae58e8a6c417dc0e24444bad93dc345d1528beecc97087899b7ab7942f7933737;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfea1396b3e21ed7b15cdacfdafc4a14bede291ccac08e91a06aca0595f6b01c2ddc3029fea42d469d10a51e92ec4f828b6ae78130f7d452708c5cc036f1955568ab671683a811bb6568a5ff620ecf6473178837dd8fb5879616dc8c58c01cfaf3036482bc23b3a8bc6fa43dc9ad607acf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h804767636a98781b45da922e6af8049c980e6cb09b3e14ef539fb2fcaf747ea86ce48e15f5f825d0ce2c38d946743e5f2d3b73fb51dd58aca6addf47c22f12d07f424ad73a36c094cc4a450be915152efecd95aefc151848c69a89230532d3835692643aec6edaedb94dcb2b6d9bad33b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f03d2e1e0fb01589eade1757b8609f0d13ca2edc05b0232fc35af832b18e0b495429568ba160cb2d4b783f67d33142e2062704109946aad4dbe285014daea331cf5630b3dbc1057b18c43e68712220e6af6e5dc7ae67ef06668f7a619a83c1cd83f87fcee94aa9a0cc38ec4056d28aa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2284e2ccd29065cfa4b3a372e688f7e16aa830958c2e5cb1bef16d6533360cc2b8c32006c41f67208f390a79aa72fcd204b42a669dde08a3b7f7acd091e79a4764b889b9231bbee46237511db1ca075a04f42a93a612a422ecf17a78fc2e6c18ce445eb573b7869c3f077e90ecee45223;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha16c947ad6b64813ade9b8c767ab4d3d5777f206225faf2a1f7f6282f555adeaa27605a2dc44d702c038d0e4b31dcce6369a7c6438b992ea5be4f41cdfe2a2cc3e9ed541eb0525c3046e833d328b28e28b4b1dc39b49db0a362b7b2116e299c798cebf7af2312309fa8b42a41505c59d0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce98da0b679be17dcdfbc25e88a0c98f4a8a2913a6ee15b6fdc92d097154442050bb31a2e53e544a9399f24a4411bc9b800025b83a4f230465be10381595d7cb54e0e8ac82bffecd7b376c9daa743e732f70ab4fed89040908ee7a65e3932487e0d3ad88cb45adcf4f18a8730d496368;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9132f722ae592264766531926ec951e25d73e36fa25038475a70ac48fc1b1b474956cb03ea948e56b0fae21e4e4acaddcbcece5adb9f6275f9ab204a3362bd08703ba2c8498c0171b6c0cbc236bc4ae7a29c87b891ef34c88148f4ae36dd2d6b8d42605a156bc14eae7ef21184d49be6a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf6cc2a36b885d3412256903dcd0981618c5291f7ff2d47fe285797b6dfc46ce34a81b6a74d21cc79bc8aa1a5d67c37260b5b4265a4f1a0ece26324d88d3bb7a35c32adfae4fb60bbb5a251197585d864889b4e4cceb69da09e295b92b415814a836c91a5a67781985f14a2e00cd1815a2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43efe8b2bb20510a197e4a710050db31926a878c724212f0e967f9067196554a86ba8e927c54a1cda5e1b15fc4849722e2ff227438252dcb5017de867c9573bb10bb35986a88066eef42de0a024b4eb5d059fe939a41d087e934336dbdedc3f6d551f5bed35e5eff20b0b7165c3476952;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd5fd079b7c0e3dd4e4e818f32927774ffe18bd3de3d8c86439858a909cf0b99750b0c11649c71dc2c71091947920b89e98daaba0b030e4d2bb75fdf70f9229ae8bcaee4730d25f2ca50712ba93bf3204e2ac4eef920f88ce6efc9b361f488aaf0c5ffe133e5996f28989b4ef1b44cc7f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h148ed842ebf3ab78ad3b473080148ff7ade91269159ca388573885d6fc43773d61f191233ee48c1efa26cd0ae4569bd3f4d3c9a7155949d9a9583393a88aad4c76370b42a20fcd97e627b39a00a4cb86da9a6dc105192b5e07c120000ad43c32aa3898608d5e681b94475fe9f7d623d0c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4632ee3ccc71fee4af4172253996a646bfb2654955bbc67634f9f77411adf77263425ce0062a588c687dbb33737b8ce9d188515fb21a12162fe6ad5291c4c6e682a836592003c8b53e8a2c4fbcb73adf3e50bf7de39d810280ec81523c935b3fc009319f33b27f3e45d2a4970bd4ee41;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44ac098464df65fdfe9e33bdc46f00af5a8ced4eeb3fd7f1dc7b54a4dc2588550e4493228f43d1f57bfbb164d2031ddcd63fa30ff9212fac030e4de3df6eb4eb65a2b61c79fae102046ca8793d41ae816293204d1dad5f71bca38b055d096d369f2010a31bae037aea961f5e9dc8f2d6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5888f95191427640f8008452dbfc5681cfe73834f944b1fcea7cdb80c79855ad3846b3ccf503982ac6b30364238a6248ec04daf3f356078f8f75a8e50d760d3e3b6c413e651b995738a64783b465bf2cf53074cf24b5cbe7d376b2646e300b13b4710a0f5e10cb5836075b730c87f50f6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d69bf36d5d3f17ca6999d491322891df8514d30061aeecaa42f5b91c7200b509836d5a176078a2d4ff3db1422ad4dc8891ceb8617dfed829743ec29eda9a3548b40e6e34834529d0fd951e05a3022473572df327df512838a784a820d3152602703574b84c0db1ae32bcc0ae2eeb993a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9bf68e829d9efd4135af75798ab9370ea05f9ba88d0cb0b02e7df1e30206dd208e7f802f5ced16576ec7d4951c6b7bcae6131098e45c24204f36c6542ccc7af8eac79ae0875c29f650002dde52f9ff5073caf3d00b9d9a086053439943caaddb0628eaf53d3319f8e3e59c15d43ca81a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a5e88e731a07440801fec1509c5b1a9bcd2410d9f62237db19cf0858fb3305b465cac1cb3c404e0fa6ba8d34cb05f483c3ea6d8c69c2453e9a31eb386b2189ff3e4df537235ca4d30fe35b209434a5e334760452f02aab4f772d2a9231055ec07bf9e5de88e6a911fe219e17fbfaf040;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h966f06929c7799f3f5a14992b57f8817ced152a3f57a65cee8638907fc77f17b212cd4e06f1e10c926d9a0abab82523030f153efd1fefe7ab84ffd7564c94c09c5943411da17d26a270883f745ce2546c528aac04f50f4b1e7421e6073325e0c8e91731fa4397f77f746a4c7d3cca1575;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h536b08eadaaab54761809f0f54b66dc9e088146f9e9095e4e154c8e6ba82e3089f7756372573b338ceac42d270334f28270a032373206ac8007ab8fc23f896b0435cdac326812641058775e1c904deac80b4aa0054064ac3c172814129fcbbc6ea14908777bf82af5b7dd1649f294400b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h60da0100b8db41d6264799d8ec81fb8f5eef6619b35f456ef19baae452b25c0e916cf43073aef3d09fd29ff45e8b5be9276235abcc118ac2bd002af0f9b63a75f62e26bf7ea42669fbff4b79491d085d8dacc770fa4b0f976f7892c7968973dfa0edcfed3fb7abbb92160dcc2ddc861c8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1da945b712af4afce26a031e2d734af340474ba5a0cc938f839d9fe727f1380b0c150b0b9ab5377dc679035950a7a6d5017c312576e0121ae3f308d30702db465f3fc0376dd76923ce4b6e9b7d5fc74593695eeed456417f46a4d72c304cd104be471717f170b775d5a3be6367f4d5fc1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7499a4a1dc8871ecc30ccc3a27461ac4e7b621102bafa5b40c19e361f408160687ba11ec3d49aa15fc5a7b17a6d441a1dbc29df9d0a3f582790e0a8aad20b7dab4a44c49d243d76cd65c8002b1ae880851707decba4c240a2700881133c635d86b581786753cff2544bbea4f54c558c52;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38ea74feffe010f96fcb74395cd81f06304686c705b06047ea2e7f805af390e6afb4e98951f7bccf3f7b4d84b34ac6960dfd44e85b76124024df87a5eb7506d99c16c766d0174f6615711727b8f2fbd1304c2d030577319fffbb65df752b45204c91214d9345b0b61293f814a3ce65cf0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc79b30163256536544602e64377bfc785977df3a2cced4e97a16a2bb31f21728e9eb41b257e0e4d47817dc2304ed36a5ff915088f3731abd50f63dce30b80a64a201769dbbad22e8917b5cb1ec7b7cb9535586ee5825385039a7aba48d77628c2c60cd34a9c2b1e87dc56eff3c909b228;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b49841a07e295d3368cb385f6ffdb1b9fa6f021df4f93bd4c93ac4af2b7421cb74e06f3920033419b9610c1606ca81d493d912737773b05c4338655c1ebed38671b8d6df25ae0d7c35a9b677465e7c6c8e20caa7dec7ff184cbc7f2c7fb1d3036f061831ab554a84c81193f784ba6c6d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7433d76611d4b1c6f57468671a05ae1f813df3fe4b47c7dd7fa5390e9da0038794e4a176937d6acd960dca887e49d0b845bc7820df196afe7c4ac650e687c12304e5b9d460dfee32ca41d1cd4d53a3860732363dc31c8815d77e460077bddeffd3e5a058746eec5f3791d41ef600f3b3b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe03d15eb54b13242257617cd41788fc3e10380758af2a1eb180d86e85b764e3f84b8af44570df68dc9ebad185aa97e6babcffe6fdbdbc5014fb8cb2b66145caf521220a8c9868622de2e842624314c947bf43fccad32c2a7ec7ce0f901ec8265439521f23ba4913443a7060d7ac7304;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he83e59de49ce7f7e7397aa28ca3dd7b5e03086ae82988937c69db59b05e7d225712823615546e609c926ef77a8ed8d90cf6bb7641a11ea62d3de9e04b61e009b233edf4123811173c811abdb560575a057ec7d13beb6fc7958147e1a1f9bfa9b349465085235a782a5514f68c8473f743;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb71f02e474e9c310d9af9b2641015655e94f8b5262a7ec5aa6ddcd094aeca9525a753bebca86969c3e86acc3caa0911c28b0b3f5a22007d28c316bfebb0e18bc3331f4be5d3becfa1e2137181de63375678aa77ab012ad645dc7a890a7762494cfd0ab10e7a913e7f687474961555939;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed143b6b47c63799c42d4dfae09575071e7455563a09d17b7c9541679f754ae8be2c01dd87217c40bc50f69f4c8e0ef562debeef5026b2fabae9197fc5ef641915d0f2f8fc30e98b5c167a8238b7acd3984abaf21bcf4185db8a47c2910bf45831149f4b237d71179b19af9c63255f3a0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b82ee2c0cac0025fff885f97182117e54827a9cb10ab954f29c54539c0ba47e232d732f50893302d1be153bdf1e900df86a78d58ade6182c7e31069a8d5ef51b2daf291f96417ba42baf5ffb17d27ffc4f9e67a0533eb4f1dfc402ed7605e843f803539a261df0a82de2f50132ac91bf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab48886fa1b00cf4a34b3e3588c08686720a1921fe235456557ca90cbe6fee13188b33ccb1500db5480db301b32e98ced20b3796e58fa17e9e1ee09d13552b3668819358e9aaafeb45f334b75b7c204fd82ae7910168b607c2d1054f5cf99b0c0db2e7fdd33a9fd7db621c0b772e5be3c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9499993c663044da1d2340da2dfe27b9962eaa2ecde698a71449ef047199e1cb4425d3d3340f342954fa4bd299e914a89954f2b27de620d9152506692ace06b2cfae637af99f99961b41ed6459a9288b815ad14fc3c24d1de8f671cd90416b3507571d6e54ec27230768dbb70e7025c68;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b238ae37c69b4511db51ecdc365ca3b8269c8c08569d5b17a31069f8bbe42030e9e2c07410ed1396a13d08030d7f7a5cd2732442a6a30cca976b71ef43b42b4fe86e0f9128ea6f82cab2d60725273245baf07a3580f5dc6c0b3fb1819e4b127b5ddff59289204465e8a8d428535cd2f2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75fb3cb4b643051ca6322850fff281a7166adb66714e613cc2ba2991c9283f5408da9a9726be16dd6c7fae2bfe399e72b8b18d7e2e5fd13d4843fd4663b795935dd5a1e8c64e1465a35efa18b474def0dd493b05d4ab9e34099def002f4e0ab3fb0bb9b83b39dfc34597e0a912bc087de;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hecdb2e9767f922a1f74665c2f84d073412bfbec63f992440c0d39e5402aa55c347b7fe359d338cb5e3e5cfde3749c13969eadd5d9bdbe6f4e89dfbc17f2a0e6fe844c4e8d82bcf7aeb91a85d73674d0b3863204941a0f880a84b7c6e448ca79682c0990cc7cd130d5689a0e19060c61f2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca1a935d4dda3f7b2e7bbce4a359b69d3ad50085e3a729131c147518be5c89544707df9d8c45a1527432b0c069bebab0c6a814294a157ee07c54a7d2a6dcc79b405a41cb5554ef64df0cd69ec47804e7f8e3499204fefc12dcb90c461cfeaf8a9e24b4800eca2ac896002aa72e0ec0732;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc01670bc2da2fdf5f3d826748e9fb48d7e42aacc30c416a6b10a81bad877b1c835eccb45b88bb711d91b3b0b6cb898bfbba62e6ba913b47c7897c880a669118eb445443cb4bf2e75ac12f76dc77de13e19efe42672fc2c3c18eafad0527fd2c57b950c6af7ab647c63fa4d67893177c4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcba06d36b8a475212495254cd4841b48e9ddcf65b7487180c91b9ed34f3374fa2a3c0c269ac97bb942c990ba29174a5dc4a33f53cfc78288532dd4cb4f6555247c9da7ee29c40161e70d2f1685ec56f8401aa23ac7b671464a3538319dce418667afae96dc38a1033e9db57b668495e22;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5be78c4dfa4bfa66703d71ea205c4c0ebf76ad043030e3e944cec8c9f31bec282117df7c968475bebc4f41d026979a0c0cf144ab61bc8ce497c0145bdbbad92ee381d6dde156962e2ba76b44ed9dc5025521e0d2296f6678584d696c4e35528bcfb666c7e076a43f3ebfadaf2975bdfed;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98973aef5c10e878c6d467c8cf327dc580119b89beafbb44880f1aded4571136e80fe30a56afc0c4ea4a89386cccd2a8de2963a0411c8eeb3f8803189df41541a3a0e50fd5852a136b05a86f31bde388eaa55cec7ba4997dcbbb9c7503ff6c78eee2c4520d5d733d15341a0c735dbd8e2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38442c436ff1ceb6b0bf5346cb7e7e839eb517183c305a3ce7c6cc36195cc1690326dba706918c8584d2f0f2b126b75e21aa2ee34237d1752ddff65ae2ab0fd1ca37d86fa0d0cece62d024a1f5b87125ff621d51a5e9324440c82a326ce10e5678f160a633cca6a46aea39bee1f7d538e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4976a452a6305e51bf05f6d40897beab715968a863f4aee8852b22f34b3ec3f58b340c08cff44a59d23656782b8969b51d3c78b94d8c7e730ce8fbd0cf361d58cc02925457023c2cae482faf92d756199e6594c5ef81b762dd6080adaaca99c54567f46b1a3516e8e8cda5737cd7aa37a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95b586d3826c02e3ff94cd42c49b7dfb6d100cd1adb8206c5349c2d09b0bdb6a806fc328ec791cc0bea14112de0aa419506041246484e6ba0475795962571352ac6201c6417e9ed1e3ef34c5d5b84ab926cf0845c6e58a3c5fa5ec348afc4647e611150b4da1e44c0a5a13a7b8e41a21d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2061bc27f57b699760715064bfddaf94316e621610b38df32d0f4fd22a85c0885f7d09add7aa6bd8c01ba4de8cbbc39c8315f5f536ecab6a36e71b2fb219dcb2a2fa7a680232819d62bd79a7bdbb0ae67f6bda9cfdfa92200c9686ef34c4230eafaa2c0e39e387bdf09acf0903ce1c882;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he63b925490ff38ef99d9bd1d93bd950a77239609bc047a20146367c8c4127b94b120b1e9ab82c119c299f1ee7508f26efb7379a214a94fa6deda850da7b201c3d152a4ae9e3b25a597390816f47ba442e718c079cf58b62a5c4390cb10b701497f0bc646edcbed2a44f1f23c38dfbce3b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha32cd3499e2117858c5b585133c80f67967970561ae301fdb65ef4b72caa2769bcd45aa849a2de360f54d4ea5901b33d9c226db4dddd80875b0f41cbda895d12423c833a0e1af440e38e873c4c07486d226291f1738d2d0437c325c97cd00ecea934345dead425aa66e2c8e5e2f92b642;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h18bc749b3b88fc4aadca267bb94bdfeb79076dc6b1cd107e8400463f798b6cd350fff7d304e1b20e3b112c23ef2c93aba32328a49362643d2f68c919f43397734d92c4690d4a8d2a458495d822f433d170a54f40ba4bc45da57af4e64e1ae2b7044b13570fecd4f392e4a492a6f5ec764;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d470ea33fc0b866d3410e352f8c63acaf8a347fa5d01a3d51440dc2e35c3916f13f3bd5111eae6bdcdd95c8532ca929a2cf23a47ad770ed29505e0bd668ca612a859f4e8da37a567fb3263dca78aadfbc5f9fce7c946d849481f14a0738846c9efb4e8510b3351eeb6290fcb3729444;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h782c58c72021cb56f0ee7afc023cbe35f3467131e5ba95c77bd8a083126c8a847000eac6841f5a277628a57d2bbfbadb782e4f58776b041103bdcb9d7137aafd5a4f6ad79a1407ebcb37c63356745dcdca8994f42346fb2d2ec2588f9c28862a4a3b67ffefe0cff1bb835f8fa47402889;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf50b38af868fa9f4932e3a61edffdaa61366d8908c7d9848868bd5921b42ba4d16d84de585248a791d852261c963c65268c4e23b29deecaf9dd4f64cdc627426b6870502d0e43728a7a7d5a4617b2d511e8c13e144f64fc8c687edc3d98837507f28029932735d07924dcf967e0bcfab;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he202f190a40c364ad1f03031081e3d56e4b9d4758581aae24f5f99d8b642704c73aaf3569fa4b8aa6531a97fa51df305a10b1c60e3ae93631d55e2b4f8fa754c02e59b2b6166c6401032efa10eea946606875f141c4b8be2331fadbaee74551ecd796f9252cad2384519fd646c1f52326;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa0d635afdb9686afc488382d657d3301a8b15eca9839f164bb01fe89523fca8c4cc90b66b74cdd73d114c6c1e66007a499ae14ebbed4c22463341c6ef66a35e9fef6271d99f2dc1457703acbda2edb0dd9588650322787ccf4b00c1b4a4c90a9c202f50c56be9a75907bb2205bb27d5c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h13ab51b7a3ac8bab8c34732d8a6849e3e00c2b523f08c60213eeca10193917e3af14ae7e5004999435f38e0b445ddf6839403e5821d377d17c36457c78325d08a74de36ed7fcf448346917b8921f7b82637127558a07da5a83654f2f47f55e190c6e519adc1dce9b37542a9490e5a23d4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb681e16dddd12ed8e0e9b41b2c5b047d86b7e63f0cc7bc4d59c9a25262503a0cc8ce06e73b563c55f12480fc154a8aba132a652e6c3ceb383977fd2ddd53622e4d16d50517406189c14873546b4269c53e675b416dc2e076f596eac51cd8b5013cbe7f506e7be16c833585df4f46aee28;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h468768df24d47e8702b1defc4896ab17e04b46f26879f66b443fc8d4e8adcad37a2261675ce265a27bc7031ab340752461b2fec23cecab7e23a3fffeb733d9fa1c9b88185438fe6c4fbf040805f8f43aca964ee37a8483e1511d6b5bddcc57429a3b00146c0c9265a86c180040bee18e1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd41dc51b495de8ad0745293892f90482b7aa8900089404d152e07b8ff330fde7e3ab388074b947f4be7e5b212a86a1ee87cbc788510b91b65ac4aac71507d2db31d5a4f5b4cf5a4dd7970d7cfa97e4c960df07d5c8bc3b0fc51104271296e9c34c7e3fc49330b6f2d13eab431b968b9cd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3be9e1894d19e522f7841a3e426718f55ffc0caca6ff7ebe6949cef191cf59e03269fc955b1e833de6616c90be933b92afa21202f2fe70f9922ac260c22e18482223b5bc93a3516600c2e851bcdae7d3060071aa1a5936137b479550035f3b217dfdf311f3dfb2a92413980647180d56;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed5fa8d0a3669e0743bdd2d4d42ca419b66c21701a11244ec0f49e252d7d1e2cd8c4493cd4a3c309d975518efd5a6919c1746cbda701c37e61c0eff74fd58e740fd86979b737dc90227bc31290c4889fce049ce3b4d3e1284c8711cc8be0d3f0adf826f639d284dd5ca0d97600c4e408d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c7c35c198fdf7d7b21b43565642ddc625da5d24bdda247a30a3abc2d7022ab6a7769fe10a45d500a85d0abd3042fd4ccf1ad37ad88e93028150b58d6832da1a815712874de5b5484efde59c126a5e090d4585d6f2f995c9240eab1d288e29e74b5736db55aabf3021423fa50ede6ca1f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h339260643efccb171911c204d8229d4075d164ee292268bbe78337f28ca7da5c76c50ea2f6b178ca05b0dace4d9c8e49fb49ee9c8883bcb0ab2296f6b4c5ca73eccd8a40b76d212c901e5d02385da14cbf87a59a89fff77868942d40b0e7518918ebc8f87976c67ef3dd1faf4d82d41b5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he907dc6bf5ea07c252d4af5929dc90fc803c9cc8426978c789b9d7968ce9dcd45161837fcb4b4280b3db8397a8d1485a721322044df20f8d5e78bb5d261815725da8f223600433e64096593e656825b541aa7b9dc971d775a323e2ce898125f28ed6b493353b834e6098bf3fd39041037;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6d48b8d776a84882d8ba7dad5f789b367f96fa0da68f6f1c067c9163e1d814cdf2d7b261fa984bef5fd4cba8260da87fb5dcb95c3bf71103262824e43e6a42bd6191aa4ea7318b84388ea9c9f4fa644b380abe99588c8399710c5648da4f1a854bd0e7dc10777910834295b14a09bd09;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h63f873eb2b6fb978b645432f7490d6a751320d4dbc1b6ce0a642ea499fdc32635463b3610d7501e84004905bd8047a9023cd70581ac3601743395d3ebeb19a872b430855f1034d069c4a1d1644d62041555fa782786813234ce88d3732b5486df46c786087587efae7438576d6a8f5435;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50bc26bc2106d90b135352eb96b5d88dc36132773df01b3f17623c608d61ba07e0fab229430bc1f31c8c9aa87fc339b148d76ae90f13b44c4c532d3ededab5e08a8bc76374fca6c02be55a1eeaeef597730884c5e3988fa94e3f2ae6d846c41847055b1a3b95fdcc83f2a35194dfbc928;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2467ab22af533bc2c79f1e87d72e8833a624f872fb513f04e86c0340daaf0b00d65ea30ef6932c3b7ff937c2bf660b39005170c474d633b529fbfce5927fdb6311bd7010ab957d1d6319b3651f08822e228c826887d1df1eceed62d44a3e3d352000ccb325b2ac4b4845fc61b2fd54cbd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb85e82a761178173e25c1f62a73915874ad5a81b50f1d89c6872c730ced3806b0448d5beb0079214e9c6b66e0a98fa048b68bf6b7d013faa9158ff0d40c2d010d2f5761986029f68d6bc7b4fcf4d1592d80827d143d5ad786cee85a969f895b3c066998b6e40d5d379242fc20ceb53e57;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd69ddf1accfeb9f77c87ff3373075e076ab3701a3a27cea98e605d35f958703191367d78d0b0df271dcf6edb217ff104b3187909bfc9496e78144e415b60d7f2d3b7c143392f86829dbe041897bd7aff68a57cd1896dcbc605c68b20e7f11b9ceef702780b3d835dc2c115aa7b1bb6da8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd7515fa73a8c13b724308b7ed5589871811e5fdca163bad601923f40f16dbfdcfbd1231228940efa5729c66608619ad0dd4dc3cabed18fa63195e7310bada145c50413fc003c54928fd2d1eb4939b861d8a778c48e91809ff6550c8d7f2eacc5fea903ef0307b771e251705a4c798de;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a0573e49b9961addc9e4314e87f08d021a1a0f42aec41ade16101160ccf52712e608f4ce34f985e135af28876a5415806aa9b3414bd64d35bb45d42797553f3943d005402216fbc988b2a2df57fd20e55f9a899ee5d457e054aa8a370579ddbf3637135f0e9bb608de5c56b19795a86f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h177fceaa2e3686447549d2b7ddee8657bd80f5e87380a670e4d3be1988b0477957130bfca9f0ec02b52975dff143116817167a0e1ad8bfb20ca1e165dafe9f3773d42ed035e576b96d93bb7a10e9dcd1ed76286736a27fa1a90b8a7eb83dc08d13249d30b669302d245e4823f4abdbfcf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd742147d9078e7826908b3d3b64cd880ec832ccefdf0bec35ef04cf890faaf12fb09a954485f0c71f3f54c622f6a0a65bed6aecc84ded428a7a6b4c55557fb64a0300cac3af027cde3182ba101ecd57397eb2fd06673adf941e7dc64bffaea8e396ffc70651b74c7dd378632f82440484;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae6ab31bc650258aec148972bba570e94501fe5966f40be2f20e401cae5db964d04118eef8333456ddbd0fe0d569cddff88d63e0a617dafe4f4f55583e21c1fa90df3a9bcad28ba84e1000742ce556f52b019b1050d260c908323f784cd5f2639be119358aa524971c22608cd2109c83b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97f895a05e6fab8d23c4c4dc0980d4a4751702bcf493c7ef771d5dd6719ba191d80068c0f56bb64f0a08ec1e815370c23b99efd4f753ae0802c3d9328847f0920270d8e29479ae56fa377a3e11eef706e4572e234be690add8ddbd71036e3bb5a1aaed3e3e9fc16535a34a54363e3b9ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17be75bc5289242aad882fd2e066f1cc1fb8c1cd8eadcb70c178ccedb9d77208439b038859cc70930437a2b0775210739a85262b14098316b615dc9c334a581b85c7d6606405f1ce774ba6651e9c2c117ba5b588436619ab5a4dd4fa91450a3d8f8466f058f381e42f1aba44e582ef71b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8a7c13b4ee2ec1d17bad3f11d1e37bee487089b6534d24f46fe65d9790235b5b31b3ca0c52b1c4a2aa1a63288c194317ee2ebddca1ebc8faca0ccfe3865a7a409e1a2b07e0b639aca3633c6b96e3f5537c0d57df0346b587384d610c694198bbd5c9cc21016ee1a6b434bc89153c8c66;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfeb19ddf426f09690810e3d4743842c88c341880e7b9b11a2748a18baa810a5aab0e08f3a8cac41facdb30269a824219d69f1c59a0a616a1d3cf53368171cf5820cabca09713e40cbc6313e65303a662f65eab1be51783aff76fc01a3e47fee28c3cdd21ec7b816d62b77f5434b31e545;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h687cbdd0e8e3c8b777eb3ec4ff65f1f593819f8f632fb021202e4d4cc8e720b1f2860191d1a8b26c820f6aaa90210b7a0a00e6a99753f27217f912d650b5e3add7d3ad3f21918e167c66c5af239b82a3da02ae8eca23e744fbe2f2521fead15fb144c16d47a7e78a05326b7a017248330;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hefdb37e78f581106378cf5268951c9ad8e28301ec8eb5892d1019525f658e206cec8e63537abeb721883db984d5279546ec81e459b6b711f95965a3383f44fe340677507d70df52f26adbf1317ea1f0f553db3b178fdb8eecf9ecf7e7ec1182ae67ab5edd5d7323ad84347fc32ae5791;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8cdba1a123296748cfad60d182fc26ec739c386da8dd76b546a83c60fe1d59a6bfef6feb45d859e5b29b2e720097c17ec04453da28f32a2872139d97bbb8a548050ccfcb2bc5e9caa7759cbe58a4b6b25702f8d3925052659071dfe94b191c162e201830e75138b3f6cda82140975473d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99fda6f73310fe1fa8d07fc15355d58257952b68b119497942093186fee44190cda28ff47281a04ee5306d3232a1f001b99e94ba687f319f3423112bda17b61cb4611f8adc7d7febca87a514024215f2e2440a1e7367ada48e76cd2673ecbe261f92d039c5c86e775b77a8147d3ed8c32;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce58d8869dcbfcee8c54f7bfb4d16a04a3e1eb96ca9a1092a9b4be1760361445715b8e65f9db46bf2567c10d9d8a95af635872c4500c8b0242ab3fd1a36481ac03cdec6c2b7a6c5c80a8b4bf5e0516f03c778d29df9014d90755f4fcc717e53fd7f7c7822022e857592631f30a0d3b914;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75edf63d66167e4fc18498c40204dd3b4490f80cbab5d6f61680ebf83a0cf16c2a0e29a1beebd8a9ee96804b1501b2468c6176d597f52f04268879925a1a39a5274406ad75b9d0e628a8a89cb601f97d29dc828c5d7eee9d29f8c32c1a9dd0c062dffd522ae62c12f6482238453ff1fad;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1541a1b2154bbb013036261e062a312e3ba607fb942c98db5f750fe7ec7753937a8aa9cbb5192d311b4a8a95f94b0e2271eadeab0f793e4111739425b2d2f28516fad032212e40465708f6757c03df6ec4fcb3996e68f4e2ffcff7554b16d0a82301a183dc31e21eca0858573bba41d5e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2bc5af97622192a37b830f2ef6f2130a79bcc3c55edb944f4f1b0f6f746c3fe599ab06c696a312b968e2d31b1f1003d2ef8678f18c73663dfffa35836edfa72243b32105b9df496dfd7670fe766ed8cead2e5e0b3a4b8512a45b748bc1261ba92cf88bc819ad715689de9702bc37b76c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hba0af596ac5c99b31ca86ae11c2bf644866100eab34eb9be58fe0f5903d7cba1711eadbeb5f3a991a46c8b2fd738c7db7b8d254414fc1dbcc7b2af3cee00bb92f1497a87dea9eeed80d6927cffa655d54874f3ec375769ff83b12d55b72611bd30ad300f253d2bcfd5f84fc89036cf0c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1a4868fd92c36d0adef6a3eedc295845e476d1fe833940f18080dff1772620557a2dc2daf8e804044e61c778ff0f381aa2c5adf26879318606be5cc5c1b0b95e289e8a4d84e7151bcc748b99d81a29ed1cd01a0a33e0dbe93715bbd0baaa71b8bcb009e7695bef5a43e9d7d14ca472fbb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc1d979f4cbfca62481fe92e4962a9137fe6680dd468bbf4fbb56ae5caa0fbc5027d38f89f406cfc61d3be5c0eed8d78983a1e1de7dc15250955fc52e183fe6e74be02c1d3aa89d7249b8d93e4f579696ed9a9e675c99f5c699d4d5d5cee63e93d74f5041bc0ed09b5f500abb886bed39;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c45c1cb3e83f5d9a06bae843d2047f53d8dc02cefcca48f91d3d7cafb422ff201e7021b7b576fe09ffb3ae60fa7216e3a5a67e652a21ee71587e197c6db4c8ab2fc50394b2c40e5c188126be9cf5adffd770ec97ecb686f6e7df60015b48ae4a1f5c8fca5ce69144af26e60d68008854;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd39bb53668a4474ceed9d3a81b4e0064de76429af0650a2ed3994d558241f8a231ca8fd2ac216e3c02226c3560c766a34787403948ca57ddbbbe5401467d01df921006152e3e628c93ae8fc4fd93443a20aab30efb16d65b6932781ea71464ead6a68077ecd0b93024d9179f26bc393a5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h689b0e523940e2adff4d0b1ae56fbf9c2b8b9541b22d4be77ae62cb8ea8873d77945b3ea81b79efa061c8b43fda3739fe2bead2c370caad7ee2dd6f5192fd09f2e00a67061d3fedc40dc11bb833c05de413b52f6ff08d99358b23ab411c6c4eb595c7da8baff473369ed01c9e12cf9fb2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78d0fd97cb5a6659c7e98ccaac1bd5f49d09249220feffc6d42285ff702d9621de9531b7b2d2fe5e36fc7225cebff31550bea383195e4d9dd2de297797737414469e732a3e54e69dda7d5e3823ad0f1e413a6fd37bb20ce440d99ea162e0731ba6412328201e09ed417da5e4c324e938d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h79d7994064994e47276de7ef1c3eef87d96a671ab723a9f8dbed526ac502133ce3670ba0006d20d05d41be070657477677c508e47dd09c8129c62f884f5141eaab05f0181f349c54e2ec484419d5ae132086a3d1a65dc576356a605b9854b3f6a7be8eae60357375b6c98da6ed38f6ecb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha35fb688bec017acad0b3c26e5b15dd3da348af092821bef815d56396040b03667f665acadfee4fd1c663d27dc90676ec49ec3f2fc4b25a969aed41c1e1dcb4ed846be83b199c77efc41087f291b5456b85ae431efceecc78142e731dc898cd633d62293fdf03e5dec586097db8fb922c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd44b3ca7577b89feed2c4abce9394308997ee62dd2dde98340f9854d84fa60aaee6246a3855ae9f05754c05ddf8c10f3bfb0b9d7b02feaf669a1c4908fa70d04181f0268078d76c5fc1c04df2818b0f20501e05b2400614bf2476d86ac37822c495836ffb7677e1e075d5f4d65563a6dc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4715682df768417135793a77798a63cf618e425b970547cde5ea850e77af822fd84201062024b76534ca1c9dbab6bebf74bddddb944e326b16f22ad62f2718e6630152d73aef3889445e8482a8c2bdc615733477beae305a1536fe3079cd87266bc2d315d201936696a47d32dc169e59;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78bf75f3d595a6bbbf179be2c0ed4cc6891b3beb0d533d6ecf2c9ec49209162ee560d7b959bd3713ed0fefb1493d23ab292319371ef87b8e7f5e58619dd23c904460f6586fa397182aa1cf28ef223ecec8af3a5c0303c6353099dac02fb7ba3a0a7bf3a8395b3677ef435abe4b5578e70;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf92ca561198a3f4ea9ae5abd7edb9953aac6fe6c323a9e23db757411f3be1b3741a3232cfcfce351753c012e52da063363fe9f4d3c731a29c150eab3d890c80f84a58264dfa6bf27831f06518516b0545db978486015e6868af0d048e5e3df9c85a7da4668e95c05d2b3f607388784038;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6eca6087073f880571b092630b273d190eaf278bbccfec6d018416b629a3073bc90258c2c90a18dca9a95f88412fce3b1779837e68771826d277d39aa4cb143cf04a15bad1b0a4afc59092239945858e9f1111881777fea2e7349dc7539b2c45fbf3d5101c43edafc5378610a9e49cf4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3cfcf87ac6dc982a92754bbb649cd6bf204f283fe91a0a065a22f12037bf4fdc1e8d13f5519169ee68ee4cd49735d8b2b329992c15e4ceb7dcee87c3852e2b1f39e0f808edd7165755b3878cb30c20b94fa1eed137180478d32dbcb3a286e907747f2c253f682b79f94b762ca6484e319;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4d4d211d058f6e6aedfae5ad5c043a6d9dc0ad5423470d831ea265b190a3b8b895d97f6a082378f6244bf340341caca87f60a3e7ac46b7cf3b45d3d083ddddd3f87e88e40366f3d812d5a75ec2878759c80d6cf041b9e3922423b3316133a3224955f1f869fd07bb67680915bda237c4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2efeb1b7794c3328b59e1fcbd1b4b6e6a26745d901d5532a3599e9132cd115ec38f1868b46c62edcbe4c554da125fe1cc016b7912a62296878d08c1eb686b1ccebbd7008c02caa012867561fbfc0b69a31a7c493af4887c2a229a2c4ac9a68b584077ee817c36c2cb6a2ffdcdf53bd970;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hebbd21a9f90a086a0cb70a38350d0ee3e1e6d1f9f3990d2af92278fbd5cee67862f48ea79eca8490cc79898608c921eaf9c33c66d995e81a976208aea62f0b36d0d16df4aed2a1a574c068039f19e671ab8e153e51cd11d54580dff49612ce5b0081d9a87d93fee3ff002381d45347386;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc53fefd7631bf2f8627c063f5dd7b05e2f7a21a7287e20a0654886d9b6fdcabff09195e6fceec9686610428284ab0157a3b30a6b3c3eecab6261742afabc5d11c9e8d2d557e24ef1698d958babf448a66cc2df750ae7d25d8a6eacf986f3e7cf1b2438cf8d4f852e42891b1b62223f2d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c71bc6d30e0236d2e65c2a1a7aede633d65bddfd2ec65d40390e2f410d5054d2ca9670b1f501d71686e7d9088d3cd4d990e9cc87726b566d29173df7b6d0626283eddcf74ebf52204a2a056e0171612653bbfaca5c5d5da565b9f313b62158ae45714b90c2735d278c7c124d8e346bf7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha1e37b10c939cb1e753a32a1817bab20766fd96ca77ef05127fe669b51a21af11fa08a745d353f09e6217420534fff84f4c3d4755fbf78774b0b3b90383cf0208e27d408e80388aa62b5e59c7f45ed32122023e555db14cd81dd93bbbace086201266e36ce7230bfaaf91338a571c643a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92cd3aac4938ddf03de56e7c8784a320f3a29dbfa4edfbe1b14764e4f9f5ac5f10b138872c464819005f2b73e2db28f98f705ed6a06e9809ab19a758caacec1d3ba3a6587e3036f1d54849a2c75ebfc0ea2bdb035c80d8127181af625930e2613fe9669269d736b3aaf20ec9e6de057dd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e889cf3a7ce689550ec8e55b2cecd28331db253f5eebe0cbc1a38c21ffa9b093a5b9c59afced6795e2e9dcb21ddf61aaef08513da1c024f9b16b926e8b129d1af8a512fc11a2b9d8f55ac991f74f16c454a04374b9369d4e1e9e362158db6676c1a26841d33fd6c034f7293f812feeb4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa6509e5d81e2cd5410e199236f3e6e42495342236513f8c94908ef97645c0202d2d41fe10d5e63fae44ed8ce5f96cac8e9eaa5c2400412c5d83dd6e4baa74e792237d54aab043bac6e11c0af59ed5f68b3ac1241cb06122b4f55014e2e8771816681cd229119d4ed5e43b97277c8b883;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf363af544b03cb1bb2426aaaa9d2b8b169d07d3cb284d19611b36b20f0da74597fcb8666d7c53754ee35a37bf56f0742a101f78a165ee7c4329c81013685b3ddebda57125dafc676175a12e1f672bd93e9e16a5450699efb198c585027eba1b539e3612d55e9504de6aaf9e9495c1cd2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb2a0d3a4aca99b54e6837b7df6e18d7922bcb551c6ceee2a2f2638fb82d8ed4996ff8262235b3b86909d82157e3360fb13e00b75d5f2df8b0cb7bdd85e79f82be10892a310ed6e79e613ee4369f2447bc48ab9d0f1e2de94386e8e38dc48a37a14a557d418e579589c9e691f1d942d3bd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd206129411e7d51f5f8c4d04cb16d2e8d405fac5d00cfb9a2b636fb4fb10777a9e4d20eb85d9a470ff7b8031a17c6010698e94fe2e1dd9a4f954beb955526e2cfa5fb67b05a181d4fcdb53844e9af9466b74dd558a2859dd61ac74d9671f36bc2e825159c1fb81a173480fd61e48cd886;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e2434a15d7e740c2b99781e83a1100c666e4e71456bd13c21d28ac4f201750e4f6d1b30621d172b81f9af6dc40e56a5c3a5c51b149a6b4b9e8aee81a69e3a2a5d332d47f818805cb9c51a143f7696b3175b7029c9b5c0b66afc762cb057b864954eb83ee6dfb83aff760fdfb14c7d552;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1a3bc8ed0562dd37feef47fb17deedd231756dfbc9e4253a321f370bde1dabd11e4c7bd44390de1ee5d1acbbffe91bb52924a9597569ccd7873aa884c18d5715904a65067c62f8d323b2427bc937aa2cc06774ef322745172ea951701e9d6e31974b42a9ba9262d4e70701d55ad1ce8b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71e0a7c626e652bd01f17b240bcb83025e8715eb9443af464699e1b6e684116bcb7adcfe14182afe1867f02a4f04f6c78708553e27af650a69c25c2f62063c74d4f090a60f416a1d55f7d74acebc8b8348ceef6ffe3401dc6f3e0a1738404c87ccd61f7ecb1c90979d4397a4d2cb83ed9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c526b2c795228e9ca877e1de33202a5c53fb02f4bdc7257429729b5c98b2296525e357e5f0451bba762852e868960462ec1e870ce0ad5e0f9828c2ec081986d0500f750c074e8d7b5b2a7e07b52a1dfa92c7183d8ed30077342ee093038d1ffba37324dfdf0868a11d721337101bf441;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8727426e1b11b224128152ebd792471300253ce9ffafe9078a74d4e0b358f011e8ee88a916c0f71edb527eb4a381f4a51f8ff6839ed1435ca4b27fa645959cdb185d569a3df57ec6a0dda1033db52ef44413a71bac3c6e91b2b342dfadd4a494641aff63ecb8462b361762284bf6dde7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90fe1ec48c2f43cb871d087103f936c2e9d3f5911bcf241b39f1ee21b9fbf6bf20b55b6a7bcdb12279be211c38d6e5f0061d1669111064dad7c9382c79d990a60d18c345bdab078c2fcc5bd3675056c42cc99caa510c314d0fc3624edc76df423802b09c50d890c58b1ab4654e9ba5f9e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d8b76c0a8b71d453986081ba9d908df6a7bd9f8aa7189b3ec2feca49ec2c1347e6b5a881270e16e8908976d3bd07ee4c46ce50c7c2c8bb3484bf9dffa64760ee04204f818021c8b3a064aab1a2e27b46b7ef77ace391a71c30218e5ba166af7c734a5b9ba884126e5ea22ef00114f372;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43f7679a9dcce8318175a16e2f61aa808a9be6bf8489c85c9bc4203947742e1188073638611e00883e23bddd60b6b007e5e9057f10515d6c8cec9ab9b3c0053d3c51f6cc7b68223477c26113d1bf7bc2cdba96f36e695bb64d4884b56de9b8c5c93333283f539dd46817452abcc002e2a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9529301be4cffbe6e8d6546a309449b253c9adc5b6f0e8c14a2cf03a8ec7dac1b0aa0e9b2230ce56817ce1c62b0343501b2cbbc367d76b95991d6104dca5517be66be13b70458b3b9340c2b034ed333281c4de592b9fa4a315bd30636247cbebb01e178ce322a8e88b2da38134dc61b11;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb63cb29d07e05798f0c5da72b7d6ba1b50499479a2d522e106266b66aac05a03b854f303c67f10565974786e1f9d1e09989da693a8c1321e3e709e0916c54e8437807e366455dd37e6ec6e84a401fc7720858bce4f548abf5768047c0131ea28e50a2dcddefe88ac753a44a52d150bd7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6010de14b491153febdaa4af1364706ee1fd303e249df39d4670906297b5701b41d2b9b3b825769fb43cc87d6e08e2d71d21eff1fca5d6a3e81b8fa6cadd72c23caa2fbb138c36fe0368e4102323015898f90f66f5b68c91c44f77ab8b8ed7cfc5d57a1a9249c1e64755b0e7d9c198f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h147abeb5205e5affec327353f180d1174e37b68d5832fc166703cc7c97e81735424b8811bbd548c7caf4dbc57d4ff76e457a6a6c838a5060014f2c528681952af99fbe1deeebf23301e4e0073e82b162543a63e11391c07f302164ee912dcc7ceabef60f16c4f517363e3745613a5c50;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e0fdabd29d21da0f451b97bad8429ce14b2b57953bdc63cf0ca3be981330e79ef17f6a6331a402dfa3138fa2e2bf3b800bc3a5fe7041c795d426422f5530d81b835ec39d95fddab7f8e8ac2b303d75ab90e880e0f23e27c690ab281e8239fe1df890dc6153b6296382c6b559aef858fd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92f54a91724c5410637e84674b8aa57f1695ab56dab7f3ddf706544f23a3896582af492c7640ebd198bdb20cc0a95b447e1a702c526e0eadfa73ec10a4222bb3417d88d8456bf90c1ed8bb5cc7ae206428f430134aa0184da5d1874471056cf1b9f7f018d6ab5eee4823b99a5a9dc535;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a069d19527b870c645d0218e12edad23041ada6094afa11605cad5375ae99d1a5c122f7b38f4bb1ab2a34be9f7d5fe7d55c3dc0db67500332c77a1869b9e0c89b0cfe5d8a3f6c4c3e8be33a90a79036b959c91bdecb2f3b3b0d56894a05e574b98e3b858d8d762714d53c32e4cebac6a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c93ad9d47ac20ef574df4cc00ef8f260d50a2f4efd9615f3b2c48d467439d6b8956cc76a45bb60c5809df3b2fc2ccd2054de080454386dfa7cde820942a02d933be0a2d3b6c5738e103a115aa170dd4e51628afa7a3801d4e281745114265101c36bee5fa1c598fd83e59d4ec21859b7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34b78fa059b2378382785bd193fdba9303c5058fd867e1c0206ecf902ecfc948c56df714ba3236d1d2f0b440871d60db9dd39d2c00f63f321c458a13f4f794cab45b82578e35cd1759d75d8630406d0579ef9edd64049b5265502952b434bff0a621c31f4b6dbb55c7cd5db1eecdc97b3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc85ee2c34a8091b8444fe4b8fc003d2826fb635ff641ac5b1c0ae44731eb24c3d2c4327a4b59b46b8d1bd46bbbc59f3bbbe0cc3ca17e9a4e6652357df80b8c75fb5ea3ccdd73e4cbaf7f4432e1bf5bcbccb32478048ca0a4b940b15d42f285399d031799525971839e30ae0d49081223c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdcc542c7278c2f83c91afd2b3694196d5f22fbdd36eaf185bbda7b85e8cae6fbe0e4acadf65d7333ca860b026969af9839c3d55b7f701470f18d8fab6fdd64bcbcf636eb8555343cd4da955f31df8ed388a488f69b34a3a31487175490e1af02e4ff0435af65e0ee4fe8ca6d642c25d82;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he4cdb1b8c859b9a14349a03ba2c5024b9d1b619a09f6f3e5b315d549fa64e2beeb40244cd4c095b4ec01bce382fb525cd1de0db5f4d725025000be81000756329f4d00c13fb0faeb8dad8f1dba2bf119b836d446d853879994b9a9c31c5cbef682b6a519f5520289e4fb5844fadb250bc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd87b055d5b3efe1fbb446434fca4a0dd0297ff6e844f03a17939d7e5de95b772cb3c34628e9998d705414468d7686429a7e6e6b4edb14a017dd46b9e93320a1e4e4878aaba3456e3ee9cfd26965d288e64ffb3aef47ee0db6bee045ba7c26d83fef53205e5fdbf076e5568d86e312091;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb8ee4c99feda959d5b09b3c48db261f934f7f5438bf62a65fab8a987a7b72f49c17f0ef0a9f8225ea558c3ed66ac0225fc18d3c61c17e4ae114e3d168e2b8befc58cbee995c709fdf300d4983fd3c6f81d270539a1401274cd49c4759c1bb91a22b174521128fd79c0194640beb35c36c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hecb568280150694bbe34f022f90b873e4764c48b1d476164eb25df39b1995a9c560df648dead09802304e03b55c14278719546631292a40cf3ffcc27a5f4e5bb3cfdcd139e7d6ad3428b24820602da262117f472d2dc8cab2f7f4736ddf9717bb109c165d1e22aeea35bc2680eb81ae5e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8bc81abef3af2eb1f996757aec5de44393ff682917b4f43f75415980f4898f283d33aa5e8ce2d4035a6f6442f2fd6f4234fd8e401a6e0c232973a7fef76332cfb26d02b1a50f416a8054f2f602c83de57da04b1df409e7b505af3b28a6318068cedd575d0f379277f09d04b89519b1ea;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd693f65e4f402a813b395abc46b527b645da60583fee6e2d14cb3ceb3201f7b7f591d67b92d6b18578d99afcd27752e520bbd3266033620617e155be864ecf210e5320618713ed18744d55937ceb8493c4805d5f15e4374200f054e54ba3f2563489641c107214dc24eaf476b84f9def0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc2598c09864be2337050f36a717de2294513665c953f27d84bc6319cca7734d497353428ee913efeed149515bea67588f52d5a8d82b9f965f4cf7c9b76b0d31dcdbe1958550f9aca5d76b953adcadde58c2bfe52eb08ecd93cd287fd1d076e23d8a566d1703be98712aebbccdd435da5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72a48764f4f951b315c0c69a2ca5591b1e679b88a2eabe365f52f7f38fa0d3eb2cba82d41b8da855f3942e9dd512e92347512662bedcd5c051a6cafb234ebd560e3e8a25d6a55884a2620f77fe761a34cb7aa93ef9ba29ef5d891e1ea1830754558a735aeda18bdafa328a20f615968e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1455576a04431f2eb09889161b7abeed0d2761710c90d695686f202de0e8ab73a56512d2f6ac76597a450e44568a63c63b2201033bedd0bd5ae38c8f6982194a94f45828e7cc05ba977d532f5f89d12d829337c3b4190a9c8d127d811446c72e84526987306315457e622798c0b2d00ec;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1db3c2e8955eac02515dbd51c720fe3246c69efc13f933c0d51447802137ef197ea43ccccc07813a8f5acd8166135464c9c0c7e5bcd2e3ddecb0724ffd63c561b11056edecdf090716e5f1c40bde25b95d75f0a0b34ddfb6f3854ee67c5cebec8cbe5ffbb9efbdf416ee84591a581a433;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8afe46c6f63bb3fffb7f6d2ac9e0ab7740d3459a316c14730334464f6130bc93030b4c021721a58c92dbebe7ea79bd5c5dc1d8eaadff7e40804bd74d88d73749a3fe0f75f6741144afd0b932561e8253224e9bc42f26833b052685577482c1d8723d656764e96d3ccb30617ced768b0c7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h15ded9b808b356e868943a2982907ee5f357e506596780148fe217e8b9de55a002f503cf302ae8a4d68fb035fd1e8031f416b82a57e0485dab394fb47b305d0b606b167bbce76a84dc885a6f5498fbdbb4d5441c6deef3610a8b6c08b8ce759e0fe988b368cf28a136d5a3bf870a12432;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc537587cf2fc79cee1cf56774765daae4b9406c7dfbe7e09337b220081bffaf1c1684296d07f93112df679b245947b7617057c6a65aa728f1a8ca7d4f86b1f878e02d72d61f8513b4ab6078613ba4e9ae2694c0faac51021773bc16e64bdf6c30ca68d6206fffa4c61cdff7a880645ef4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4d3e10b95ca67dad8fadd5d85db90ff4d5384215a6a8995afc7afe73904da63863019070ab0f812eca9d7eb89b2d5a5468ba14edf883aa9f384a58215c420919ea3a8d0bfc73bc272a7cf80de0b5f02571d566cc566d90d095d71f2c28693e100a65220365f6230165c84ec7f579165;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ac0a4d6167db9e399db310652bccefdc1fa37247667cca81a9bc9cceffa295ea55819ef8ead128ed5cc193c8cadd5d700726664f16b4fe3b4f2792ce4c7e86cff1b0a4481a70cb2be47395397188d1d14a6cae5a100e4e2a69aa56a7c0e1b4d208cd94da6d7b45e1ca37f9b9c54fd287;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h520e2164d2e603a0a6ad33cf88add4a36fd6a2149f011af90a764750566b9987e6778eeb28f5b2ad4cc28b0a39beec43579b3c3359a4ba4e153ca000e02542f88571d99d68efbd277b416d2e52e52c788c59254f037a634e07f6f4f68f41b762b2b13190ca51b34edb8cba0720159cc31;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2c5a8bbddaa18f122eff61e1964bba9a89c983e40802b84b41bf6ef9ff885412dfe5f4fb48de233de361432f384cebc363e429aa758f2ee2082b21fd8de18acdd79a6bd0de201a4d6d58f3caa47482a82423a7395f0a59275d1773997f332c846100984f2350d188d639a1ef671816f1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h690888285dc288f6dbc965ecad456cebe03d67be40fba425594dacf0ea8ce93d0238722d06261e6e19a66fafe19485d7ea109e848fbf23ea204daf50733dc71a3fa71be7cfc465b402dcd74285f06cb44b1c392e2532558e9f1eef2733f988708de377256301b45588c59de14c5fc2a8f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69493524fba6b79ab6b47104b78dd0600083f200df461f36fb28f37c7f2cc5b50f46229b96f7f8dc738d9a7c85b9dd94e663030803d68f5641f96d6836acc81e48187a009b2e2d427bb12715883db078e9b2cc0256968c8dc257abc90afc0d14e8a145c85da55d98f1c6ecf7aea221c2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e7c2d588816663c03b16108572e2106bfc0c2e5ae74c662bb430fe9e43c05072a32697c2f00f3440e3a88f318c01f8a53a95a64b6827e97df07cf646a7e445b70ec4c1f6082a6f9b42e3c28e6c8e2557240aca79b74ed22239c18eec1085c22a53c68685c66c53e578a3a1ec0722d18d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he957c7ff11b285fd400b139d509f65ae0bebc4adf1374c5f8189108467ee0eb5e4fa3fb3a4ffc9eef1da5f05ce81203fdc802341e6ffb6a48f90ff026f6b779e36eadae3116aec50b4338f73264d467603ef6fe6de48fbc29b6879e6928b94ec4dcc654e090fd209699a3d546cc40579a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4088bb78df58f50c5c98545c8b6aada6b694904d4d8012afece2adb6f5dffa7a1801489467dca431883439b8cb738edb98ea9f588920d8c194d079c9c7e4ed8a8e9e9ca90b13f3ba8bfc3c8dd7d85b73cd029bed919bba9f69abf34a213a55e1e4042f6273e7091479a2e075a49393844;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c05c1e74406c86c3ea044836e87bfe8004b76ea0410d81f635dd575ebb3ae9bf39c707e9b3b1b83406fb3d533d5dc72c6db2102e07a0d5d5b22d4685110c00728f1cff572dffba53d5088cbe6f4f655c8f44ba379237222e6e01dc7f15472f5818f0e19a9adadabed8964aad1cf2dca4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1391945d7f4771d1ceca6a55a229da414c3b1ce25b4271fee17de54859c9a37e3955efb2707357b7c63fe8549f30e28e81d9482fb62250ca9736e4054e0a12720519e62085dc975f968e1680f0dc47d805f2c4e088a34d09253b09a6a06cffd8b26e63228a41091848567a0ed870f9897;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5bb682d9e02e60a802ff76fccaa813e3aa1c77261408690a0d363a45d511c32de7505377c636472efe8125c06ec40334014be405fe4bd68d2f38eb4fdb94acec5ef4e213956bc7f2522cd6e5d9e5fd9595fd1bc4b289566652dc7daf185cf622832ae262e26bfd9d35dfbffbcc149c66;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2be7e1e0d8bb1e395199a20f9f4a9b0e4aaf9a0d10281bd4a849fe19e7895a8b66793e2fe3e85daa6fa2bf54b0e3085258336d5a98bca1632768f5e70d948e49ba8865ba4ecad1142ee58c6e12dc13e32fe6a71ae79ac26c7ccc45d6b85a0b595765159d9e75b4e63f26af778f3da59d0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1a03b3fd5dd560d149acf45c6702753986710994282cf339ba45a24afe29b2bb2361be33a132cef6797b57c68167a749368f3276db40416e077047fdefda12f6522b39e4c8979a65f700f79bba96e1fc225912f91c55b9807e8cc38ad3666cf6d12e3f2a225410634bfa63cf5ed7067f0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a17a05b8044767b0b033606675dbe6cab7c84df65b1c11ce8e052ed30e32d2bdc6db6910b33093bbf1abe365d3c8edd3ae0e83345b94d3162ce1e486a1ff01f20ea97d3d57dc3d64d6745f7c9b271bbb5d63aa50e173ded69a0a66ea5bee50cbc8a8f113d98a39ce339a6fcf626a2c58;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb8e068ca78b98916a41d3c43aa94f2ef925dbcd311c8dcbfb5939d6aef57bb2c87b9a5872ce368993ae34d2e16e97ed623d019477ea8359c4f08e90f65a8d4c341702926ee93f28c514371c0125f89573290980d98850a103b99017b5670026a3b6665fa8bd3df4bcaca9d7e83bdc058f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h206be0d40e0b2272baad749494f7dd7663305174ad5c2781d369f19fc9e4529e23cafba654e31b0d7d1a38970af2562bcb8f53e6cca9f3185f94f416c4595ca83523ed814ee226f50fdbc44abb85509935a8ef6e0ac4999ea3af57514b2c582eb99bc75807b042e899ceb96f5cb920d93;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h804a9895c48acfc0436ef318b9376d3104cbabd7aa583a5cebb898d19de5eaaafd8194568f60da9865b6ece5d34a90d8c0aa2d3f877831d184a8a8534a870edf7b8118bc6d29a7ad0a4d6a326f2d6094cf83010656e84fe722e7fbfe8f97f5e1c7338fc4efd629a64eaf2767cc2e3721a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hecbc28d8a833204245cf2f962132a10c7804c76387f32d17181c973c5476ada420be61a3b5c70ad43ed143176b98e5bd77f60187b28e850cc62eda13e935972cbdd3e01bb559640ae704da7579a36d0151bbbb9c202b6ebe3704f7f829a45afae0ff1bbf2bcad8124908e1a674862102b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2be786dee16a2367afcb3414e9631d224b067a3f1ca1daf1cef2c339acdb60275a9f8999e8093c6d19400116c32d0034432a7cfc53e9ed0c60bcab4dfebd2d943bc148a6276d057f1859e4eb8c344becb0db3e55f1d48e5d98352e96fbdff575b51e3adb3c75a0cbc638ad40938fb52df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfbcaf0b4206ccb1ea5f811352427b1d8ece44330e489fc82c253015c150ede6f18c392a799ff7faa7124fbe45d0757b13c23ea06849e1a8c7d9b1f4038435ba2617c9ca3e450b68573b20a120cd377ca3b419d490c911f3ebc1dbe898ee794587f65fbc1f644c503b2bc87abf10555275;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha921f8c6387473e03d923674d0b30ad7668efb180fdf2b1e86ab8cb95f1ad39f831c3907445c79a238df72855c1429cc19a51e0c1dc9eb94f44736b28be318c7383f0b3c847b3ebec3d72592d237428893eac392197d9cb445b92005f496ab20ee879b026964e2db262e7ff38fe6ce6cf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd3c1914113f866d9594489b01b05e32bedb0056d5c1e045769edc490cbca5e1b04bec95b47eab3565b3ed55e66fbb10b65497476c46d999e635d65bd8d64042b3fe004e8c180ae50e0794698f21be8640a8d5fc6088ede5fb365cfcb97048f2baa5134d7bf7051b0d6ed36bb1fae52911;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haefd55d899b2f3b6363134d84f822a1223ac1987a8c537441265beb516240a6a540329b6c2b11eb2cc2c30cff8940def6eb7e17f02751687f8993b326e83988b43c31bf6f233c13f685143314e00f06305c6f564538d273f6671257735ab7a3fb40039118fea01eec730088c8646e409b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57678e3b21a913493043e0d11df85b93346d6c6e5763f439b08ff22376cb946bc247b601c7d762c8493feb49992bf2cb53fd980c69faf7fe5ae6e2c2f8e5ef83a3cd2c6c6b7813fb67da46c914ea7c494bdc270bfa4ab5526beaf399354526eb989e6d66994d3d98b7e86611ad78b50fc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69cb231d827640988fc17459fd71182c50cb1a85e7ff82142be0227271ed2bc88b3435533acdb5378b9815ff9317052984cb981735983f6215aa45262f8cac98e0f4e89ebe551f6d815bd497c482fc87d9a56621e405241d5efab014a1e663c7f3738473b8b540b0a62643b0d67e1fb5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf803d85b0be833d4c667e29a03567b0c185964a3b687b1d4f3fbf16defc61b22cfef8546d009df2a4374a8e516c227bc577cb42e2d3866175126feb3c1ca447473a573ef7fc499b6eac19567688cec39311b61adcb0bab3ff5cada48f7ae284d5336c6810f5c743d12246c48aa45f7191;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h378970a1a19fd4df7bde04c2a29d0c4882483d0dcbb71cf8740d79c7a814cfd34cf48ece4ede4c598077013557d644d21a7d3d421f5bb8e1b4c0e007f4eda2c5f62e10469e2f48d1169019bf89d2e6712f5c31e3c1f5435915557f6777f633a91504750149513e5dcd2112daadd92d3d9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25d4eac55af8702d80c3a127770036997ec554a41be175e898f34a0e10e6a851facbf8c316a3d761425bc86affe2db39af8920c8cb1ff8dfed26a262ba93ac92c8fee27744194f1b0876b76b054dd30ff6149be354cb2e9d3f4fcea8c949eed28c09a12c3cb114b519a66029ddc62460e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71c9364f97f46f502701067dbe47daabc1aeea6573fd61df0917903cf7970c12566d4fe9e26e2486fbb68f9b114fbe06fd21133f7d39f1f0128e246a7742583043bad3781d06c2121db41703443cd2068eedb400fc81d7fd346bdb2cf9f332eeed005175e9c087bce4a4161f7d62bf946;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h622524e28b1ff542fab6397327a11c7b3671f07e919c781bba3ff4c03edf67e066f1a32c19ffc7ee2f27a58cc3d5c49cfd3002a8eb8d978d1b27454f88fc0f5a5187194b96814741bc72c6fc4d70c92a312e25619ceec6033c95811424be346ae01bf6dc55db7cbf14664a2de5cb8a861;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69ece7700b8babee95d82cd5e5496a518d3a7a620ad9f28741d5c508caf3d3d32c395a33846816bdeb6004ec5bc4965868af5e0c3a20b5f1e55d7d185f63b923d956b7748db47344c722f75a0f67ed78ac1dbe08b24e4ac89b047d589c2f9a307c8c49bdb94788eaa789640e4345ac238;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hddda7520bc3030f44e7d7c9ec1c3b6ca7ee8b58c11d959849e40e18e1fafc65a6151ebd2d7e1e469b8073de33363e14b7eb1d4375988c1bf687d03befadf27239d760581fc34ff687e92a9824e2ca32c93309c01ca03ad634b2af6be6ab54021616be2b07c02d98fb812378823c8fd936;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8bda3bc2df65ded64830b827614d7e1b0b0eb5c7a356c01927a0bd208e40679f2d0285c4b1a4f0394b789679edd09ba9a0fe016d37f099cf9eac438bc5718c44836e52d2f23d08a36bd6fa3f1e746d10e81a1fa94dffd215371c66cb83fb41a22ae095dbca7da5cdbc000be5989dfb886;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4814dda87a16d773e5dc6f6e7ca08f9fbdfd9d760a5cb839b8e780b7df418f9ff923bafe648241dd65ce5c1bdf0a60cb5e1a037c9b560a310754b6e51470f049005c32a76f7ba2956d79fb192219f26766124c8b9f1032b1f0a75ca49cfc0aeda92f6564ded5a6f51d2eac4ce988d5423;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h620f15e615bfceaec609179d8bfc85e1f22346d77d32a100ebda986c9283c31433861be1e7363864d3f7309909cdadbcf171b79bb7002d0aa2ef8c73003e09f59df06e088e8ffe9f2bf490088808538f45e36f509180ad3bf068b43a22200549a90b635aa91a232cb71cb142a4882cfe2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2c1720f03692162dde0ea6f1055ec974e1bdcb67f276015f055a411b2f5f8bbba05567d8e25aa009ef9d15568112072e79bf69b23c3964d3a978af3c40a0c2886051e417446abe7f1c9eeb9b306a2f1e49c20997c0636e852a2c4f173688a288215bbb7dc4ddbe6358b332ac77ba86673;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h35642043934c18f7f91bc07867f854b61a1eafe90deaa96100820c48ba3da2ce3e5e5636cdf01a6e82e67f6cebfa25b1dd452d59d0a838c07f3c0f6e2442e9782370ca3b14ecd699493686cfda556e58b92a481100f408ed54cf67fe35339c18eb466b288077af3e949624324fcc383a0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h696189ab05a5917f6446cb7c785d1455b3361ad233c9de428b5f55ccf116c5463715ffff1e670df06b368203dd6c1135731d0fd838a0edce736501ac1c1162e7c9f87e636202a52abb6046f58cb23fb9193477fd88997728e71c421b4f9596ad8e0659da4420513115625d194cadae501;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f4c4833d314071a3f9c0f74d699bf3dcc1f0d89535ec12e25427188628b0b83a79bee632b4f8519ce7e22c1aff8689246d5de0681dff601fb50f1d03160c905355cef9098fc4c07d82272ecda026227cc38536f0a1af550269c25d85cbd891eda6eaf40c6ed4a2a8803b6f4e7004f628;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22574e1e627fbd43447c64b009b959b0b5a2a3952e4f32c48957a146a27e47d04fd10c8a2ac26d0ad2afa53a0758626c8af850e812728559deb0b1cd1f9555b17cb41ec57940aebe0cdf1cff8195983ae2a3793ed024ccfde1c94af0315b8fbe5d0c458fadb567b4188bcccbcff902dc8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc50cf078a096458527c020a2ccdf64e8a419825ed073c524dcb9ae069f6183d8e1c9864a6a6a18cf2aa78fec5c3fda935db1ffa1a0622f92d73448d3367140b8f02311356a612fd093b6e25700b5f3f6a0ef786d49f8a13f8bc03540dbe1fbfbb00a8b9b740a0d92e4cbed548bfac24a6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5d0b8f4b59652193d345ee02cba819bbb9a60560c2a2b47e01b49d37c2e98af7cecd0290b9c4d487478fddf0f70576d8b128399042fb4a27f5e440457e43ec4dca5986abb1f8cfc5ebdbd84e275e4a755cb2880e7d818b2ee485c44c914f765555148ed945dd5b798bea4980782b9292;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8caca41865e507155f113086f4de9e09e6bfa44f70a5d4cb804a0ba8ac20b6255a80c989c04f2519e592e1ec0d8dc7413043626f47a6fa465786a78b34ad4aaf5f28ced8d33535424a4e5554608c4263e2a3c7344c43b6428cd6730ce3710729627dcfa05581d5cded6bfd7d077330d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f8bb5e4735f6164f05fe0d7aaf989ddb09e3f68cdb58c477bc3f1259545f178d4cf8facab28731683b24e621a5110b7cd65b012ffec1e2a6622cb6001aaf11b3a4a8ac07ef878479312d5a1583743d2555d5ce8412869395569ac454c6c10eab28e862955b3da1ca3bce7ce3aa8699d8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbee48f6db16c47ca6575db7e1c545ecc2f8293edac1ca6ef7711ff3e74c939808265d42f310aefa3d73eddcf9a7f922a589ec8d81bc7da7c6501bb90c0d3a15d3deae1c52b83b38cb51758fb7059f854725724ffa4916bce6d3b5ee36be433304e493fd66137684c259e5f7bd97fbf81a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54c28ea054ac06cfca43e9be5720d8abfe671e491b6752a6f7aa87c0bb654f59798d43a4b3cc7c0267137089017e4a76c506ec515cde132def4ecf482c9dbff798165e30c813dd74d53fa00c8dc556774da12fffd950b95f92121e502270f4c8f08852f5ace31b77d70014cf176f436d7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h428b992d435cf527d79a108fa07cd47790d9689fa272442906963a3b9ee4dccec44ac16caa61958fe67b1434dca12a6c7135cfc417b5d4160d06c6740f3402d557c3c5ac193d24dfc5a6d964e6aac8cc3d34da9bcbfeecfbf81c382d822bd3848e273fa73b32f1e9974a62cf91f259926;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58bd534b038289a53dbd0f1cfc3b673cd93ed21eec3f55c6216e06cd39dca91b37584a0f0b7ae7bf251aa3e3394a59b138d62188dfe8fd5037b7996eb2e4f97c643c90c572bfa71ad760f10306a4d3a40195c173b75bacf7ec843654268c6ab4ecca8661ab36941015da81a0565ebd134;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66e727c0cadc4b8f3d2ab3641c200ee5fc27cca88b560166d83255367114e62ac2ad008ed248b2e2e24654e2a38ac8976f1922a4f3f6fc197f0a9f1bb6cd7211d889488bfc186e67db1b1b303b02816d21749778ac1147cac74bfe26fa865b6cad93fde078d06093b5ce3d488331eaa67;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he09f25aa4a920728cca937afe35f951c4a880cc4baf906c17cdee0cceb4a45c6c08b31ccade68405b0b65238e9b33d2eec4c34ff2e61525edef938adec00195d97b5581945e3dc9601cb4e9ad4327d3f0c3bd7af779dffa8b2c054352eee9a9c3829a659a03aca2c8fbb69dff2bb2a178;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87ff265b87cc0c2d743ebf01056205f0e1fbfd69ae3d5fd2e85eb0fd71fd9de40a334b72b0c4fc318c739919639549774dceb0e410549c825d7342bf4ed6a3e4713dc11805c15be5694127bab1958f32538db0df448cc5178afe6cee3afa10fc0440d666741cc0dbec8d97d9ab87805b8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee39a2ad48d54110203e334170b716940240a8bc8e7d040a54d8911ea67337b2b6bf0d4bbcc5c443539558222808b3e0e2ba8cf9f9b6801809f74e9e1a602c05fde92eb02cd1987614ee30e30e76af10e56445e007d66960d318f5f0b078ddf7ec90377cc7f88e3d85255460af634b764;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc57413121bd5acb1db3c266f8e583880ed45a0b68f95ffb3dac5a0766d01df5a192a7f6f18d65251c222db5a172a8cf8c6e7926310f824caaf884b060a758802515ebaa028bae5606c03a33cdd83f3cfad881903b862ced4a9735fd6fe86ba72898f50f03c9fed0fbf1de2062832be317;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c692cdf27e934db8c74f964c1ad0a2633e324f55d58eaccd4afa7780901aca96d7b095ae699b2b733e34ea57600de4442160700ed9efc41efc6d9d3bb7b37f72bf06cc84863b4d32aa9263eb52c6ce50163399650f84b024691a5e518f556461b54ca4282d6f18a3fe9af88bcac7d9c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50471ae2ff93518c394b4868f305f1a3c3c9cb86262dec9b9f785fdb8392a660dcb8fa2b8f316b3aa428c1d1ee5bc4c3c2f6f2b30d44a944e3f027fa9a6711eee03ce738d71e62b3bc1da0e5c98dd8265045df95b8b02509aa992de17dca1480f95bfa3c2c6d4b06ff124b615029075e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4317faa164a460fa017d55fef8a0b1bda8829192c06954b6dd78279dd45ec64cdd0ce275519b5150c7ba9342b7bdb93209410e87f59c9eeb69761f791306fd099b62c6bff39fdba9e103c220a9397e8d274aa688679741e3c7448fa137fea5fb460fab8a8700cf697f2625e6c6fbdbb88;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haaade18fa90614d36094921000642e577ad8faac3cd86c779223b50c3f904f672b3c3d33df55fe33cae25d46112adca678b9c4be1956473e19f7647541e6127b397fa5de537edf1e2ee7b52aff3843e78c41f15c932f665d7579cb26cc5e14faa65ec3e344eb03c61b464d88f962bc8c2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc0d08d175efa739608d17488ddf1d75ff40e128b483a58a9830b66d0ad89d0f30735fab88e4a5424d500238f3fb0a1fc71046baf81bedee21ce4a6bef0c8e78db1311b211b155a058ca8ab964eba5010b932620049f6cbc5e9dc75a6c49719c11ea61dfba132ac84b7924717b6098876;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b3a943a93018544bfeff3dad06bdafccf2d27c751f9a6ab0926fa28b607740d1401159f75eedaf031757c2b3c3709d70a17b60cfb59ec334d06817b04ed7134ad1be502eb7962953f8f173dc13320b1dce4e1f39bbbdb0cdc62df5e1990b3547dacab77aa6669e9574d2b8318298400;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11853ec6c0cb6cd02a59adcbb6a44af167f1a37fddf769bc72426dd7def86cbc4308680d29a06ad993946853f4e5b04ae46ebbae9f3db07387b54d1b3955b090bc41d7b440bb92584124a9a6c41d3390dd063bc1c879fbf5afa83d308d5195672b105b2e15307f3d44c78787c9ca37cf2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d81f1f2ba97db6c26462d1aec9af9a97af943637fd312613275c593e00fd8aadfb8b07e1c1048b4135edb5482439a77762914edfb820d72ebcecb0107116a9d210a9bfab5faa5dd2624169c0546265a9d88738c857befc4444e409a94ddc99b41a77056e2f022ea457b3e0276ca3e985;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdedd1b582ef734226013b50a1146b62e6b044ba78c782bf8e1d4ed7f1bae017dc351c27b0d80098f657f63b99e098e92adaffd15e77a5045fca65a3dd1b00140a8e0a01c0381444f40b5fce1534687a9d2a66be9c25e4c437fb4530e44beb57f8610e56a2f98238bd64d7657086c7d252;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1445d1a99a7fc74ec44350bad9408fb80700c23ba648a373cf7d34ecc06ffe2ab9c5262af7c29319ac3029020125bb8f9d3314d94f7c118841ccbf2ae90724dd4b70b1b73083096136f16c2284039f78cccb8486e466fd900d0ef6ba032d4d2487f2dfea0f3c0602c14f744342ef0f629;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb1fc9ffa71177bc240bd7041479c581cbad3dcca6238c3d1f9637156b47b8e8000e2f3d7784b6d745f2852e038410422044b9e5b64d6cefc4f921b11fac4653dc20dccdfb7a64b6d9e7c7a55d3da127fafe67ff536591d281935f9de85a06d0493915b493f3b2276cfef61573f06ecacc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc078b5524273cda6ead8a91f018f42427531fd0fc8b29f237069e10f647ec0032ff852b6d5da17e386862e71ba71d9a1833dd39ba104993f98f7d316709742e56437af6075498b0e1ddd75c30816fa86d8d9b0eaeb0dd117025b8d41e9a93f2a8fe84856c6380eb52f64778a27180268;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d57e0cde4d601dbc188cf1dac1a1e0bd4c8d8b7ea9c6f4f00eaefad3b6dc80a901b9db261b5a25cbc6ae7ce34721dfa7d2955ede7750cb2bfb03858f1085aaee3e97eb1f52644693cc1cc8e8893d398e46986f5f2ebb3706d63ec2b3ca71ffa750b0037f97cab10e4007e0202ccbe9cf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1e73435facb57b3601569c67bf0ecdbc9c325bc613a128a2bf89b28a925e68ed8cd8c7c4af421b762d7c31c51f04f17630d43cdfb62f1128b1338e7273762e096fe064a541d429ae52aca716efe17e7a1eeb797835dd069b79a229a592e09f51736109b589e2318e4ff16c96fae18665;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf9855dd301d8007e7efd0b4bd50fd4ed033a1bf724da3f5b903dc94df23d3545261022d1b8d62dd5baf7feb05763f3f613f8f0fc3183c7bf0465db58da74bf099fe944f81c3ab024fb09d17d56e55e26f1d8d52648b9194275d3959a5fd2fa629fc65607ca41a216e7e4349e36df757d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6267c877e5650927ad4c884e5cd5f37fcb95da8f9b027d1505b1ed810317e668b684396afe43c8046272b5e51ffd39cfd20cfee960d1f4e56ed9e7e0efc8acee4a932fef9ce056e94d078d564ece9b537662ef4221f9ac97465ffe6644afe0b69e2fc3494ea06aa228b348f0a6531ba0e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45c3f96603c2f1042ed6736b090982ae575b2d9d1e132af75bf1be84c4d44a6a83f25452c767936836b92954e1d567f6ea5c971d4c7e8efb292fffc8b9ccf341368435bc52d51feb636a8955b7262ec61968349d669eccde27f2410eabbe83bf4c237553ad4b8386a75d157aa944fe9fc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he89208c4328e673e0c5acdba8868a261219ddd8184d287bbdd95e7b6d9ad20fcc90bf6e63117c60529803f9b69e93b27aeb74fb142f80ba2df88a7a6e2b497c5ade29ff884028949c63f4f6aeede98e152883415e3264f8e83b7d088a524395ec3c8c7532849a4de2d2b4629d71a51217;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c5da0fd4f0f9c4e2c254ea7b10ba8dd14da5f475061b18a21c31216f9c44b1f63dd0789f496144ecde91740ce81e57a5e57f1cab3183822e1ef30dba5ebfadc8ab49acdc58c2e27d2dbc65fc468abf9c32b5093e24630f65121a988e8be06623bdb9fb179a37c9d59e30f41d1b67780;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h850e76bad84d5c17328e38aed2165c51c8d725eb77559c6a109e49b9fc8a8ffa8b4019c409ace0e9707d294b06cb06289677bb3e0cd0d73c21e384d4005e4d9ab00da2d168e914b3446c333112bd9aade48b362d7e8e8bc45a285ab0beb1e2939a6d2aae249c7deb19c9bc736e548f308;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76740af04c6aedc2f2c9537362df2ca9010cd0587faa61f0258daea9aab41ac209a7d5d27c0ef81dd32851b81bc7af7e73b013e3fe06fc0dc873ba1397d83fd82ff5e0c204028991d6e019d1d8af3f6577325c7adbe39c824ea03e4e03dd8eb64ed3f1cf32e18334dfe9b74159f3f67ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4cd6cd6848696dccc559dd44fca5f866f40385b9968fcdd58d5fe92df9f86ca85cb19d708f3cf8a709053ee11e44330bde3b74dd0954a543dc389ff38ddc22c501e4681df7059de6e32a54a7b4bde28ab0d362ed067479ddbf89b3e430bc6cbbdbe5f0fbd818bd9cf5705d8b7ee571d73;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3864130933f265c6994aef2047a5edfaa97e5bc6ff81314266e7e627c39accb2f99e131ccce06bb50952909476a89739950afbee5402a632317c2518d3fb537f4eb1bd9292e83a3869233467c1369a7cefe875eb0aac1e66ac01b2a35c47b6189928bdd75918e30a21e57776042eea67e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc764d96488d8e0846978365c78aca9e1f3a1f545296c452cc5938007de1040ec036c7f66a76b33f530fca72250f94ed7dcb94fa7e0b6e8aec07371f8fe2586b3dab7ff1670b807c03e6dd252fce576cf38d4eccc6ad5648f6db1177dab92d704eb70e4ca8f54e3e405ef5071c90260b09;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb41ed120ddfefc6cf86a167d8770ec58dc1dd1477e3c71b185fb27c7a37946c029cef202bd0738196294d4503c52b9743e691e9f3641d93e71bbac876f09077842b6e39199753329708aa07c76a4a630b3ffa821c3728cbc8a621b390ec70d56c3ec3af9515777dd407c238ad5607421c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61fe64c1978baaeca03c31444be153424c73fee62f6aee327e031ee7022bda7a48f17ba632a4244f4d19573fde4b7f8150b7d7a708e7e831777a8b09b3c89a1142b5cf8c10938e66759f2ea935756dede3bc34ccee3f7cb7285de7d0360d9f20c686ea6b7026c9cb7fc09679fc1a87951;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a5a674df411498b048026a7e2348c3986744ffb395df96747fe6903ffed483002ac6bdae97f79fb3af21f73aa07ac163298c2e224b1bea61e31b8246e6b32ac03f99bb20c95e889b1571667b882f4393a97a3a61754764531d2d1d8595e572e696798a25e321342d93d78a73a64d7859;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfc772bd9766a97395f52940992de3719ff8d61b85e6bff0deebba63c1ddd55bb3eb6a266ad2cbc11b2e6eb7d65dfc8691cf38f2f401dc65761200ed12dec20dd973a1b12526cb280a7cf4b93ccecf154913b78ed6986be7b73092b1eb2ccb927aae2c434bcd0425f9c05111afac6325f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h152bf9efca837f7948ffb2ccbf835704619be24cd36c982bb9785aee9af229a1a826afde7c7ae919c6be884079afa2d453827d30b034d863be5287283a6d18843407af024d2371e102b7ce7cb432018102e00921fac7200b02801815629af5427218b1d752dba37e64e6274d723f74514;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd15650e087890bacc4ddf7f761909a5567741cc0465508f8aa38bb8409849d587c77e87088f1f55c4510aa065d064965bab63ac77a019180339812115ee6af397f3e4b3fbdc6f8e004cd4670eac0d1750a3dc53e867d6c0307947092a32a6cca4cfbcc808e9cc589b4c90a0ba2a7054;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf54919d5870a088e4fe2ccefb2f7d8a9389a62693e7963c34a5cf921f77656c1996f3c4e54093c1d54d14abfbb4d8750fc4f4c6185b54f4d459c4dec3d9b0f7b25f5d642bc4f5e9a0191adb8a3b4fefd68da60841a281f9f33bad833f92750cfd48930dfd2e427af5f67709acd2e9cc00;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h596cbd51e19cb8e05d77b8304d2d42c0dcd1b88e1f7fe7028b704527ad022025ec9b156f90e8772ec1bf188e36a7e75e08365752f4d96672a3b0d2a831d129bb1b0c9541e25724914237c0f1dba33863f0399b356d3ec99450ea0cf51c8ee3bb6146e1455f7649c5ae7cd2ddc735a454a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed6b0396113a5e197a5e78cd6d06c49e08adb25ed17126ee8d079b9842f0ecf803a7bf9ad58ac65a32ecb39336a51b75454cce590679e40f301c1500eb4ebff40d9f85f1fa60a63396bb796e2914a591169f0d1c1a37904603f56b7af62dac5536da7769dc9b4610176a335d5e011e87a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89301fbd3342a773401eae29c4407bd2747b1fdfd484f68b121d9be3f6ac217cc12d9443f3f446e8b538d5211bbb1fe843f4b66c02c2115c2c0f7e9312abb3131b71b5b0369adf8a5b12f13c58c32438ddc2c0135ae3dfe5def6fceb605c8baa257656dc7f282b38799d31aa7d131be02;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee1724dc627a2959094d79816f19dc0fbfa7c5c00fa8bcba2315625c695205f15a1c62c1419b0a067e928b7eec5d1b9dcfb52d7cdec762589df903c5365869a796fe95d942a225e57a9738ac1447029899391670933fdd8b532b1dda0ac5524dff12c45083766774d4ae3ffd0918749e9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h640c805131a39f6be03d1ce98f51ccb1a8fc146feae75f0cb09960811f9b11f0e93fabde6828a31592b214dd1c8706f843888efc1041139b0cfd48dd742501f0708ffe9ba753aad224721f8ab9dd8691654fd26cd7e4be1b41fffec842ec181cc71216f2b333d802b3c2865473e958bab;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd413589c077f215d30c212844212706ea69a91fdae69b5ae7a920f7c179a6f5096057f5333e6a5503572aceb554be6309b350da6e690a428ab0da5e5e5291f03131c07c79bd80d6117fbf83cee1c15779ff2777c421b2d3ac2edd10b06e216f2880ad63776cb214f6536eebdb950763c6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h63deab07ed93fb24d12358b5b8b7977f89654312f4d139c9d9a4cfc966f113942c53509a35ff84dc25c553f9a72d0e12e3032d30c0b5bb1d8e49fba9a07cac97f83fa96ae5266ca2ba5063415860966d666d5ee987eae6ea612fe6e754c27a4f3396c46e90734c19c7169ea0e3846cc9c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f762d7a172ef23b51dc5d3e88d6f91aecdb019c7f2311f20d8ba0e2622fe665b53668218b97c84f67ec5d9dba623db5bfb61f1cf943dfdcf4733ad20c8814e6d4ac3e5dd31a7dae3492e9b3ab428ca25f247cd043f961946b3f881017e7e79b55ac596966a620b4b146e886ce6cf93f7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43303d5e6eac58105fe243f95f419e79b63b87f590cd20363d6b6218e50cf465539bfc24f7bb87044080844c68d9839ad4fce27b8d61221f031ac5b3040d73de3b1f20f369fc8bdb01c737d426616ad28b5ea395ca78a5b3c1dac803eacd41c66fbc926de83924aafca1b323318dd63c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc7671b616e1a7ccf08a13240622d4b85314c40fc50805dc9b3b13c208c911ea766448142862aaf9d35ea01a8199d953aaa03942674679a5a3dea275217a8b825c9121996d1661210a35d33db5d5bb6288fda89af6aca346b15167224d719d35631ddaed5b2305b678f8b6beeeed75811;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf31add5fcbf782a8818df6ed8470d9e7f03b32651aa120ea85dd8bbea3361ed98833c355498aa05229f6f63f8468fbb10d0dfbfcf2e40c6c187fd9ed5b2d3b3fa135a9159ef67f172e64cfc826660c850bd366f2439d8820031de2b374a5a01a9b27ceaeae130aa0a5d7c7e07769ecad1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h41273adf92a71c0ba3cdc0504e9f6254beec134a9f8e0a7e075f7d9c8fa263cac0b56d765e7f56a917c17d98170ee2386a831ab8bc2d832596049c6cb2f3ebd3c2393addfcc855635de4627fb91963530e097b199ddb9cc6dca3b86dd3933d6a35c893a459ef80417be66f492b15fd61c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb8019baa92b743a0912f8edc10d5746dd498e3b13dcbd50b54bc3cbedb00a979d879071d56d5c3bf94d4bf16c60827d92bf1eeb10d0a946d7f703a4d386f786d091f66f2bbeef8342baabe6257a7b3baa55bd4d3c44e2c726f24cd4b85886e1336c25faf6341e830d7d0f68a71f91911;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90ac5886101d8c71acd2812f6e4bb9f452233c66d4b8f9c83e9519d924c9b5f15cb3b2466cc554b07a4359dd2ffbfe2c9618e05c63c5ca89e913af60d34e6c0b471cde36e1ffa7b46c0652eb70d528647048d6c6d742ed525d226f57578b8113d657f1c966ddf45e127628b326fdf6cab;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h19fbe46a15d3b9949a205e11267696c146053c1f728356e610a17912c4fc224d3c71fa5c6192bf6b378c4cdc01abfabd4b7aec580cfa08ff7fa8ff28fbc21086b463e6892775ecd9de6d40263566e7a7b8f68d88c7aca8a41a996f9e840f6a8dde2dd6a52f3ab12ff94a828a4e22f8704;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf26ebfa6908171fad87e34fef8745a19965c596fc475560081a5834f20051594b4a8dd482add9984b54c39d84848f37c07317b2236ac6575e547b76bcfdc8428dacbcfb9adeeec9b149259c4ca33e5ea6d8110e8ae25d7784839303e0c99d73acd078b4aa2f9a61609792b47030dd2464;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h124c5fb4755f8a9d594e10f52e72e3458b4790082c7038ae0ceb9cc5a7b8366a4c4ce99b348b63a1585c139fce3aee414f5a80e143255ede048e154f849a878ebaaf31104aa16e78036b6ebdb0f1bf5c6d76f1144b2c6670a59287b2bf34ea7074ce2d7c2da497411e01c5775043dc38;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4756faaaaf1b2d8d18f9ba67c975db646a59f63a8f29ce9381e7943cba279c33e36dada9a69fb929eb1d7185b826126ee2b57337564a922752f3a3992323ee26167359f5cd1ffd41989107d1c2959e673263907a11fedc175f8dfbb693ee42c595f6113fcb15097e3b58d86dc46d5d4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd739f55630ddfbdc2da8f4374805b48858f221d8aeb20626eedb2e4ddd18c77b7d423fb55f7c6ad7ba83b330aee61fd026dfeaa6b88ed1aa3a799b59bad45d758badceb97eff03d4dc0b91fc564a3023228705c3132c8fcdfaf0cbb81cd414d25a9ae4bf86e9e5c477a95c3897dea44c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56a558aa78ef2c361a37d1f4278c2e279cc68e7decfaea7d20f7efcd6936521ee95c9c694c6376d88126bdefbeba12c77a9e7dbcfed8005cabbb797b1549195fbb629d8b61832cf2c620f867a3d01ad5bc8b83fca7e02f37e6cd5e1d54458392d7c5b2e0021befd68bcae8adbfe5b012c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h742976898bee2dde46407ccbf0550dd4e48306c2f8bf7375c9c5a69a8ff3049afa1eb894ae193d9c7c3150306291d78e6380ac833013d1a63783236255f397b4f1b3eaf0ece4a646e8cc18638b702c26e2a843d507f2ffb40e7920a3f052d993d0995019dfca3341ab6da059951b081ab;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc67a660248fc984683400b4c83a4ab7427bcd8e4e36a85dc82993b9a8db4752462b0b811590c7660494b813f269d98659627e97309f1625a2f5497edaa866c7d30b0c53391bc8e0edfa0afc4ca1d0c3a8a6686fb1dbb12d26a3d651646ef9861967fc239b963defc6f71d7e2d09c7dd90;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h243149ec28935a1b11fa16458d2101e6d9c4d13b75f200adb3f4cd2111291e995e61412a91ac97572d373772ae4bb6645e67c1cc25f8cda521845a8268f44536078c45e3365978c6aaab4aea9fa259ef02c9c7c2c24684e6f8d21fedc5ab620f7cf558915a07c405b603cf58a8d1d3aa4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd9926c9c191a3701183bc107d75992e2dc7c5f1d2060f6f6bd324276728b0a444a553b5b969939fab8181b3ace75be657b5cfcbe3a1317bb5a1eb7779627971767a325fd5fd6ccb8c418a8fc560782da4d482e1538a3de9695117941c482dccf904535221f8dbb96ca06e136f5dc00b1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b441ec721cda34188b177c9c32c638e99d442d1c188a12ecc060f2a5bdd77f3be44f113998911f68b2b4e53378815a5294ec008bc5d1a22df72cead308e0d7d1562c91ae8e8cafd7747dd4563e58672ded2f1988b57c1495a89fd8ebcc228d66c41aa470eee7efd31647eee64b7accbe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e69eb99edbde4e3739e0994dae0911ab59f89b7038e5acab61cc472c415f8473f68f5f6231aa835651028cb6ead605cc2f67e798d46c2d8a97fa10eb527eb645f9eac4761f480af42fbc775e40569fccba6843e0a7d0e69b5c2723329428bd2b9875a1f98dad3984abda9496c88c49c0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40916b4893ddde2b85a431afd640301f4a6865ee276ca43c63168cc68f17c513f3e511b39953a38246d7f0913c6c5208da35127420e069956c51fb93f98d272eba2505dbad2cdf740f7dc5ebe542353aa73ed744fb3d100f42f538afdd8a56b60208fd941ca0bb5ebede03557374bfd6f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3103bdf533804e68d6496c7cb5fd98772ff93aedac7d2b8590539566e3a4e4bb36a4c27ccbbb6e9df00045487215480c610ff696e44fa9606d6e2b86be1532aa9fa934d740148276a522c2850d15d5da6fb9cd9545bf5e5642e4b6754f2b8887d8bac71bea43fa08b2c0a62929b25cd83;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5d6862a0e622f9acfc4f2cfb32079b7fdf1863a221e1c39e9f691aa1097e465a44a2b7dc233b511cfe84b924f067c496ebe91d954577577738c672c1d20bb8e3958717101d3c603bdea0778716bdb8ca8418b22fb7990f895326eba3df69092fa41419f26a43cc281943e0f9212eec9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70cd485750bad789c4469ec396f044fc9812e4c55035d1ed6109ca54d71d1ede0164fc04c63fb5f624ed6c4bc9055da7235d6e728e0cefde98e16fcee232e4597bfcc44df89fd87941b0e1a914df7340b3f2f85b28211c9ea492ec5200ee1845bfdd61cf0d821375c210c4b4cfe498d64;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb939fed6967e74af604ed88bb92be3cf0d585eb12ad776ab6a6f3907a2f661477ceda144d630544580b5aed23f320de703bdee2ebf99b04cecdbbf3aa444c5e14c0fc3b885e5edbffb4a97b4e80e896f3cbd100f80c67a3ecaef0bf2acdc2a150f89601bf56df9884c22bddc5c471372d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce334422bbd436156562ac5e4d60d745ef80b1780ce3a2f6dd7ff46f2d5491dc00a2d60dc94efb6ec63304f8aa0ac2e330c18cbfa8419b977739a8dfd410599b2be7f669a0f94e54a6c6ed08e1b32512bb9d5faea9df4de05127e89aea9238a8206f2f0e152b7d31f6033f51766e4b84a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h387fa62b650019fc2e809e833677e7436505b2e7ab5c54188c23398c5d48cdffc4b1ab418199ab9eb88c09e5f518b9c8ea4aa86df81c8f29b062df05f3870206a03884f73b3360054441bc143d812e35b5cf6e405635fa317fc663e656b4beabb11b397b7bce0a0c22c2af2b244630bc5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h393937270923cb127e6045dbb3efb20f06de121a8a3b78e2912c201357fa7a935f3f378cd07c3807af92a280943357fada68d23861b0ba58977cd24e974518c3d2ac8a01d15f46a5e955d19a30ae440a5fba4f7e607758294dafea41a32d1c04f52c6947ce3476437c8dd52030613a49c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he54acf30f2e0cd506f0b016552b29b88bf5fa7b77a0856bf2e9dafa7c6a1b9412b19ae671559c3348d51d118d01d2565b71dbd62fcc56503af6f0cdae09c7edd8ce1482d0600afc1a043564ddf0e6bd758009994067b82d44c75db5ba3ebb815916d4de081e23283041fcdb9946829286;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b434111fb1695dcbe9d95fe0a73830f7d6f252b0e28b51a84ebd8fb9544724dd1f76579f4ff7522a645b18b61aaf08c9c478b5db95515c0dedbc3c64adfdcf4d99a92d7bc683111dcdd3fcd4b4d363fbd886c5375d2c21f483bd4dc48d0bce4608f340b8584a1c86b4d2070096553f6d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha08643deca147ed35286dee88bdba1790fe03ae40dc367235ad5ed4c2a5188642e4ab75f064cf47b384943d1331e84801fde0ce944b50e69d82a857cb546ceac57e9e84181180503704245f9339445633a8702184ed73311dd0b3e091fe5c5ad4db0d4457b447eb343b2eb6c94b6dda36;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a85a09b5a32f57e9fcab320242842e34d8d58f666bf27f7fae9de90fbaeda78001680226157323bcf12b9f2c8e0d59b13b7283649a72c3e56d279bd3ac576e7016937d6d1b2e57760dc56e77b96599d3cfc58d8ed46626db9a4b40561d09038af5c0fba23d233b1ce8a3a9be9c5f3c9f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fbc009dd45ddc3e835d5e843815645dcc0692c057557c1426d7ccd426ffa5a873b053f69d044676e984fc576916a0ae1c17db940912ee9f69d6f37a87a15c75f3ca66d49284cf5267a9cdb3c8b7bdcae9e8dc21ec7b033f0fd418a2e31b7a4d6b07aa88ed71ff7d0d0033b607c921daa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4dce65cc0ebd5680fd37cf54edf88da7768243df8fd7818a711f209950f869db30157af7de2cc4dee3362a8a6db3f86a43b1a647a95ad54c7d21d3345e488b53e117237d460daaad8bf078eadd077ba9e8c465c06d9a92f703a5c5f4006e3eab2b648fc804800ee49d5effdcc293c7ff;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87fb40366dcde38c9dcece077a7cbc5b3e08d24b871207eb4af8d1dbd669b82dd155b498a16dbe5aa470f154211228251caf76f87100102573a51b7aa6bbca28910f3dd1aea2b8d08b89025be103e68ddc4c0dfc1aff9df55bd9deb75c3e97b39ed42656510570f006aaf224eaa1433a9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4ce7ba2d06c3e900f6e2fdcbbcd3b6f895266c135bd766370469263d30e40fb9edf5547ea6e66ed51797906a0c02c4e678b14f73d0cc03f44b0cff8eb6abb49b8cb24782118ff91eb92cc99e737cc1a6462f37410f510ecc19ac678fa4383d415d000154d45b75f2dbda3625733ca85;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50b65bd25f947fb95050591a1c3f480be2d2050dbf4a584f8baf3e979b65551cedc3868e1d9822ab6295f3c430ae359b48d38a833bc1ccfb78cb368c0939437a06768a0855acfe44538f6a2f1e30bf7b4d9298c22e3a91f0105741973c59ae6018b481637fa7f1ca79eb7e4d35259a732;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50ccb404969dea905b24e749f74bb7fde8f4812c8b96d9c40eb831f80b7b52e3cf794a01a65df520387e9acfcf2155f6e1bfe609ae99eeb732af0c7ee211a4e7d50a7fccbfd0241ba5e2b3022855ff5c0353bdbb4b8cbcd9e69136e0d8223b9ff886414c27a5226b77849f4447664d87d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb821d7e378916e9f9c564489bfdebadbb873e4db6fa50ebed6c436ac3a131aa15ffdaa8a70631dbfd67579b2dc907ab224e86fd37144030eff5b147857582c0dd3f0c36c11bac4513e23cd84c3b2d73bb9ac3ee15e81c9e9cb6caab062460cee33faa8552cf09e5cfd574441cffdfeb7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h33f31bdf7c8dfa23a5898a3401baa7148e09a07590e3223e291752992400b273e19b8d4beef098bebade6a5d08c4b69a459410630fb6987a0364946a54836975e9157de4268973919ed1e04358358b6fb5258e627476aa9f1c6f5064341ab7a2276561367eb120f944db37a4164e91fe5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h237f4ea56ca3f8c6b16328eb7330586afe80dc6312a249c4d67d9d65f48e1b3b2f7fec2e6ce8b5223f3213ae239889288028717dfe552f8a20f014d9afd8facabf808b1e4dcc53f56ab390b1a0833f6b4af885b2b219b038dab83e70a4feebca6e9a3177b23944e6d4a0dd9dd49273381;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1227179f5842029d3fa8b9fea13c3ed2f0a55d928bd0c44caec367ba60e785aa76a014aeaae62727c4448836dfde464670996b0d85953338c84393ccdbdac6c4a21da36bd95544b174af8f05a65e38957f988c743b76c9ed3230146e33dcececf26ede2359015824f976a5d7e63829a81;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84dbfac78e3f222fd50cb7cbdfdbeabcc0eadafe25489bdf5e5b31392c9cb4328213e59c789a7a48bc9f5c8cb01e8ab67d7b23ad08a39842b2c5aa0fd46169b51f5133aab21a7623886b894f5cca1c18be133b9873362b8c5e273d4d404c4c2bf22872b4ff0df1a7219372354197399ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3915acc4369ee78384097d71c7e5c10607c1361ccc5e683eb5f2ac5f33a31d4209eb9b0315e061c14ee3300f9434bad716e8d9ff4ad61b7afa73add033c62064085fee4bb66730a805dc72f93389fda3362a545cab79b018e465f29839dfbc5a81198ff78a002d0b1ab40993a28694852;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf62588814a0d0eb2ce2d5887723386901979ed8bb3037d24ff0aa58c78542cb79acfbbc6e00d7542a49f403042c6a4d7fd795999aff32f042ee83932c320ad5584d5f5436c04b83523c1354eae4e3a850c2ceb2e8fbb91645b091a4af97f98c82c6f823ea4f759c513345be94f198de03;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8269036e1da910f914bd6c7cbf26aa7b09694bdd18f8d231da3f7cc1298e9d724aab71cfbc741d7d58917f34ef540afc3ad3fd792b62fc4bb8cee2cc1e5eca009fa76682ee86f0a1c99c8e4740f9c70ab3dc04886a19f5294c01cc1c109ed0814fa63dc28407caf5575c3477b12ded8eb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h67d6a38b27c4e4a09541c5acbd0c3b2839fecbe770f764bcfd58ce8da908eb3d1de17eec18dd9ad3777ea0e19908f34abd3b1ef45f330300cc49979337d4efb1005292968b92adadcfb80241d0d3857b9cff87b8991568bfe77abd358bccf2867592f97a3a9c02cd2c5049b3f5de0b036;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha020e27879eb672fe0cd08ad1bc7c60f5b723e9a66dce2ba7d04394c4ad9c2ad484ee7c3610ddfdb1c0bc9d374729213f5c143a3cdf4ebe9f2a845f495c751c1328bf2d2ae0ce46419cfa745bcff8ca24f227900b5cb8cda5a6b17f74d79a32b2a10064e22ed33aca159deaa2f94d5a23;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc264116a51e9fbc7ebf035004c5d92a4ef505da266554affc52e12a2c97b74a4b676bd9a9b868e4b95a95473ba4658a0d977e377ce43f18fb4bafce58bfde17afb695c4fa210ab6f3e390ad2164dd4512181b0ca899226c52547784e7360545934cc31689b8f7768b44d5bdfba07ef560;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98466c0d5b542b4295c3c8a052178657b6a5d4683020f4234bffafa64eaa682d625508e779b9efeae0173a440161131613bb3d9fa446f9039bf86bacca8510a5ce4f7ec0458310e65711d833a1d8f0e780a223e51dec8199fbb2bfad8bb0f7f891e689124ceefcadd3ad8daa29a2afd15;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81922821c38bcddc83494695d1870b2fa324c0d3570cb1c0509b8278fe35f63c97534ac7ee9dd45af08eca7b0cf326aca2a4c48da6864d5181272b52d259699bbf13348868324f5e77fbad7de1e568611947683137e7f74f9465667c0df10ed1ac834cf2363baa101fe0536b798eae8ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ab09a00af3d93842bb17486938bd3ecfe382c5ab313be25f3328cf0c2a411b2f595304db19d65bc9aa1744ad161c348f75f9d6054afac83314533f80162a3add82cc545282d0f5341e59e7589a010eaad1700205fd88c645a14fa811b3062042466992560718cda5270105c6af9a0c1f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4058d95fcf4bceca7e0f27937cf16ff316eb0fbdcb31a1c5239068c78954df557c2ed34c42f2cf7e6d2658406ebb08fd171b08825ad071958f9e148e109329b2c0225f86bdf7c88d1729687be44f903a2145919380e3beea748092731aba9924ddaa7e9e09dfa0c202895b043fbd6ece5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce887a1aa737b95d2ffb031cf1c7f5de8fdeccf1f4841fcb493ce0f0fff0f3f493052f1084726f6e93871858bf917a2b30b2f4ee8fad3987603ca71c06741e87388d856e92fc0064ac1c4e42d125ad94b500c9dd50afd95f9f535e574e9ef07253db100c6412e293e7306faa8319c0222;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d61ed475f15e2027a4b6cb5f3c96574ade1590f45c85c7012adab469c5de6c25bb1029eda8bbe8584b1c9fd420e2c48a3bdad781af4296a837803184118aee49e12308a1db89a70c9fbba7586cf8aecef90d7cdd066ae56edfc32626a6484753b93293a541f6c6de37ef62cda1eb8a9a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h53427812e7abddebf88324b78d6e56b96aa651f5691a7265ec201e88a5eb3be10c1286257fbce510c175f7f1c696db94bbff0f1ab0eb46da0d32500b501ccf81e2ae52cb95a475298c1493c485c20a179806a40c776a5d7081c40dcdcee792ecb87d92c315838d91d66f9a9b58fafb199;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27218eb588864d5b9ba67a690882cb9a2ec7fffc5cce90342d2c2da569c466cf1dd50a53aa822768c0fc8a2c41224434b6627c96cd8a9f021f5e36d4202b4c0c90413cece4251bc78d292b5475a4c7f2d97a12e792f09c27f32e004da75af2d871be9ab14df2d53948de8ef5a82e60bd8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a3e1c376f49fe5914ba2588195f035154059831c32f918ba03b0f845b4ff6e86b7094bb633bc55bacdc2b56c919d1a931dc3b28f427c07bdfd3d7093914b2675466f372f8fdff55f00beb7f290b979c52a777c7c7750efc650b31efb39e643611063a513e13951e806a2e4ae0a081de8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c7817c8985d9f6652ecd9f3ee04abe5ba039d63bbeddf18b22436457e8e2a7885602ffd299ae66642cf512df760a911a871dbad5c267a4b27dc3afd1d7da1e6698855a1bffd7b4eb52ee93800ab8e85dc88b01e6a6faa915bdc5c8e1dc6844bb180e54d815af4ef3e0b2e07193340794;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbde0c6cf22092391699376cb1e6e4a6ac9b003bfaffe36dc7771d7f774a36bbf8d45620c07622661751fc5fb6b1ddd6952ea0552797ac1c835506a7c495a1b5ab89afa6c2c0ec2fc7d273bb8ff1805846578216dc2e4b29acfa7262ee201ae36e653f29033b4a51d04fa48c0d86a5d0f1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h193d91b7289841efd326dbefe8fecc3d2c2924af6dca2e134e4214966258b6d58ae82be63cbb0aed96f17c9e3eb4304483d9c58d5be752a71127acff17d72bf8c4cacb15c17cc0e5a1b894a7202dafb86804e4cece82afb8df4f5f02e3242a6224a292750b222255eb42067875bc4b098;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7af805f09abc8f96180fa816f01d9b8804b56ca0846a05668a8f0751df41de9baa7371ab4f451aec4a000a3e07d82a7e69e4175d331c9d247ec23daba025473ed6e448a3ff47ec7ffb78d4ff87a1e5f3e9470f4738f25c0574705d73fd161de4bd16aff261e711b20905e8e81babe684c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h391cf62a64c43d6f7e7ff9e3495c89a4dd45b6fcba4f7bfc591412ed8bc882e8b9f46011057e1e895a64cbb5097e11dd17e9276cd0a54b4315374f2233c4bd4b5bce9f4317180bad717da4b9560dcd5615a457817a87ca9fe278a1924f9964e14882afa536b285cbed6deee11b34ac96c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99799446b40af49903624e3f9ed2e9cf776da13700bc3f1339b670dca6502263722e9d01a09ae4d60a0f8bd2addbeaa882341b6742f4af6f0d4b76a014f59b36f52612ce3ee339385c597938e800cc5fd81a9704ca820e3a0b376a809247f83fbbf7ed7278f0ea06db8cf40e1a88fc2e1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc5b1fcc465696f099da692cb58b4ac3578872b3f1920f387ad008d1c832797ba626acfecc736d467f350eeaaa729f406c4c54ddaf148a96d62bec7adee76b5a4b542f84c77f84d1a39e0c14b88e6bcc41749989214a891c65b86a90c7d12f7bb4f1f3fe14d6a8dcef547cee1ad2bc9a6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef53e24488e5662fc756737fb52b43670ab9733693f02e5308f8f71a8ffdb62f3fe74d75cb8f0a7dac45422a37680ad66384bd820c6b12f3272a8526c769a47d1b997ad0d265902349acaa805a6aa31e5c0f334c504a5a7c19dcffac2d2ab6bd42f46ef867cb07a8954b52dd88af6271c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h53614f5bb658e8db03de31ed1d2a702a730d70b1a61028d172eb7127125a30cfad1782c666952d92239583a198b254740779d988bfed084386f84ff18165c574719abacd41dee38817649d65018829d2339269d2139e6d578bc47afd83382d06670b6a12fd188c7443405710f499810aa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1944df2d4c6f78a61cd9b757ba1e749b11a19f4947f4ff24802c64dcbbd28bded6b1ca1caa02b52f318f38fc19a2b5f3fa2cc79d4ef9f5bfefdedd692e0fa3dda3934cd4992ed76e36df99bbb3d51fd25744fbbe8f773fe0f9b09cdadd905aa74ad02c125800df78da5eb1df4777f614d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h20d8248aff4798f1073c147c8ec521cc2a5d891193545e513454b1913d7f8c46dd715d23711907da526988c833335b8b5dc46185d017cb0c7ceba5d695bc40ae601219caac746e320c243de75bd43a879bb3ad7f507e187170616bea0bca0a806fae3dcdfe60f59d3ef9c3ff254345b91;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fd6f2b296753e11977a4456769ac6a058836aee00fd94960337c588c7ed8126296e37795bcbc46672e991ca819408eac2222a12fcdbe2c918c983a74563657e2f293270f018e481be9d6882bc4defb8c894da6123c30b05606518d8920d51ef9a1c0c65ef5f2e56806b91200d12ee860;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28b7dacd8053bbfbc1f2210095e1f6a25acee1518031d9293f24f1ba34a851e4d2d14214bdb717f24ab2a5957fa43588a25ea44880be86fc854b4b74a45bbd5bab23c77d464ebce106a38413de88923538254ad1c170990e8d4aeba2b99443dd2b46d8b85473636f2c9027e1c1a646e22;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a2b954e692fe530842de19d9b185b5fb84ecda3177e2c3b3fa8d8fc72ede4a08362026cced9e8786deb6042eff79a9272bd51e951d27d6ceb3cc0caf6991be800cce99d3c10c2c4145c4bd8d08770251919b31bf964cab1dc585b7e02d309eb29b511872f68ed021a7052043e0c4c9e1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78391da6d1b145016b645d2644b672a084175de0fad6be045214f99320c9407811dec4a1abf9263621ddc3767c5496dac8ec0cfc8c1e09f603d2b9294ec0d5ee6c317d0fdb7c6ada589327bec402557313f954de5301bfc6c31c62cd14545d98dbf9935e22caad70a96694e46f72b2a68;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34f9008c6d2337c82273fa49ddf8d827c30db13dad7aa54521a5dfa9c842714f0a3ae8710434f4b8972d44af020afa32d15d8f2248aa147757bba4ac8617220937713dcdc3d6d77d6b8f8039c2aa203f577f032a3fcbeec5b147861ea803b1edc4dc4e17c2662b8ae0fa481b5b2744903;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c3deb9b489c86ce63fbe3a3648716f92e7b6240cfbd2b26cc38586222147afc4c1ae173fb967ab3434a85494b8b922fc0be8578273324e763eb80b82e3b1881372604f1b07aaf12c4bdfaea83c2ce1e38f359cc56fb286a3c08f8b07089349ae4079390a954ee505d481269a30d7a52d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59af232daade04d79433af9a7f4f3f065d20a6694ec7ab5ec1dd67f5381b84b268b88d2b585c2e2f26945b6d40e922cc41e70f55a2ae7214e96e92f537f37489d60c95f50e1135775206da99249a080b9357f8c19c1e105e71f57866e2a052c564746b5295e394eeb4085091e1e7a262c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4252a0e9a1bc1fab3f61da3012ad54085546c98e26e9202ff0118fbc5d7971ed57d5c7036323b3535b971b98271526047c3a46a9caafff5f2e42d2d3aa43b34aa9b82d7bafbe6550565d862c5c1ed15a79ff7737a336754859762c154a81438cb3122963410735f6c7a71155b54107f8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1202cee830614db97a0f3099ec8439ac50a851c89a142dc8056a9adb3d0ce08896693ab1e91798afe9bfc5998372cdb2481a38c4876ed460785a0c16c987045b233a6ec17f4d3bd7806e126377e1cc8077eb6393afb85a419728cb7bedda47181f46d4578fe4edcf7573be44df724ed96;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha46284f33faaef46fe20f9a5dcf813e1bfb8c3c16f249daee6015458870ca4319bdbca7f6cc299447d07ce994bc2c6398ded7db9ea1ba37527078395ff1878cad4201635d27c93d47031ed2d4ede082d02a561be7045deb03449b5c8a32ec200aa88e06a02d47c565be3ed2cb7c571dd5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf93c62208bc752bac13168149d947a609366db562fe376a5c1e0b8746374e83dde54e07117e6892c7e231af4d1db20390f7eef6694463d1b42f8ce327bb3c17e018d4d0941c07a3546afabf87e8c2939fe70bb300dfae8ccef1b00472a045397544966c0d1306b220e283cf072a5f3f10;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12eedea2db486c8678a24a9fe647b46b985b3e7d3bebe7ea7f8562cad0d2ab50afe23ea89833aa21c129bd956d0486af7afedfe789e53b08770c469206698fa473d5bdf9c356ff4a118f951151178a1421ce51d3857b5fbc98478735e04a5de68cdf7d751272638ae982c448788ef472a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb906b048fd8c0446d4e2b00218bd57ac15a4363f904a3cf2383da1af265e1c16468a392aab443e205a30fecb710f7a608d11608f71e618061275db5fadd888bb0e79eca8d066fa9d5e309546b85060f6b7a18d4cc48272945fa2b2234cef86a5674d2d156c5b8536d1e6f0acbc7164e8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he348d17f79b44e66d66249372d4c28876b06ebe58c19ecb2903ffe048c321ce6b5ee2668e50ed281edb5e5d62d7933e8a53a029a31f167d44912edc9a3e5d5c1e94fdebe241562d3e101e681076f2d2edca5116d24f2f07f59ceac3c430ccd7b97b13348bd82d99649876664b740e62f7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7b7c5b4e00a8a715f4373f7d0752d30ccddbcc7a46f9a7b1fea0da53242bce26fbe6a5364fd30abfb0c068f12299af3abb7701fe94adc633130e1ef33f2b0df350cac41d60b6881523af9e52bcefde153e8c7c5791da8d0f0124e8b48eec328b8c1b50e40290b0f9fd949a57801649a1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h133181e895956cf3df3f38441d76880181ed1f31abbcd82fede1e55445c324978228fabdd5b62ffdb6e03ff87d3dfbeb836195255a846ace0b396d3d4d384891228b21c040063171f470ce82cb6c083d89588f70a7e92954f044ad6849f8fb31fdfe26c0a83df9284afaa5a34e862cf7b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf96fb48f0fc7ad1b4d6b9b2b231ae8c4c50c3090e5d6809b6431ff95dcb43539e3d4351644bf1f49ab168ee250ae0080fe0a71dc96ca2d3bdcab33ca829a4897b53d8f8b4b4ba53454c98edc01447f4c975254e322582b4f38a9ad3bead459f37dc8f42a6c35bdce89d3361395fa6d38;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59e437e0633e93fbe7e7c247e63fd0bb2f1e61ec4631ed823c00c585486926f5530277d7506affa0d3cdeeb6b21f01897a207ff39c09b8b23eec50ecc1fd31cb8c9295fbc4de9bf78ab8c5c9408f131acf788c1749906261665482c53a649c3d986afa6e092078a006def687f2b1983cf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd031d0adf4159d1ea7844d0de222a8b492f0960088c887cb83e71b13f8ce06ca97b9b94916e1213184f213ae2dd30f8daeda79b7bf4df63a92f019e33fc9e188c3038ddc1ed489961bbe47ad82f6b7342c3334c70567db428b16644939af988e7e71b735a6c54f3e5fdf9b1713f4d98d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h302e3e0440b8189b1a11f3f8293f87745693b7a540850c37108d35965d9d40f625f759cad8fe8beb739796089929084d1b40e92b68a54eff58fabf3ffee1b787ed36d001cfa95a1543a0bfc2b7fea1482f2903a2b3bea70d7eebaf8de4875f5b32cd0c3a6252ce44c8b737054dfb4b92f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b4ee555af18d83b7a797fcb76fef539e102227a280b2145373900cfdb3d51a3f1f4bda70da306269ee3ad5c7e9e31fd12dd498771cb9cbaed5dd0af3443050061ca97f4a9abd66e9797146b30b9eca55439fd32bf90a77aab9f26cb208b491ca5c20aec5232d6d0d9ce954652a27dd2d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde39dd8a94ea870d6bc04872eec79eff2c52e158dac0c76388f79b07baed9ac6c2713fdddfe720e7762fe653867d3dbd5fb995086854212a20f403dbd121e70d8908adea33ff7074e7dcd068dffd7e37b696a2e3cd261293c70d4cd8e1f82207bfcb1686927e3c1f2fab9f50f16452867;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8920cffaef7e064119cd4b8c44b798729f41314b4a29629c49ff92ddf2b0eed0c511e882a7e63659abc622db59ac797fa48e7d1c5e8ee002b8cd971711df0efa6bf7b336b4e875445edfa373475749f15ae36261d360fc10865936101ac01f93d44db3057e3baad5baa2526131b5ecefe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdad74397a5526a814dd544aad656c068ef3237146ee445ee7d9da7c4366fbf83e61ef9cd8439637b421f49fdfaf9b78cfae4daf4add1ae4ae403caec1338714fd1a3f77447299be02bd80ec94f73e1e7144be6b52b1076eee7a8dccf9883eefa5f42c82169af3cb75d9fd8857e7e470ab;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb67eec43f61fc92cfd6459ff07d3f508e66d1a07e252ea0908d7a7c3eb9ac4d91a93862137c8f6b820f09c481604c93d59d17c34ba56bff8e2322d44192eb1b9065298e4381c96e8cbda08619178da0f84b1abdbbf81f14a37b343d81ba810b5c6430bb96272b75abb92d977c17a35e5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf30d631c9fca6edaeec7293b9801e3657e546ec4c79269a92ae31c4321bca5fe61bbf721537fab703fb58c2ecb29de51e744154d016c152bada0a76786324a9f5513f1ea67f63145c990c0e12c0d8803f24448c290122df9aeaf6c6790755616e119f17dbbfcadb1da3787d4003c7caf4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e3be0a5602a1426dbbfc2171e9be180542f912f9bf7bd97ac781f58477e65f3bf603b9665359f9a9d148ffcbffbf88404d3ac65e4e77deb59801097c5df68491c6e1bd70abc56a470ca3bf31b0cb04d8f4c88a2fd1782a9e1bbb16c1ec4afbaeb08b051e5345d5a4d31e3674c9642873;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40b5767bef81b7c53b4785c52838a1ac0270aa7b35d1f873be439841e0b79b7a3a16710c50631eb2504b321409fb22eb7e40d343c88aee6fdc649704fab439851d53d5cdaadd1829cd66f96f25bdefc10da20deaaa733af0bdbce905da208b547e7355189e453edf38bb862d4a3c81d4e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9ab64e35e4f4e244f2c4b4fb5da392e16ad6dd5f64a8113ce70552ff0ed6bd52514f8dead59354e0302e7794a8b8254b14acac9fb09c8504a698dd1c1d58017c7874f6205f3d8030e0752a099c6f13bf7edb757fcfa9093fc6aa3a12ff0c05483c17f841eec18341e4f8ad99bd1bdac2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h142d09523f5fa764109ae3b89ca4da380d7fc150e7f4d2c77ae0a16c4bd4ea72885ff87af5f12d224e90ab774ae15e3057b8c6f66cc169c5e3c96e67c4b5ed5ef887da7d4b37c6f4239ed1e1e703df3d33cf7803b211125b3fe13ade6acf92dcba373710f2cb3032230008eacd11c3218;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc08c100870405a07134c77efbdf6b9c5361d63cda8088695459bef396fcb0af721b097539cb893a05dcc892d0049541f3a7df29c49e6ce35b11dfd8236b75b7b624cc634d31ccdc23b51bd2b492e0d8e61406ed367ecc7739500e32897bd2a2da298d6a952ea63b7ad3113560b225c324;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7b852930c279f864df6a9a9f5d409b4edd3f460d7f920c79be306956c52b80a8d8928ef3f4df631adcc5abf734cc03e295d684d1503358ed5cde2e4147607e9abdc70f9714274051c71faa8fff8cf63cd17d4b7d3b5b674e61c70ddd8f1ab0bd19f184124072e85f604c25ec06f2a2ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he64af6c1473a4b0d75d59ee6e1b64e7a5694ed51c3334a76c37ddacf96ab5c1f03859583204032bfad1a147d0a0556b480f644493c6a5327b0222533ee6e5988d835714b743bb0365e902bcf2d2601014ab392a1c00b5124a429ae2d152279c0de203795fb70918aa055fc1b84cf0a948;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8a8899e3efea7c1cda4ad26eae0d71931407f886d3991ab8bb94f2ab1a46842844b2b0e35e218054f4257523f4375a187c7d1d03e4d1715e3dc5e954865ef84b5ba61de6762cb025fb50deaa4891807cdfca9720609bd870aaf8d1478034bac6edbf0aae9547675a1e7066cc15eaed4c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ec21723f4ef425d1de3a38876ba1f70eeb4fb162a1cc756bbbe4756f9f396ee458fc795a276fc98b3128117127eebed20437e7d88713210b9549f98e92997ef79d3a37cf12d444faf69eb7e8b015070feae16a777bd45ea36cffa224e2513236cdf8901aede1fe5fb3a846ab787b61f8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99739ff77b4f52b9bcbaefa5efee9fa0da06f0c115010e65d8d7d12bbb21d9475d89540b1ba1cd88538fcee785d3f47c2dec91ab2ecdeafb21e72fbb07a549da268c968461265cf55f436d6f3ae1039c7a67ff5af3111d2714ad5889be8eaf0e2577da8841b76d3a2206540bef77c816c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hafb26d5214dee6cccd2e35e58f7a5e34bb05e96ef8bccc6c3ea26b73f4ebc2c2898684aa910e852fdc06f04640e98a1bc425413cca0b98d6191ad56ee0abafb39d5d770e4ee3d314ad017e77613e9db0f6f693b21a78358430b6104ccfa24ffedf232f9200b7af9a2af666acad4d5dafb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9015d50d42ba14fc7adfecd531e19e2bc3551e1ed69a7e00c63238b801456577f3e428baab73c6eb24c7ee4a54b8a894c119bdb96546734f7d7fa3e69c3e59f8f0d80ef60a8d6e045d099dcae166fca9ed5427cf88f3b21a47ab1c8632386f48b0447b492e8f9e291f7637717034b13b2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf5e1d8d4a7011b074dd57b68900d38aaff7b863f3dcb5a16d5a4c21516e4eb880beb7be3af27f5a1c6ec4454d6562ecc0124c04e6062128ef28341738466ea80e7a11c2b17642f9f5e9e13b795aef24493bd021b1628a446ae150ae3718c608f26c2841b3284bfc5306a99f3d4ae6244e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49200bda5379d2e7513a90261c16e770e1204b6c6b90c1d9720ce736a66228278c3103a5f155042bd13c49cbd3606965b7fcb649d1de445130d20dcc4e740f835867eca16682be5f42fb71ff56e01e4b29de0a36f643bbad7771b95bcf18297d2b0aed228459b4fe57fd4292061e0375b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14cc1774000e4760d2596f6009670267209f311edea59a89487907375e99990751e61ea630243e6beb797f3da3d4ebf3d9033237857cff527f6633ea4049839344a678483f302119b68a0784908bde1994d89f09ae76b177ec6048ec9538860885514895f0fe460fb1973171e5fc3f8ed;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf754bd6f99c8b99b02c5dc2781adbf94426162bad7124697ed45efaf482c82510510e902358843867aa2fa0cd44e1242b5840e7d184fca20211619d06cf8921ee8ce69d2dae391acd6e598063592a84fe23329ea489db71c448436dd9a1dc9de8917aa68a61387dfc9d345438c0292d3a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h425885c08ceb6e33b478a261ac61a792ea6e86345d23af4412343710eca438f4a14fcecf91c6f5fb0701e03f767ea462a5e2c3874e31529d08a02d6a535c71a73791bbe03e03145640c6ecb79eb309526fda1a862540b8781afdd08a19c8027233f9a4a3cc6cb3ffdc7e2df5a2eac6dd7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf73505fa05db478a0c73c632f4492f8b8d18dc44f5dd78e1ca30367bcdb81d089b67007cd1ec1cd6fd54edb7c3457fd1fe8f4a4adf651243512505e3be42dae30abdeeac46a41dbad11769d4e354e92842692badc2489fcf7b06efd6ca7ab18476900951f25286f3f56ecbef4af151472;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44288f11ae673e61fa89ee830fa72206e138085b4d54e551df766e15b13e039e7a96908879009b93fddc008dc3c351b8fcd7cfa8bd049d01ac62c60e831f288b300b565718e19af7353f0e03652da0d8fe2012cc3e516d530969f6f77d1dfa814fde71eecd79da0956c41a78c32fb4f41;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ed31d0562deacff3a7fdfd46ea09f1d210ec78196b069219d365a0f52e3136b3a679eee75f9f80530806ef27a0c66ddf2fd80c762991b5065a78bc87e008ddde14baaa37e85beab2b859c98edc153f1d790652a95580e6fdeabac91bc71b169a4e1704a9d3bbbefda35b407d09b45f72;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb1667ebc94de381ee74f696b76ba72705d45142b3f851ea71c9dd5f15016f6ac5a33afdcdc025a665591515e4673b3ccf6ce39935141bc9fc72e5004dfb696044b28c2f5e3801a22d9bb4dadad0181ac40d2620c7059999721e491f924e296f0f5fde9d92a2838ed3d0a4ef552a88c9b1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14c07e0fb779d67477ebfef96328da96676d30ef6b0eccab4f56960aeacfb69b41fd6cdf574c9fa2520c43392c79e948c47cec410528bcb1f87fd437ab91fb1b4010501e701b9a1dcc2b650a42b27c5b064bba802d899b61b7f23ab65aedaff3333b9b92762ba748730d27ffc39ba2c4c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdace71c64753d9778f124a4c73cbf71f30e5a9497d16bd38ac0f9b95c38b3c9c5ef382025e0c34b7d363d13dfc64968f2fa3cc71cb14a96ba2ad1309663a42f5b5203b036514ec139bb750806d4ef2591029658616421ef8a1ea110f7f78cf89d9ce8d684a0de0025c2cf02b40b8140a6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b943ec4d164afe0c52d17ce8389188d4742bd8c514fa6c994f1be28e022932c5a7ac9f2f9c5931b0389297904b36e49f01bf63fe1f3af1dfadac71671fec90e0122c671e943885d13f6cdccee7d05a990cf746d196266824d707cc3ec5f87016035f0eef69d946b8ef6bb3e794da27c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd69dbf3c92b3bb5373a8b168453089ca3177c12c5c5ba7f8d3f8e78c15e1add5b42d9a81750657f9ae7b34561c7e86eb640b532d03a701a179e7c053e2107af56f22c9e84a7f1cf398466b55b40524bc6207cff7ec946fa12e0686be14efea12d221f65b0326834512601c4c746ecf324;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab9f5d1c337283b30e14006690438347818995dfa9ff0e3d2a81dc798b9baee7da160b7a0a837f8106c59bece2df816e0eb788df882e235e9eced203d918f2ead248a335268dd2dd4d2bc39d89f3631775e13923abada462a36da94d2752a6c76cc487b185bf4f2444aac94730c722666;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2572aaec5d19cb4b50c7f4553ad688b0713bb458c10d8ac525d3464679a29c0aa3cf92cadcc4bab29ac872cfeea92b8e380d4b1a4e9d93215fa85ef8826f473fdc21b41928b270289f3dca684eb750935977e8bc46053c550f3d8a3da63dee6c09d90754afe5cf3441c304c891096c7da;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h934150b39bd667204396329a2fa04c9670b673e8939b9f49c64b6d2e4689f397da3027d3e50e82bd0ae834a0f7398e649e951edae696010a5bd151af748ff0c4e9bbba3855d7a4138dfb1bebb7311c3ebe8331c5c4c7b8e1d493682078bc7963c6028798e767af194be4496c15c92b2b7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf37741a32da44a79fa42bbbf34f85737b797f7c9cb27a1ef6ad0473d27fc7c2237e1d018f61a48e6ff128b3716b1548dd858fe75e4d4a47eeee1582551b5406a82efa1f12be51148dd8211b4696b8070e72b899325a05f9435013c916aabd3765890dd0bf2d59e7127af12f12c3ac3d89;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9dd41339df8cced4275e3d8c854d3c15018488c96c0d0da519173f5a18484bf338951395a76b1c9d9f97540d3f8b3e43b9ef6b1834afb619b257e0142071ead9bace3bb2e3d75d963f7b81b8f36e7e1644379ade95d86bebad827a76400a692a579f595404d3860720ffd16c37932aa1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha397b4b4d1e8f99bda847df980c972b68523dd1f6e74a98f6e579bc30382ee7edd8ba8308bfc7bf054e2f8980a33280d538bb19206b8b3e23d7e97f50411365aef29b2663ec3218288a7e26a8b786c47780302beb99ca4b40f04f6377b176660432b09bd1d7cfe810129f574295362517;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf3755a648f240217048baf2d3255809a211377a4a476a40a81b92eff9d63fdcc0bb26a52174f49ea2a3ca66b14a716c520ba11e3b2cb2d57cc73df6d705a9c936c2ee79fbbf703c1f61a6035a0fe2c75c61396782083aa892d9057e1aed08463466263609b5e080b6623fa84003cd2eb8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11802eeb6eb4d6f47021cea181137e25a9ab23562a4ef6b91ad6da42123fea688d64561913b7faab2b5f8dd80c127891332906de34b8047a71342341c81f766d3abfed7e63aba5911051ab34acdf09f0689b5d6fe7d149061b561b847b32f50e2fe83bedecafc14bc29f89a34343514bc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had11b713c5891d75bd5ea3bdb018048554462d13d2fef14e129021ed2af890929bf35fb1c0a10d20a2716533cbf3ee467100b35bea17c71cb6fe512622b2e68a037b9db5e4638dba710fc869ced2665a8d28f9fc304ab8b015ff0bcfc73080846db7b59cc78bb53bd3a49473bdb83a678;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd328a34f96ea32ad768d0296cbb88274defd4027dcb5e0faf888b8fd619318602b3817e6b7eda7ea84c0438e78525e02c3b9eaae2a9f7fbf0074031419e347a0bdd71397fb8df8b34ee68cebd49a9edee43e29ca455f66b822f2a4245b5b6c4a6ca917f47b33e5bdfc8996c3b2be8654;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1cacfc849e2a78c7d94e5033ef30cfb8645edb12bc883ac0da333556d481ccd87c787d637e0252786d756ef23aad4ff76199d74b9ed748087542f8b4357015e4a2b9a29379a76869ba7416a5df850fba9b084fae6fb8ec56fb6f9a30d0a97b2f702fb4f1e3b4e7dc62086f8f4c7c49b7d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24d5c7fba5de043d397b134da832cdcf2500491043231e2d768de351a2de4d99f11e13e67d233498c9e89f502b76652506762e5fba931c4cbbec00c783ae0dfe283f3936b2da1370ba76b81c778a1cd96c5e5af6f27274e0c5a8e5ba36be158ecffbd3d064a49574665c5dc0cdcb047fc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h752c29da24205687996be06c649a84883e9d70e5d3f88b31b7c307576a3afeb4cc566da9462275aed341291bf380f674c9a8b31a0925467bc1b6997a1980f7b13285e75ea023300e81608061c81a2b4e205c9fa71c16def8f33a3c17606e5fe96a356f3d77814bdf248dc9953e68574d6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85a0a84c55c05c97215dbfb299735f3b035928019b9b10db84f3533c409903b5146ec5e01b14f1f7f8309252ce86cde6a18a1b4ce6db810cd608dd5e18562a5cea89ff0d491783b0f9f91a15338356bc2b0c639c052ed3b44b3269850ba804edbce4a8610077bbe0361ce42c86acf6bc2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7ac36a90506c0f94607187ee5e7785587bf20a7a38ca3026ef651cd0e2769e16753e85b8691b4540608143ca8cc0d03fb34ab8a860ce4e2e952925ee3745d45de2097d2c958947e0286eaca3551ace6c5fb08633235ed986b3c734906c2f471423b936b6139161e22b8405f983336e17;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae94fb663e3248e8b663f862d577d21366f3e4eb91513d471084e3d81c76321a5afb723a3385ed355e3598c5a89e22ed774b6003baa185c3ed192fb0e3fb72864459676c3a5d117735e58bd982772016e2ffd24598f41422428235c185405f299ef83345903c3060f6429db214d8c465;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42d46f935ea0613a1481a56e7da251de11b88729dbbc208a0d0669e3b7587d78ce8e9694c961936d7e0954b4112f018509eef78b1c34a1f1c89d896bc3a4696d37764aacc14859202272a57ccdb14fecbe689471b15615461d88db79d788a6d3d89d9f916a9d21b7907a9f33ddc7d7b15;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ad0844f8b539f0456aefba76d05373fe296eb4efc34140ca7fa0f34d4901b04fa7c935058d9afb03f5904cb299b7e9da11f6b5afeab0fd8afba1686d35dcc817fe8c99262845b8d5bbbd6e44535628805e98c363c18ed4a3fba4813f80ad5cfc8cac5cd78e709d60ba8fac13e03d61bb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4897050299003aa663cae8146de57e697939d2c9e72932fcd7dc2e2aca079a2f8723f1214de91f62291f3859d30cacd857b8743c4cc8ecffc7e982fbd47ce1130c95cbdcf144c714e3b44a562ebba174d279acde67bba9308cd78e94ab456e7c835f301024da21c175f96f00d588b2679;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb9c2e98c125e92aac0ad55870e70068364c4d94b88a59f84ff69dd967b0f5395784681e6f28b4c03b04b9313a6bbb84b8e8ed57591080661cb52df5fe979c1bc2025d1c31983c1cb61fbe30e495386b37dbeb8c49e273e1eca86c8e45e63f82e8fbe5420c64ed6c2382740aee027a5aa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7408a73a3c11847f0b71959ec66d7a20ebc01cdba559c06854ac80e7f6b4f6147cdad05e0d6d4dd24009138fb3de94ecdbb4893f1991794c9b20cdfae47f73a0c2f563f5ed3474cf3c1bb553b15ab03ad37c60dde14ed0171ed8049f7d7f527e3474d5d7c54de9afdfc3880fa62d8ae7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h419451d3c161ae837e6e6d97f2b430b8ef18112656a222832c9402dcd74cc251c43a5e22775d91e2a513afe54f7b0ed55f168e5c9d8396b8f3088c9322c5e4d141d691c1def76abd1e3cde17ba69a80ccded2a1f031e11c897fde70cf0e5fcabf8e15367386a93fe746f53ebb1de71cb4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h783378e0b474813104204aae3906b75bd459edbdbe27cc8883f0cc19afe06a5e07932e02652a1b61feeb779722993483d155f9facf9f3ffe6b3064811b7cca0aa3d4a5b88b1b87c74568d3337ad48d6cade7764d28d866ff49421338e31a4ac4763ca4c72002b9ac66b74463013a2a5c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haed225c8dd994c9901e988e3c878100013f220b0004dd90af3a63006cb7c2a68b792eb06449f581c302457f955a1f77cb0629741f7cff2b2602dddff7cac9d7a7b7ee4e41f01a534b9b28fe4c028df2f2cafc6b1bd196689fe066493c7a2f737116f34278846f63c6628fb7f38fabc4e9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6c2297f8f44356654757ad1d8509261dbab299846511f74479e09167aa6c78492b00a8da6959972be68637e3b55e4ee38ade36188c482011b6dfc3e9b7263a9305b5aeb4912709775e77ec3379256a5937cdf9caabfaf55de83fa8a59e7b14bfb67f3af74245b7aef87790b9d550be83;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e461ac73e8df9f5919504f8715cb8b1e1607433645a929100462e7ece731dd4eaf9706fa41aefa5dfec7ceb56706941cf00f1c6afd648160f5ed1557b1dcc3029dffb6df63ca9daf92dbe61b45784e70a3b694172c5f3ac05e673659b802968035f1f53b981d5b767e9c1d4ab6b70e91;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfac388c44e6de33d5c42bc5ff1da1768ff58f2ed586a42c1f773e0f8ce99e027bd425d9e991f12fb0fe0e2bced34725d8bff915760fad9b8f7662a3740d2b1b17d34a199927d01a5122da31c47dd5ebf6492bed55bc4cbf6df77ed45e03e75c8d3d4cc648d2d6b8643c9f4b9adab0c47d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf98d2c3a4a3e440752c0c7edba36750ef49ee482e521293ef928125ad6e85dd39b526b55625e95081958fa4e1fd59a32f8d2602899430abfeca1636f10d395e66041674f8203f98a1efd3e0f47d93b597e99e7f1998e6aed08be2e0d900e43a48532873cc62e1153b2cc45592dd84728e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h19a8b0d4a5bb45ea95dddcd7c60c283871a2a61cb8c0ad76e853ae5c1db720d0cad1d8daf8ac8a0037a54400b21f4304b70da957d4e4b4d6534a7166f9abd2e04ac2d139f088ec0199ce4461e52d424be095e286e85d18cf07975680f52753f5cd2359e7db82ac00e4ffc578be52b93a0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b3f197a665c3f719be6aa80e05604d0338db265fbd7e70f7a1f272d27eb5c53c1ff2af68acd43f2500455460f2a31dc7df26f4535131ae1c7e5944017e683205d95d5d5b2429758043ba13f57dc86dad4732730e670b8bd48670f6fa55ae5625858a0dd7728b5b025b4d2dd7b474304b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had3ab65f6d0848077ab68acb8b53fb7b1f6a6753eb696be34eec085cb1833539da223ea86fe66363c228f5afe82e1c1a4874ebe8b55d16b33dc68ad08387afb601e7381bb23eb56e50f28c0bb73358c9d539acf2ee90e7544043aade9c4b5a544f0ee371fb350cdd7fc78f69b532ff2d9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d9c8a9b22c8eb10c4ee9c48c85c4f54224504c512a36faf130a7f983b23fbd58e7dd21c4552d1d64794b9a4876080bf6a0b0920fa31a4c907433bec930469905768f159850299624287cfa7afd566fdf051f4d89d5adb6a7a6d186eeb2278f2809a02b89fd4cefa7ee325136a91f02cc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc7a4592e9adc5c6b4468c7cfdfaae080e47db0c7951e2289468bbfdc9c04704b8371e0e6d6f7bed1f50f2b1651dceb818f5b42df6907660a4a7a460e89920938b34793f062c33ad91f13b0ad746b450f52a6e54017dd3247e6e4d263970dea239776bd7638937edb91d49f21fa8a66040;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca4ac555ef97b4500f76fdbea29458b1eb45212753f6821e5ffd3b0082c6fc4b9b53ade37ff5c3bda7aa1b1cbfdd26040c5f21f13e2b2acf266cace315105a6d31f7f175180d17356d162ba525b11050d443b615a9bf51e9d57981c1cd54e84b448d5bc71be94f9c856d1c7874119169d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb001baf9ba2b2635feaeeb63784d4b337db34e0d3625e29d874e43d90947a322a967843b87039887e9b6af01739f1cc3100c7a8923ccdad6cedac73fb0af1cd476a30b477c5ca002a4319ffbe0d6450a5c084eb0b062c50cfa6b8cb1be449237f592096bf8a31b623290a205ed136829;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2053409415935fba10d293af4f963f897f7bf66853f516491eaf7caf6b6afcf04a6f35025140eb4a17f684623c235bbcfc88468d1c29ddbc6fd9f9a880524751cc12d1e3ce65b6212c6d71c26bd2e3e5acdb204451be8095e033ef85e6d662d8ca6f65a3d3652ab1bdeb484562032c9f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8646fc78eb63bcdb0b7cac4b2d8c89009d6cdbe158a0ba1e20159a104ac6e956ceb0cde51d0fe7801e90cc12e45f7b546a7d4a7fdc1dc04c36c8dff87a2ae196b5a6e173a6806e8c9c9572c506d1f5bac9c9f8e8849a363b9633bc8ec7fb5734c8938a7ff8e2532d840bd238146ed7c0b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66c38b9c386806b8ca07bfb50b3dfbdd2f1a13a3766ae05286350f8a8d9b2f8c0d2a5c5ff521d6609686d42dad6bccf510164fadfa080d8bc4bbc8bc93f7796c8a5f7c9fbf937eaea461501fad0b646a66f8e4260d7b834bdb4e5652baf63b6e99ab0b2eead5e1e2e57d32253b8c10d6c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h555d7e82729c24e216f9787952311db05c1f46b161ffcdd60558cc1396812303af39abd8a79d113ef710c65b011cbb570812cc32ae8cd897f7b5a52c5b5e1306e87cb20b8b22c72cd30fc4657283c73178d00c426c9c36c844596458fa97e571a9bae98f02a7e16002d66f5de159071a3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h930a78b19f0a9a00e17781853644ddfa580fd4a238297bbe9a063c49ee1bf2c41988cb257e4b6c1b296d4f95344a26b02fe6c76100e62133038df39ffa7bd7a9b5345731848ce5fd29d3617c21be468376bcac160b951dd3c9c9c6517aa2950a09b95adabd90326ddbab779d3a88f2895;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9fad3b6c446433c3e2c41f5ffac8252db89add8127f3644e61b66985d111b1b83e6094fdde1a74e11415bc286442aefef8c1f3129b4d0874996d09b761192b15159ea0cefd07fd615b32edc4c4ebe1c20aac3d09324bb8a2f0ba76aef7a1430c7ad41c18a3d5489501d051789cce59a07;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf5409038a6a24c3059f1c74d08c59362fdb406576f92480805af9f3d31da714a55d1386839499b47c1bd1f67a4ad55364480421e89a3bab9af118782d370ddb19e096bd9cd277b2897ee1fa9c1bc42ed8ac1503884326b7668642956b7e6c4b59b196836b3f105c01b4fd7d9f49476b9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a6fcde2d6d29f5a330a6187dbc3d044ec97aed1d1b9ee99d3f8d1bd979fa2ade6008b3cdac0df662ad21fe59d909e4fb5c7e0f16011c26f53bc83808017671f2009d5fb97738cb84d071db5f3dea8c2946a22b6148894e8257267a56436b3a632d06aaa95935bc3acd30e4543a91a412;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5009345e4b584a47656d35c508deba56ff1c3bde00d18562be655a1a4c871f06a08a863da2bfd62fee54a8d865aba85a0ddea5f821d04998b661abdaf44bfac7cece19272677100eb8d79507c69a7cb9b2636575842a1ee9a89966cb01c86e8b5a419e3fc5d915659112877fd977023;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f41ae134c6105cdad3c89dff3a471c209a31da2398e4a9cc7dcd14b079286668014345cba26edb170ffa014b43c0a90cde403a63ed76eee5639967249447938ede580f1785e1c1cdd31f9078ff6a5bb511df1c83069dc97ba9cc4d552e4aff3aed9fcaa613a8e9efe2ecb4301d729f66;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc54b4e023b2b279b47a571a4890e4afeb84eb1f9128fce780f6871b4d5dc2cdf85f9fe4be0a53fee93eaa08148670e2c5c7ef415359d35b3a62b298c742f103759ed25fe729a32e3881fdf85c1b730d69b6cd5acd2366e04145e018c94426396d0ba5c62d45c7d770972ee21a0a92ea9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a04ddc0561cfcef5aa093423a7139a41cbcabaa63cf0e11bf87ac2162028811f587f6c2d87cbdac058e0ab54339db3fcbcae6f62c31e488f0e0033677bfb36844286e4f307132e0e64f603455bb2b29ed203efaed5216d6e572b4539caf364eec462a9ffbe3181982a9ae34a34ad2bad;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc3b2af975a429d1c645521fdec7d73772dc3dd0a6ec92a410909324c1fa5bb6b01ac8ffceb29d22a66f24747a2d69175e8128d4670a3637855e05a37c7e41d8bbec7bb83f09bb040257020ea3e351172a8042cfa77e83e16554d072a8240ca77680b4bc694e3f8c15d4c3fb362d1d045;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fd5960a783010c9a8ee2505880e6df378f6378206da63caead0b73661a9e239c9f3468cd0a9a9f552e6f3c08c15b2e07505f753f57e3849c44dd727bb9fdd335985960527bf533da6d40c2cac312638522d1fb06cc8c7f06ed495ace7cd9a8658442c8ecfe07588fbb303615374dd4aa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he284f49e3e984ab00d4025d4c79c9e22736fb07b9dbb0a784faf65515794debd812e00eb8a908db3859696c8caeb4a48aa84032099ffb6365e271d142e8cc6e8d2590019a89775ffbac1ff695cd62fa8115bcffd5f26238dd64a1a5a2a298167c51e34fa6f48f1219e998e5b175f3dfb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd151889b1bfc0d8ee13365cf9cb1f6aef2f299df8e1bc74baa6fe7e33e35274c1b12f493b581aa0a0b4f75da0342db00b3c2b45b7b881d82516a4f29128effee9f8bb9186afe89bc9cb3bf43ee6cff6c09b4d622e4e75f90232c24d00b11c1c47a4b3f5de0a6bb111397260f89a6ce85b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h136ef5eefa2ecad26946235cb2b1df772796fb98dd76bee2909b6d0622bda4650ae788e41695ecdf39d917515d91ac41dd49799650e3f52a430741323c4d9f291d2969f256d315b881888ffd00bfedd5183437cc0a01f6778d02733cf1b946e08fa30e113c508c18bb89e698e0551b3a1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1a9623d0f9a4414ddc9db0966ef4e9f8f426da37a6a7889e71d49b24ceab2a5b8068d96ca352b73142f0cb77c8cf4a287c95e6a2002510f5aa94014740ea0ec03321638ca162c821419cb2262512db67bb7ac95f42de6f63670443add37968fd9a155dc289cf009e6d795cabbed87da6a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9828cc2f511bb31d0f15864b953ef0ccf7458213f408de975b5fcb004ea2e9a5f396706da1c7432a1c337e066e342a6918038c4da8139f8358b86f897091cbb5e8c81d857a450844de0e11418b124a3800e7b4b6aa4fe12525ce53b7daa2628de364f9ac46010d1621277ab97435f5b00;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf7183c5a0c3fcf40a9c163eb558e12a742e22519953c55a9dd8add85f540a1ef1bf893057edec29524991e0955aca0f14720690a6ce08b8b09a5b53fb866814ca680aab74ec0720770985cda4a3c63ba3ba0900d652112f84f671f461df88f2a4f4fee391b6ca32284a85a56614c97aa0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc282b33c5448e1581abe61d3a87dccde11a8348e82f648cd9050f926e597f9f05483fe57da38cec8536ebe9cf5009544cd56e3fcb29702fb1516798d10f4c070c03eaf637da9a0b3ffc84576750e1ea2967639d2904ded5331a797f056c3f9ccfe3506a53f5b55b43c0392691d00b59cf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbce6327e113a4c736206fb4c1486653340cb129b293807441562a387b97167623d9fc275f1416da57884bbdc029ae0dc97eb97983eefb54ef0ed5eb13df1eaa6d9b0e1feefbfe1ee754e3d4043891a41c023832cf89e6f7743614f7fc0dbd9375eace7a0bdf32f45e94de4d2cc5632ad3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1db2feed82ced6dac89b9b96e8ccd96d37ce24dec994a2479efdf686fac5ea6feec2db656332bfdab3da62176375fad376e1acd37dd3208834252afb20810e1d2d0675bd70db79684fa155aca680ce2816483b149454473a1b5d07eec6ee7e0db45b252d5a3f453b42d90c9a00a0425e4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1418941680908f5cd013cfede7f0f5657a3a528361a14c4f1b76cb148fabcc0c5ecb64d06f629a2db67708e5ac6525a4ee703b28d92a2bcdebcf8d252ad9f25946598aa2ee444f1d832327d66c2a6573b0857a3cb05611c9dce79417ae566952fec990dc2250f06ce4c69003e91fd09b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7034f307b7dfb47af4fb91503a15927e8b7eb1b1191bcf60f8102c2edb74f3bd19e075c18b51142c431da09c30d278e638bc0ea387cc414471715bcc6d6fa95533b5d45710b89200015b04bfe51a26cd7ca66372cf3b919e6c10e73a9d116beb2204757099cdae7184de73a4013e52a36;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha924736ad7ac60b6877db024976d635ab4152eee14dd6bd3219cfe32de092449aa6c7dd753c4b482697d49c4bd0f251e8b8746bd4e5d205146fce6c14ee2238f6725416536645188ace15085c26184f8e0aed4da1261306cb5cc9aa09402205eeea509e55709fbc53219f57d65f5e9b9c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ab8f4f08e4eebd13e98258f2114f66025344ae3aaa24ce75e4420fe12f2e7a2218bb39e4a9eda4ca0b139612cdb757d930594985513f8d8d620315fb653105de788889aaf4b665df74b3da652d63385736b78aca93f066e19cb6bca46cbf0b74f6a06a36f0c18e22e64db88c1b0eb9a2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb3f940ebed8e39aba31cbe917a91bfaec29f34242f1571e1e1e586a85416d65e72c6b700fbe86ed47433ba8f1a2315b76f73d90655822a7a354278801d5c19ef843ceac1522eecae4e240fa6a7e5e46798ff00b09986294989126a96814578d72778054e6b0f11af05485c625002ecfd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d5eaa6bfd788f69873301451d51f38d91df69c9a3d05521039787c2d6c1c6c18225b53f2c18976be930bc132c77b1a6973cb252054ff74ca7adf2f44ebb32737c00f42b187447771b75555283859d5784af76499e1fc06469ed0957b0453e8bf9d15244993b6ee2200ec94949598928d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99978d7105c92dcedd14414b09c0487f8246a88364b5214edb47d2bdcae3285c1a5a48b72c82b0f3082392b941d5612415271fa21d8483a5260f66ba491d6b61a10bd9b67a64952757fde30fadc6101a1c4ac5a10f829f25e6a877a42d2b551f67f81313fdaf8199b1c5ee4d628f29382;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h86429f6326493435ab7d5d9c504d0933a89ee04b530db4e71e008b46f5046b2c7065b92cae65ed371963edd1a4a4853b18f7cf4d01df5c032cdd87a8d50e6594e24ffd8a124dd8c8c01dbf9e6730e8de1fd40647d63192e1ddaba3af71f0d1911c3f48a5b314f47ec81c61d6dc0cbea8c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1885d88b4ddddde6f3ef8c7e0c9a7f30ea4dbe528260bb90498e19401c2914515a66b00cbe7cf80cf24310a675e71f548a10f1ad46af5f4dbd633f8adb0236fa6371847026fa7e0ccc34a32e97f465af0806313ec0d7b364c11789e592b20a082f80b1baac0564b43a8d44f2a3dba1f9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8151e5a436c948f620059f4df80ea5e1e6a1d6b109928374416388b80fbd01cd4e171800c117084a60dc0c6c79cb817bf86a10987a791875922d573b03f32615040df86c21049fde10c47d3a1a9863a7fdfff5afa01b1b641fc2b5930619e91c13f83bad6c9e4329812412220640e10a4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7489a466de499f1a3c794da9d72f8f5f84d2d6f031aef12561d601834431753c5ae25164df7f3eabc5db66b9e17f5ebaf523bcb58373a14a9fb6101f16df709c01402905c257c1755df35e13d2c12e4c75f8de3fb0c008cb2cb2c9120575ace6c9a49b9e8860d74b0306cc8484aa15a00;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hccb2f9fac94890a5a52ef008e3893a2893a4cdc9491624b311f565e1aa41f01f6d094d871b2d2cddde41acd1598540df1da9bede407c66a2e3e2a95d0ff3fa244389014eac442d9dd288f94a76eaeade43fe6db12a451a20f7d1d010315d3e9a8550af294f8262e713878302296b76fb4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b38cd8c28d9eb15fbb00547ce8fbd4dd4a0041d9131d63c32dfe2f2ae0024a11735267f357f3eacce9e7d893f0e5c0a9bc0ee738b5baa963a3145d714e867d8deb4ae2decf59be5b0b7810fed14c541db71a07b8b474c95e07f19f3edb8ebd7111aafc50a67900115c907c2cbf11837a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2f7d815b77cd61e115a8d58246838fe75544c141446a29fcadca5d1fd4877ffd7c65b66393e85e4875aff2508785d5cd274483d5fd2fde9459c790aff5900e7c2b24cb1907805ae839d848e133740a1d7286ae481578936668c0bdb3de36da3d1c277c5b2175e06b3e4844c24401de07;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ab837a4c62f254fbb3bef37917c1aba4561cf6314c8e646c80b90ba6f846230e5a7d98cd6b52c0a69158a7d2668acbf4c9f947afe4efa7533e17d45852a9d80df6b66bd7ecce7ed3ff7619ac99eb4faf3a196d0b5b1afb8c158445a3471febf29bb81eed5f52791f97eef115a85908d0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f3e6e04a7e1688ba1e45fa93548fc2107c676730401df304e53e3097c861a549c4e79029d1e687e60a2874c0d7183b6502c689661a252292b5b67fce852b840eb3048cc08199393ba7625388811cc807b7b803cf6e15732d7eece4a968654fff2c8186bca5c4198c7e85d3506780a049;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91682ccff5c108018e12da37ac58af482bb7a17a5d8b9e77d21cef710a4c7bb6a7dc50c029e11036c3b841f0f4d3b54df6bbf8a156aabcba76a54017e58a194de486dabbc20ea4c974be86f7de9a5ee66d39193f12a741fc4f36d57d00f2901d6c3b9d7c1054dbd1fc3fb47ed78026064;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4acee261cc08ac500aad2c8d788408aeb28d7d1a6ed81e7c25e2a112a78ad6c84b54cc80c2d9fc8a7d72377518e66c25e3505c19e0ed2b732960492175d729d78af54c59b97d3715a0423692f28bd84537516975d98c5c0d8d2334bb7015bda827750f2c0e87500786face980cbcb33fe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc51f44fbb6d08ab93cccf763f939b0ddb4f7d287a9645b10f256f9edc37ae313a768d4e439f80bcf0542504c2038a4b88b8599c8da2e10429f79d5db2c72456326f0665c97b7b73e4bed0c90adbc54075911019db27c982bf66e76dffccdc0a30369274b3b8d5d6ee17d47e498308737b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64246736e566ef49d1858d3e044f687c59a3778c3468cd573e3fbad69525ba8b8e04b426fbb6e3af3a9956c2df48b0f38e1db1575c1bebb468bc23029b68cfb98fbc39a69615e84e609ae3da4eae5263bafbba49ccc70e7eaff35534497c9db363b582099f3770053421ead88bdd290e2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b7b64a94951cb562809e00cf6fe04388ddfbeb5d22049d2542edaaff5e8b2213da90c4dfaf824c7091fadb744cd5d4eb169b52225119136d31b6f79407f99113999d4a4e33fbcc8f64d788f5a3e1fb24365082a2e675437e44ad282866d9e53dedc7a646b23991627d5bf88057787a9d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25b7b27ca122ca4052881aec48195c3aec26783f052cc442c7ba5bedb3d5f48f4224158205daa53fc06d6f9057f3e73c3a469e49cb720d1f669c057f56729ce43f2bf862b8b0d4fd0bcfc836c5e32908c34d8718205322cfc587a39c074a4830428f672ce31d1f20952dd8d841b747bea;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb3e11370d30fb527e02a5ab71647ac4807b0440539b39246831d968cb5a5dc15047bdf11b2397c1cd285658754bf1b160dcb597a3fb9c2500089d81dee3074143fabda45f818ee2183d09e97929ebf28e47eee31a1a3ca5ae8f0bfaf21e98bea531e5f41ab2b5e34c433fca6cf8f5a86;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb5378e4ed966c5123bc5c5e73fce501b8999631fa2c5460b104c99890536fca78562c1c75377794ff1b2bad6c1815850c17ddfe3f7e93ba1a6aaaf782b7751627b76f397bb557cb509fecfb72e7fc57e43748fb8bef795a0283560bac73bda496a1d9bec0850bc956afdfe5518b09030;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2eee2a26fd1c090397f5bdb46cb6251282d473b01f0ab50cde68a6ffa022a61d6d4dfd0d445d091570d2188e9d5cf36e97076f41f397b596ebf65de5729374bd6850c73d84c852888241f1a9a9a9441b9b409b3a22888e5e60202ab8acad683cb8ac67ead6dcf6678590527f8e4b632b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha901b8218d83744866f022eda777d05ddefc53cfa186bcfda1c07425812c1d75347bfa9ba86138059eb25de6af84f3a81bee177733eb392e4ff21b60019681cc731ece6450d8d6e154fbd2e2cf19578959619f39835545ebfdfdcb0a5ad14703babc13284801acb11ff1cd940b2bcc97;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97aa897463fab3806cbba3b9aa13afa4152fcbb7465376af26a07c315e4458b164a9577603103084a0d1f0db34fe2e42242eac0648a4309c47effb12896c9fca41bd987fe44d50e9cb20df92a1c051235adc79ae3a0c082360501ad9709423ec87edf433b668d10e345f89f376a1432b3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54a7e933b2769589e8d6a5304ba622c39d97461dbd3d19f82ca3b3e2717259c2281f32ad8c6d110225afa9ce724a99002e14c59100e22b4f60af0586f6c28489a71e02532abd3f6c32ec7f36f2b64d385d47d97ac64079e9dddecc20b519a286cef01cb902c766c8254bde766b6e02834;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h445025617e829131440e260307ff2480b1e0fe1b5c1c7cf56cce1d2916bcb55422c1630989bb79b883bf6cdc25b893a0b78696b9b6976ad1b2a5e0ef5b2be197281e8630c8e1b7b4e0b2af59c9d781bb037a5ce0c81d999d40c136d8bae8529020e630fb75c39c94c014c90ecbcf6d276;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf27b03a78a069ab14c867f299688770dc13f17bb9048dfdfb6809306f44465f3fd68deab530c1ae102eb6dc4094d06c8890067c9fe6e05cba49b8f190c454f2c7f7653d6122ad448703fe823670e44f752cd5da33cbd52e3cef53e790c4bc488556abde940b18d07def0b373918c27b3e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab4f010e1f5042537490a7ab0d80da6e40bcad66cea87346fba58b576abe73e19085d60a1b36de0ac275dbbddaa4625799e3ca40d7c1e417ca9fe5d250cd264723225122acbc3cf7cf2392a4e3c3169b29236a61e45c5cfcd09f5236710348538ec10449defdca506836114325cec75da;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h699daf8d8451eb40d72c5fb82e848f9e35d5fce3481cfa257dab5a1faf6453717cc3f8688a21d1957555c9e982e63100630a2e0d3dc91bb922e329be74a51c6ccc4c889dd8317e7edfbbf54ec5d4af3a96b6cc943232c0ee9f789f737ec9896e3528b1e8ded7a8f17efd73f5c1471ae63;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88de0fe248c1b2dbbedfcdc0863e42f4554d548a2b5b1a4abe8b8ec51356150b8d8a9105d5c5a71d5b8761b02d61703b5c789869800eb7bf02919d4ca1cf0ec92e067274e0962597a2bc899e15ea184b3493f60b852285c63cb235de816b2a5b3461e6ff1369bdab6a207ce27e042db0f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8fcbee65092956014cf81370c636e07e780febfbea7964f48670c54b334f81397815566ecc642f2dfb9c50a2bfe16c825e6bb19f1ed8d9c4f3c3a6925b217378b9e62a6ef1a544bba377faf27be497f6dd26716034662ba6f6f87983f6666da65bfa3bb09bbcc5350949e672f10e8888e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51bbe6af0fb9cb7742d156c48d6b3360996debcdf37d74946bda6b6b53d29561e9f2e3c39e00f6097785e7962955f15f8ce342c4ce4b740d353dc92cf43bdc3fc6e901d3d28abafd9b82739bf54540cd88c289a98f3f2c5dd285fd943b9045e8f49010924d2702df8cc28d9b8100a2a82;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he9a10615b9c3c689ee8bd90ac0cdbf6bb82317541cf3925257834c9acdd5528118eed581ab0f94bc4f092f190176c16ce731f4030ce54394394e1c6302febf7f3deee9241daa23ce0e904e8502633c44a283900426a8f05bc3a4cfa53e690db530b9c60d5eed5a402c47f99f8ffdea199;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h46f2d7f6b8d1aebae72645b060e336b2461e6d19a48bd9c9fc46d085de13d46a4d09643acee786bbb96f51c874ec7a76e2966919c89d58a2c1f21ac1f4274901d196b2caa1ffe532f504b4029234d273e515ab2ed06f76e7a9c41daf5ada8bcbb35e784ce6010dfac2f417d364a16120;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb89db796f9436170080a0cb525b4f0603f5427f72dc467d6880ac889a7fe918032adc4abc2149de693b7d2b412d75b9918a670bbfd9b3a009810515bf7e7e0c24b40cd314275b553782da92b4e54a830804398da601c6338fd57538827b1e7f6f5d16e8275abbd36c8932de8dacc08dbc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3300fce518f162fc837a64b076ed04f6bb407a026904a5082dd110fbfe149a29a5f74f7c389c2e9a484a33ad3e7d41118230c599e27ef30459ab13b549b1e81bf9cdad4d0b7cde0e1121600db6cc0838080887836399de2cd62884b1ca64c06acd321c3c56b79341b8513d1ce5114b852;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85cd6d269cbce09a0587401ebe8cea21990bdb2ea92d1a7dfa1212eb4be4815f097c5cba5427695c0e297026360e1d8a7c770a0f89880701778608452a924e4bfcc9556c43f8fd0626bdc1e7e03b09d7fc2f529c2de8f9d4c8953a9309f814f14a8833fb4b3eaa7def722587e61bbc2f5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3f6405d1402ba833307eb86306e4de1610b1b2ed4b7c21021bf97358df57868d4930bd8eda7586bdfafaf884344e6088bc4bd8ea30fa5e20bff1446f7653f0cd9b6af966be268e846740f5035f33be0d3d46d759f98e0fc790f1b7f0d330d093b15ac032add898a75fba8423b6d166c3c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56b23bc8d5e8737261fa4652e18722d636083deb6d2484fb1f9462ea6a21705bf772771f14ad1986825639285523d2fcafce5861268d66c95f670ad258f1b8f024ba5dc6973cf3674a079bda9f0c42c8a2d64a06104bdffc11a82d877c6280b3d6a8bd7e05fc35aa78e02725c550e655c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdcb9541b056309d8cceae3fab253e0da62ef437e607b2aff3ce3f060768c9e0f1214a826e232acc063724dedacb121cbc3daad47d40050a711448ba02eb0c6847c35bcaf015d3ed266fd9f26525c019aa05ae775d24f0a536de84726a4d6499744e8fe9bb44f51f6ceadf47077f8242c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdace6e3e499d6822c086c43b13de0e21fdf63d0abcfc2d8f060df7382d160275381d6b4dc70880f5e3383e75a40e43fecc12b86fcc161edd4f973dc4f3fdd6422caf1b9cc59a1c568103e9b48386ad99b8d0640a0ba6c7c6d6e213c1c2b8a9847d327a8cc159f3367916f37ddfabae4fe;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he195824f2f9d29fb061132fa58ef50e5e3ccd0d1ead52013b542292d079aaecc78801fdc08e3504f2f2b7ed46f2e79bb82145582354b95206bc081234a6f4147c112eb942c0e146f7cfbe6ffa31fb45d6db0cbe0a7e8feba6fb3e118ed6595293be1e57587b8cfca07ebc0de9cc0e3a57;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80f8a4ea4b3a0bcdeefe7ed23eb5dbeeeb2a47dea51f925587a077f6949349ac55054750a539ebeca48da548c286b98f680ebc0b353232e47c398ab9d333e3942a72b8ceea8d84c3028da490c30544cbf93859e11615e95976d2257d4977ce16a6f0c9534b3ac5b56b226ab2b16a9d0ce;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef9328d45bc7ab8794fecc48f707c28a155155798a971dadfc1061c7dbe70632286cc8392c9aa8f1811bfcd4a0ca77acc5f280b1880c1e5de8ba08fbb1b2165885e83a897734660094c9d60b0f6844c575d839a297da5ce11b248e0692826d45ffbc1b03c298f51fb94a03468006eaac4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65b4fb8e0b4db8b62d1067d0c76a571c9156b4e4c9ec66cc7e4f03761c9c8d327c09b9689e2f5111239ee4afbe7c02ad5bcddb94758085f459a08726fc9414ad15e7a4a9a7580f3fa85e6113b6ec8335e016c0123f009d32d456fe9ad0c4b8cee22066d5bea9b927c744e9bbf60a603d9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4e9d2d210f771f018c503fbf389ca0436e2493486307650df412651ed9e8a905935e58a6cd8d7b06e7e49d769648c805e6b6272aa323cfaa4aa2aa1f2f77fce2bef1ed664f9a5924a37a493aff9d212c22efaf5b6a3e1caef3eee50ec318af44adaa3b367ccd8b9d6ecfa12395d9dff1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he9c44026b6359a06ebfced70589c451ec3c14086604f955ed4aa32f96f73a127ec070d71b0274b85e69221de9d7ae82ad00cccc72a7d486203b6ca16d452dd8c8adb443f1738fdf0e903e0586c0990959fe9e93388ae1c0e644fae8a0d0c5378b5a10a5957e65346d3561145faf2a74a5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2d75d9f9eb94e2557ea46cb4e385a9eb449a505268dab5bc2296b05ae335f40821f760197b5d80830b4619d3d2795936c6d62aab645348dc24a298f7d4cfb7b546766287922b351a2a5808afa6008563666198b233b2d27ed6dc41c77d778f37399273b023c1c2363fbef0bad4da0d14;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h20a05abc323e722bcdc764e4b9a1c96ee76a8bf8b9ec4e4aa49689062717c001f6c25bbd913247b4a7d3fbfac687a8e56101934229b0a92b66e7f44a1b3328da61fd2182adefeb8dba5449f1bce0ccf29af9a11cdc48d6bc4e85d5782ac5590c86bb0793c5e13872521ce2e6cc4aa5cf7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25d45d7dbd566a7811f832cac0e9f453902fd6d88d2084cc54165067cf22163d54d945c37cc305a64d620232284bdb6583a05bd5e385c3e83464a5d6e1066f5478982fdf08afeaabc3da4a4c906c9cba07725d785888f15bf9ce07cb9feaeb833059d3f7a5cba5b71c58cbd831d7a7410;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he80358e964fb04fc75efc131aeba77c764ee4b01972818f1901dd29762518cf471470e5e21b0bb13c5cf2706037fa6327adb1d75177e72090937fd1ac5eef42795310036f54f8302b01ff5d88e8dc291a330e3eeaf6ac20d2ba548a4a9288c337be640631d4b458c88e1379bb1e2a41ba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb100a0b99d48c361b430a9e96df61d6c00a55df600debd2a8d61f064746a52276e62aa3e81aa01426c4b9b1f84d7ada74fe4b65b1a0697837d453ecbfa29d182d61043e844e67ff7b65ad0b88377fb1eb3dd446ee246da17531ddc0cec8a47cf511711804c4a8051bc7ec3f47f965a6db;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6aa49afdf382a70e880b75a90939f52fca7278c6fd6024eac17e7f5790b75a9d2e0f137b95dee45289fd43afb6f9175433f4b490900ff277c751e3a6e779305bde94443bb95103e8f2383586f9ef7fe06beea35b7501319518b6dfa1e94aa91fc55b28ead1938edc5557cad1cb227203;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9d364121fc3c0e14806bb3579c5f8137563ba7862b2e0d207792a0b3bd0757d01f606fa6883c6ac634c7b84478e960804006a3977212f581c9975959521309d873c725c3a340356378fa14aaecebca3e3a3e919aa9d98f20279f75d3a0866fbb37aa853c9435a682521fd41d2100c7d3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he786fd9d33be1eab6da682dd314b19f5c1d4ab4f9d086d74ceb9a4a36f1c8bdca6102e070356c89f126804328612b9b8dd30cee37bc330d69a68621ab61880af3ebe5265878235d763589ab0da96e47269ccdf1cc3cb1d79a63ebf4f58787a80098b0d1e9f15cfba54016876d56bf6347;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f7c0d6247763b12d5dd2022c039ada28b5d63bf2d8376186c6d472409c254aa4adaeb881b1e4ce4af1ec10220a2f1bb35c32e30fb05120a5d359dd3ade1102ca3ba9cae62f85e499a409c7b62f2a5f24b6393ed1153a11d69edb8f57e371a61f28d90f68b005151526e69dffa4d88b50;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h949e62c8ed37695938b909ec7b10c1b2353a54a930edd54e499e5962863dcc0aa6597915632b9d7a1840fa3f9d4d0a7e8bbf69e85e1054865002e7f549bc441759ee2d6a30a53f91ebb58c478891fe1c21e3dc351835a07dcd11ed501c3500c299388ba4e022a539b8ad257829e3f5f9c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h687128728d78aca25ea018601ef89a01002310a8e96f592bb43abcdacc28d3a0d74a23c57cbc9439014ee6a6451e4a9d0570fcb61e06f5c06394b8d72facc58e6786b690e176c7341d3ed79084a9e33487e099c51f360d6d0853846fba26758a603e6c68a6aa73e15ce147d91db9ba0d0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heeee40dd1cb97b7f12848f1d6505ee5bc5fe96928f5a7029effcc52489e07a29f9c5ea9d54f67cfc5ddfe4736ce09a3bf4b76f933abefa333c92f335a4f36b5c885ef90cfe75800d18c7836a40231bca8d5f70a24b87efce90deb9e92efdfe4c852caaebfa4b97203e0ced07e1709d324;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h493893e9c3b7ccb910eeea360b6184074b396b8002bf3abc4878426e413caefb3c2f2dbc8a1001186c5677bfcfaeb9e985f4b567e3e1960efc70b6cbeb82a2cc33a7004c7093aa3ab638e6f2bbc3326eb39ad431ead51087feb4cd041198d3240753394b5b96e3f4456c361fae3069251;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4a903bc590fc71cb13e15ba20ac52c31bb0a85a4cdf5ecf50f692452330a81071321ffae5fb3a4cb357eb28d7c7f92fd34a8ed7d0cc1dd74cf77c9617f3223f52043f4eb3db4b98007f7eaa251a9ea5cc9ec9a19caaa3e75a04f34afcce60ea637d253035f1955d6312118494a392802;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61bddc538283e571d4adf16665d438c9545487bee93b42b6df35077eb67d84f21d304d1e3aae537dd8d4882adcd68c70960eb76922a81227a0c3fc836d4e095eae37f66349ed421b31686046d7976af63f47416dae16ced67229a83f586eec9d11cdfd6ca647294e632426bf5dd3c2c21;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f21692489d4c360bb5d3b40695dd192fcf087d4570e0aa0c93f1cd7d5d65ae8899da202cd1d2a1cced29ba223ccd66a8ae50e14b704e1b49b7dc0238f02f30829a5b2a76dc4efd811368c59b6be55cdce8610d97451fe665c30ad7f199c7e764793bd451dbf9c069956d13cd5d0c2a11;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf91df504d72e0bff3c589d2e7fe1358eadc66185f38043a24d0e2330504cd0f873d67cb14c569d4ad7257508508dd96273a5157154ed672463b6a3e427fbd6a43bb042b7193b36df66b398722de113b34c43ac97e8cdce2ed88f33c1982900d2159b1a6303bfee77ff38477912951d6cc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5996029d86ff9d0800e2334d7f56fe001c83e0a942c9b5d98621f798e3a0087b875a67e24beb067f4bf30b9a64932c50c4bc1173141d7b1afd9cdb20da31c984b2826e7585ea3eda912d2defad88939217779b638f04c2ff5264fea7aaa7b9944e8ac3ff21500cc856dcaaab620a419ee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h63ee7511ab3f1ec9d65e34d2728ee104ae2b5efc4cc5820d4d79967c0cb0523c92d3d579a76a60d0de465a5fe061c27f187f26f96ad4c3729db2f0ae0a0a46448897184ab0f8b9c150d37caab4b697676766e9acebe13045633093b2ebcfb15097afc646e0adefc25221a0881e7b30020;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95715dc9e4f91b62bd8f5d434ba8dd1873e34eca94988e819b9681ba3d4bca7c28135e4d190779d15594353f45bbed2762d547987d356f63b255b5fcd1fa23818a416b265279337502959c8e4a28d1b4cb6d9e7efd22dcf99b02162cbcb5fed82d9185f70f4cc3303a5fe53f5eb1ed997;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff14c3ef9b6ba5c77167ab25aff2728b238734d74916251c6989c28b5bc470a30f3014899b6c0f1bae2dc8c87a57e38ad895c182ee720124285ff7e1953f6d41c013bf8afe1f3e5f8825cda109777c0c9ad02a7f69d699228969e4a4442c09865b4fcb3bfe3405287165c55591d7ff53;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7952d3e98bd11d4dbe0b588ab1cc8c65f94ade113567248e4849a5fc293c0e1fad8caaf79829603e0fdf51a5f70b2486a2f7b4ebd8064930661cc0ceb554a9e9b67bd44b81d67d117c39916652e8a199f3d97f482fd414ad0b67e46d859613e2bc8cd62601da28b55bbe9bd52c1db5227;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbe89c741b7bf0f487d61b72eb1328e212cdb533310fd6c4c13923c9a166567eedb32c6a4b5f2bc5aa7569d879963c31aef680ce1e540a2f02f03d62ceb9e286b1adb59c3c5e1530a8faf20c0ec2ed098545ac42057a5c028c3bed6a106c865a2b50301b03b033c0b0b4365d1a2839fe9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f7c5869a1cbb3750f5fae5ea5d870bd83b44b06f6c1e9084b2cb326817b4597a16d6e167fe93382a7d37b8759ec89c791ee889d6cbe47abffcfd14f842fb8b876e34292d3abe68e83d01de058fff96d755e83fe1bccaab0080561c479a167b8cf87628893452b8456d2c1bb469d800a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h828662c11b2bdd4570a25294db2610a997ef3e21b08c64486ecb1657bbba16cb3d9ce95b353c8b9b6e08c3164b56626477582631b5886b3f7f828f3231d2c939a2ef70893077b72cebe59cdfc55d6f7ff8b3e4d2a71e01d41def5419ba4ef1bacb5beae2b1135871f13316b44d787477d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2c9a1a4ec777be85ce2ea5c1418cc421e494c6494a40eb65fa1b72e6b8c394f1d8651f3daee2e9bb706224beda397cdb88a1b2bbdd68c94a91ea056ce4ee23060f69de0bb176f40f867deb4f4e5e2559bae2028a32fc0c76d7bbe2dcfa8245bd936425c44634108a33fe332bede4cc7ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a97ded995e73d39c84c4b67e53d87a4b6459f1c1da11001763e9c614007476e1d936f1f33c7ca6ed58f514f78f8871f14d4229b1cbe17f9e9c008c48302263371d116c8fdaca923ebc2b024081140f01bbfc80074f3267db8f69fa195a1398e71c17945002d4d2bc8557436198acebca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a121f8e6b6d36859705954b949e9fff0c66d0def278ba2ee5601bee52560f0172378448d201d6f7ca2e57977952503897f74fc83099f5c794cd61e2a4b1de00ad932313523ed4261cad2c235fdb1a084e350e77f68de638d7ae7c37447ae66f9ff9bc25a60ff5bf606aedbb997eaed45;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb342bd00414139ae78ffb5d51e66dfa8859f74c87cff0c7dc03b4aa610f1626be13a5ce9217d622319f1cd73e530839dd41f3ad4d45db7a8febaec3dec36fbba837938bd1600ffe38f21788d54feb25078425e4ea0afb993506907a74d5b94f588534c8b036dba6993cb3062732b45bd0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2e027c1e54f00b4d6f2b2b61368995bd346e342b65ecf9e2d166cd0450994505e6451f7c55da2aeb2c7d2e993df05a4d004b1d89f02fbd2b296f96ad3eb36d83db055409f0d8d2a6cd204db4a906a90dd93533b31a4323f8ec0fde7e71cdbdf0ce223315ba2df7d9cf0bd614af5914a6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h579b9b1b4e3f9c09c42bb729c32c2cf4dec4a46dd53d24e08171d4f642d2ef0f56c1f3c9de92b83f40bf1693f1f37876a24ab4eae1127d77a541dee3f6fc52f5149738bdc2920aa770cbdc1934ecad3ba76fd88b27e4285ff70ebbd429820ec9854c05d6ab82629d4880e1550a8afbdfb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71e4a8adfc06fee01a87e8fca84d9c36d921b6e624e1564d3192f2cd9f1d156b6cd18834e5b0bcef3260d308d9e5e4c92705d959d6d94ce1b9047773a490b71d4993d82b5e0f415359833c7d9b1ce268c5fad1fcbc379026b2eb3653f5da161dc009610049f917ab32de360fe0fe70886;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b9bf71deca4b76921d9526ca1077559539c849529133b84d567d35e6b42e4cbc6380e64a861fb1dd3f20db3d7912084e902778704712b511e0c6f0f3b0abf3f3b4687402bb8c12421541f00d2939d78527430d7c732fedda07bfd7e5741c0084d409b87a84b2f9caf30bd2a9c2c9b19;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca6124f9278010c790197ec5d96729da2ff3c7bb162659deecc54654f6863ad7fb43da350b00d5f0c3e9694dc0a4ce9eed434f1418f0af97ee4677ee6ca1bc73e7b998bf20f556c2ca4ddebc534be3e9c3e2eabe4462a667c1d990c36f0caf6bd1c31e44614df0a3db6c5a7b9b055e15b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5ae97e471a570ef61f4f0445c8eef86ed3310ddef41d66a9929eea01a05aa3f4c31eb52da2ad187334f7e7af683863dd96c450dd963a0f3760bd5e5508bdd219de6e6b401b165dde4f9d94319b4a41fa8ffb7201fd5aadb71bd4d4bff1ffdadfe2a92e72ac41ab4f359d1288b391073e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69cf91f982c59692f9c02bfdd642fee22fb74dac6784a0447c5d1a1a3bf53f6b300cbbcc3b55e9fa1351bbc64bd8eb3016fe6051805a8fb94e5da1a613c8800de2808bda34cf35277660f61c8e03056cd106968c70b64753ca0134e1d2e111169f2c66a21cd9177be076126929f6e1763;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d141c6c0f5095e78572ea4d06029dfd03a8fd3a82274686737ca2e67104a0fb253d4101476aa510722cc63ce8aca92e46ff49a07a0a52e9a84db3010032527f3ac55aa1ceec3b29eff374d338f5ca1b7a8e658d23890f3d8a5554d2266c8cb9e39322de2137ade7ed7504765c60c0f66;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf03bef8f81972d802069210543bae9124d43bb15d07b6969c6e0891ecb7a05e20ede912421f6c86ddad5365c04e4976c2fba6b45923466a336d1dca57b5302f300da42fc6dd4fe2806a4d698c3d8eb0b306648afe8469b7afa3398cbe99f15c98d1832153c881668ec6957fce187847f6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e0ff7788799cf0ef2958ba6efe1d18144e8e69b41dd1d1606bc5e0bc0db2c00f3a4c15b28c03979a0239fce8e2e83af7711182e6ecba6c866aff9434de92ff9613c86426d00fbffcd0e02e5495e5b174a586d4650104dac1a37beafbb7de9d86f1fcaf6c5d789560bc2da6d89fc31d93;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7756d5e0e4ddfb93de27751c06aa2da209d82a350559c7ceca1cbc7fba5e3ec75fd6f6fa877e6f369fd39fba7c987d25c219715a7b527dae07f30b2c478f71deffbd27c2dda89636eead1277bdf1608391a3661fc9c388abe5e9906cd62800b327325d49c3eca8b1f8c94b1ffbc39937d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc9095635e2da8639aeae43181e57eaf2ce7cb5c035d386090c711ce77554bbba2b41c5d19c92c3712cd6f59f94be0ef03cb8b57cc72bb94b1c48ae866c9d8b2586549d5612bf6b735e0b5c9eb5e09c859fd7826f3f8f1a18dd959173a01231fb849ee14a474d6d43a004db318ff06edf2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb607bd854743d081e7ac06e63539370b0e15851cc249dabda44213738428d1424611b09ee0eda6235d3082af854dd9adc1c73adb536f3d0ce53a9d4aae4ee3833c4c5bf45075287ebac6c1f5060d7f820ef4e1b09936df9c9193bd150f53532e871612fa586c81d1e0ca0c5dab365931;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89a61bfe0862a3c2198c22ccf02108a766b87b0683b29e093be7916fafd6f8cab7a0f5ee91c2ae3f1b036abb29c113e0e3ce46be044ab85cb117f0cf6a1caaaf71c0d04592ad9fd68ab5e37d9bbcb2c864a1ee0874bc7c070a2a1fbe417eca63682135ca6a87db880be5032c3255c170a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcab6246b31153e88f7deb85a512ed5609e78ecffdbdb87ecea393b35372f8a4ffdfb6a3ae2cab9f135e8b926dc65963067cbb9038aa5d074dd5510bebc4bb6d07826bbd5428694061a76df05b6149fea9059f3e3235a02bbfeb3e2574b3dc2fde40d1c2e1cd851b30246f4b1daf7a7994;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a5b500e13936bc508a1e5e1530ac70fbcb459a81d4853dfcab4928592feb0df170b8aa52a098b60fc3f63cc058e095bb22420f76a258a1a2420d3184bbbbad264cc67aaac6872051fa63ba01eefab954afc8f7e68b8eab551c9c26c472c32290598c86a59d831c2fee6237030ac8c735;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf977e0ef4c721b1a6ab68952338a99551f639503840ac116f0a11f54dfca598198f14209b145e7845ef402f8751bcf95184fe542b6f160fa1412cbc4d2af472395ef1505eec06b7eaf458d5833b46efc16f1f4aedca50ba0f1a4d4b4bb13221c493c83180c2bb4b4ebb6ddccf889af197;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4dadbfd4b1590facf32d1c4898fd3241ae991aab04ebef2cdf7962a74e09d8b46da4437b95e276be12932f763191ce97d7a5962ee0918eb4dd039dd40df9210c6e8f20dd70b1695d992f482f60cb5324871f6f12e90fb01605aad988191e4d0c8ea1017b765e7f813fdf22a0adb957d73;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h537ac7f551ba04c08d075f04c136ce3d5b618797719c10a08cd6cd0f4eff0da4ac5d01844592ac276ac570f558b8036e75f98ed3aed6cf235b3c5cb1e581270ddbee2fed05fdd1aaff98e0e8698f56b9a973637be0b6baed1fb8e7e01297e5e46412fb86d32ae6cf7925b7b0dfa4099;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1c363b430a1e25f6094cc416e52497ae7dd887d18333674fd28531408145a9dd055d9dddc4c29615493270fc7c25d2200af8250aaaa2e61ff1d1a6fd758e86c8df20381911c68485c707a287783634e12920456be37aa69827affc24906c2879485ecd62528078eea65c4941e0d51725;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93594b5988b66a9c61ca9c0be57872fd1a02d5f94df21adde469deaea9aee74b884b34a61c05f4e585a525f1eba0c66b363f2309d1a682dd0b6544b445cce42c598a6df05e5209f1f3cd34d6e9e73253bed4b5a2bcd3ed32ac0e8bd67b69171a12cba5d8ed059bf013629b7dd71d154cf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ced10057c521b41fbab611fb78d4a2f9e2e3dd26d202ee1e67c9798a2d671357f1f0176ab88ca050520fe4b2c4a35c6eb33177561ee4ef1e9a4540a829a9f3374c6f8d39057e903d11629020274b64db09509c0c069e60bbeb488b447da857a2b46ff1ae5603904ca7a428abf93a8508;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1dd67272d2541d46c1eb48817de824c640f9a9e4a2516acdccd0f897eeda770cca8e1312996b646811c3b258a1289c33d98c32c140cb49295b506d678fa811765ec19119912726c43835e5cd19a5c81c160b19e42c28db0ccfc4e2bc9cb28f571135fb3b3c27a27f9560238c970946c6e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef7536ba66b4edd111857944427f4e7f71d4d3fccb0f77918d7d71738d5cc2a989a4f21c41973a1b99a16ff005a6e89a6a3f9947a4c65065960b039e0ea06b9271886079d7d92c098e16af67160bd1784c9882e1ae4d21c1d8373a1f5279d381a25c816b30c4701b2d37d6445cc75f181;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69c8cd09ed935ea5e65a68104dff5c0d68929c1f34397d786777f494436b2a3f73a5fe956ec40bf0ff079585e16411d25aa87874939ca400c124c1f213754b17c23e57bd898711a54a3f2c146ab11f4a348f2484db5b8a1a3ae606f6b37cc48368194a372e1ef2319ec09936247aa5c4c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h839725efdbef83f3985eef5141b1333ed9ae50fe57fb3946bf2e0dac57fce28ab3ab2e1045a7eb453e9f199c9b9225d2bb50871d91e93bbaa0dc7ee5ad850312456367020cbbcb59359fc20037db6bc552ac39ebd7b29a84d1eb104c89a2f1ac789e349bd437fb81ecaacf69c444aa8d2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d812a7bf5d1478926b9d21c786bd131779eaba69b4b70af6d8701a59677bcd43eeb73667040a6886eb4e3746ae730dde2181ca7e26535ff9978f9f63a11948cb8fc3ddeaf7bf7eca86b2b0f24c9375502413333564584286da5d020d34bd21e22a8a0916a58eb92494435d4099916497;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd5080e89d49d53290ee0232f2e15e8a888538e6e84d835e9ae7095befb4297ee742b656423d87dd908351bdd6821ee9775bdc50c2aacce79f9a216bcf5f8029c42c969b92edd88cc69d3d7fee91df64d441fb15234126bd1a8af15a5c680529b059db616aac224a8a4aa92fb9e07cd11;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73e1946f06a09e2e4bebc425f3225c3310846f4454e9493a5b78a711e22025437be5b1f31af5f2698725020413b2cdeb3899c6292570c28d2d661fe55762e9ddf93cc971f770a00584ae38e9da99cf453e87bcfc979a35efa1c868ba0e7331a0d4fd430d4ebe1e8483748747db796f12e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he49f3d1ed4af93af64376e6f3802faeccabc3ecbe7e466ab72a21b3896290f4a38a68914a76121dc171465f588468464dccfb1c1fe2bc104e4c95d90537e24842ded8994dc24fda1103d96f807932bf31533f49789fecf7dc30b423718ef3ddfdc850dcf35527971beb0dde74e709d8ea;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90a7271466087d3777f4df1ffbcbf63525c77ee0024a66d335a7ad13982c9e6bb8db00c99b794a7e827e5f827dc74ac1c456da471351f22a4a0fef252574b4d7e86d1ec1a289da7a8e0a5870d8c82eaa6ffc624df6f4d0e9543fae72bb9b017debb12e375fa71c6264aad445721e58f33;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h432ded65d9e4bd8e5303c6b8009b3dc8cafbd7d00c83b21551f44d8408908a9d0d11ef6c0b5a52b407ffc94e291b9d05a8274e1dc5fb162520c5fbe993cbcba04f676f9838259fe9f4e4bbf88c1cda2d0b7b6655141a4a1fb1e5e300be70f35400c85162888690f7c6d37ae89e36fae7d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h53b7f74aa9950f8100e8b3e929f79b0346bc2de8c7c31e78046b3d1aef180f935b81e69fd861cf985b217c1b6c695f49d544a99e82a08349a79021b0cb31eef6deab6bafd749769a8757ed9d82d0628f9345efb28ff34e3673141738da7ec0c50913b82704e85f959390c59459e4942ee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc00429a8e90f191289d0236fe32d9444e6abc422ce64f5f8205b4ab9fc3418c7c8cc926b84410323c6ab2d86acdb4f84da721681d5cbdc7dcafbc11687b72dde2702d52257e32958df0e2631004056c461099d8c514aba69131fbff8a54b8e32831cdfaab52bd7cebf92ad64b47e650ad;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5be9a7388048677dd9acb14aee9acd62f038a1736a58233bbd7025d19863df4629aa04b0975863fdfc2a27a7f39e43b4fe9413d77763410200a8844f14c9a5104ddfb2545a91e4f6ce14c5ecda4c62004a19719e4a2ba927260afb7a7a0c7f3ff884f985942a04665415ab877254b8c52;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5eda03fbd3e9d322a7dc3ef7278a9a923072706c208a6a2915fbe060ee8e5f8abcc6441891eb7d1ada03f1bee019eb5b30d5aa3bb5925e410c1e270a787381aef95149485370673eb0520e07722182c19db1d4cc4d7bfd2dd593f63b80e5b6006a323ccaa51f6a378026f4a9022eb7294;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d3eb39555e8dc5d4959fa034930a085a9b82b97e276842624c38cf2757abea2f7e0fe624f7c8c72b0eb5e84130749c28c6320ccc60105d3950a4ff4cf9fdb1bc08f2d46585dd50e5748054bdb8c3b2f34ee413c1bb6bfbe5b1130ffc418c228f79a1622b255107a01d2b2c7753394118;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he9b8828b8140005d9b9a8579bbf7124f8f4cd3d17cca17f4581915141234a9b03c30293c834fcf357ff6fa8c8cf894c210af0a769caff7866ceed829d487e35d1ee8116d78f005723ad1cbf22038ef1329ed279951048ed6fc3789dbf1a70fc060fa4d5a498f5fefada7f14c92d7b2b70;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb25b1990c2c868f269fa66fcf9631c06a8794f926ced5a89465e8c2d3b1ee6588cfd17c9b18161db94c0db49b03f80f68e916cdba788bdeac682eb5fa0f954778518deb9d22946db35a693916100e38f282e0611ce2f5a7474b11beaf5642d2e81934e9ea5246fa1aab5116b867e20e7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24d9d572f72e004aa9bfeb966fedc488621a10405f3e365eadd2551112ee963a75dfaeb2a1d45cfe39ce7aeeebc078d9806bceb0d4259072d90ad7c27ae008d715e1219b517b37c132e183d1154b5a7124a195fc831565f518db3bfb0d6dddc56214400fd19f8dee76f93e6cbf0bfeb96;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3be33ad1afe6880344275d8eed762198f29abd30cca48bd0d64477f56baf3c7b271b716d77094b4f839f4a85dcfef39961801a262a0750ddc0dcc5247640a139f4615cd778ceb143f09d89ee2c7110e20ed6bc574694c76db16464f45a1f8d6a3b0900509d08c38306aab43c9a6893dce;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h35c8775ca2a47877cf5803fc0e0007263958723d02d85b19d22f2a0a9d53de19c335cb306dcbb6910bf9a1d8eafcc3282367c874d5081466b160f84e6bdd0a61d052950c4a022fca5c4bd9b62a8550a129047e9828f9733974fd36b417ceaebb01525572eff2961d850450ab966cb095e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43d58a3dad2bda1089eea666237820da58f71e271d5d9053308e81e6d5d8265881494dc98cfd726202e6db5f81fb79fc36cfab0969ef05526f571e4bef832b0b44341380d194ceef287c3b6126405e410089cd8343b324df37e023a12928e97b3680705e5f00d71dde85e158395c9092d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h219872ed1354d4da105c095c167baaf407db81195935fa90e02a76c7a126f1059643b80fe0a8bb1b34938aa97b61b1fc433e12d14f5cd5742fa6c019ee1a33d30a5cd60f1e61a707b710fed35cca7f07af46ec23bdacc67fdcec529447304d15652e1ef59a08132996abec6b717978f3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f2baac6909bc75eceb6c81aeb413b2f4c0ed14bf96e452745c8cb2ff24dd08b0735748ea87e9504b8f08204dadd8e05bf5045838d7c887e55981e0380552ed26658931a034d109eef26b844789858104882a338854b19ed37ace1882dd1ea1dd656fe0fcb9846c605e1c0d43291e9e62;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a6fb8d74458c28b669bc0d09154ebd9f4eb9f25a11fd4077568d33f22e17335a877de49bcc485dfff2353dfc1cc89f662d834c703d2e96eadbf1af7f0893c29295b5ef2b5e03d4158cf3c31cd3e81e3c8d6866d79281804b0d2d64501c48068670fcd5aec476196c16b7978d4d2281ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1fadf2452b5cbe42804e0fda9bae430e1206cc7feb131974f637110ba4ec1ed71bae8c9c4f4f8295b12b0de58dfa2117de5e81b1ecb3a5fe49e57804d72c416285f7e60e6ba2ae230ba5e51a9a821a4156480efd2bff93e06994c3de459f370da8ff2383c375e15235b17aeb4b06ddfa7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51c7790f82165d1b56faf8db3ad5ac1bc28f7a52e96d14b72b3011d308f38cf07521b5f21d810050f05c6ea3770f4f691da0008ce0398b9e5d680c39e0d9af44047c66ee95156f8919e0e3140ae6b68f532431b80b77a17ec1f728c5597aeec978e6b42185992771a54b1f64cef793b84;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf748397feda3ac5d833ef9183b5a0144126858dfe7233b8a612bd1dd5280c80174dd994894bbb673eb6af4f97052a20b4812c01d9eb2dad76d1c632e17e42c05c4a79cecb409ea1b11d20cfe386a5541cf522f9f87e0023e32ffcbc7e0846f4c0d69de2f49dda131e8201e19420d926ef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h123fd6498ea9749f98afb47e808adc8ec0b011fe9def65e14e6f299fb911ba34568ade271250a183d92c3d8803aa1654943fcfd1bf473e0d61bbbfba77015d96ebcfcf03e7671cd14ff7341590871a81f79096d4623d724acf56ff160be4a86cb54c1d1614061aed3a8909bb32724dd1b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37d90dee6b1635105287c9f5839986a914d753507bb3b9a0e8868305beb7b91d67e419f2ca561f76dccdceabc9a4eba2a878c42ecea87c8d6d7736a2d31a3542585408ed8c1b86183a4bd7fe138887378ffda46b5ca891a8208ce753038945b9fb71c78e2e7da1a9edfef8617a16ece2b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdadb132a15a9e38e1fe2ef7b3fcc80b1ec1146748e467026a9403ce348545600b60a2fd1eff185c939c3f641379937e0e05e368eea22b68682b031b1fcf59f035ed02ac8609c66ca88280969dbdcf2e13d4d5613714ff9dfc7251c1fa62a0e4655921dd6c6ce4b1ebd3a8c822a14798ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdde6611c7dcf1c4d9436d3d66b30a56049011ebdacecc42a49d2308337eb44af8c6411e592a14cfb8648a0a321f1914ff81a718d1ce5eeb06a607fd91f9186724d8c2d415747928dc55f2fba78c4b6a5a55bd0a40bb48f6e6b4b285ef374470380a185c7956f7938637fde2c1946ef343;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8ea605a547550311ba621f0f717efc583502e7df5cd6f895290c631bdda14468d892ee8fa7591262017c850118d77e617d3ed8f862b946cbd84f93667c7e4d8dac5a56f0fb7103a5b30931de6c85913320da7655544e1d64f74837bc521ec40aeba3361dbdff575326d8c238f34147e1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43ad4f0612a0db813a7d16cd39b1d2b9edf5b5f87f9f00561a4c7786e7be0173909fe8a4c0530dfd65b77f74d80e847807f83e7e9f10d0aca27eb8086d080337a794ad402098e1a0c10f87ebf53420bcf1452354d0a5293cddb7d2c30c844fdd52b83e135b889ea210521ac6b9f672e77;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb2cac5f81d3368c2904003bb0a69ee8d3a19dd086a9d1dcdbf8b704b89838da4e33c765362de20bd9524e8bc8b39b5fcef31c1c47cc81bddc3d296e7b389204cc90811392ae6497c9f65249ef8c528b78cd9d143abd70be915eb786fde77f4cb20b2a048fc11167afdf3568d2d3668b0e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a02c17bdd19b7a83aa18092e4bb69199cf793789bae4e1e23772083addf3fac93b1c9d9f50d0975c9a622c0a430864ae78c6f1523663ac1fcf2386aaf24509c2505dd1d6b267eb0fde569da88f9aa254a102f9ca5ce8f74dff4fa65ea290edc89ded51fb5b474bdd646a5e11f880bdec;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf66ea025c7dd9210f93f091dc7853abe8fb75b44804fb84f97581067bf67e2d5a4606d9c46ca0735aacdedc279ee65dbe45c115566976e14a2b620ce0e7c859d4db6e023f9d47d4b18f82059b8923ef237d419d7fbadb2891b95a29633a39381f6e30da6a6f06f978c33c9bb05ffc630;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92dd80b69a77b46c1ae171702fe372e6a37d2ee483d6c95311752c23f22703d283a61da4c9db6aa508db4f6bb15a4e093df54a2a8babd2b5ad1a2170b40895630afbf1d6034904907579c95e0b463e36221475c47f260dffcb67f07a696f32b291b3dfb34d5e4c35a207654c1f79fb839;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9449cfc704174a96b2dd3c98342c7be16fb17fc1780d12202dff4ea2bc18dced3d1a9da972ffd492fc8e0b765d868082da74f9f8db2dd2ba44cc8a8bdc3477db8542621da85b511220e9b3a9d5b39c5ac92d9424f457ee52f497666a6ec3fa868765d3029831ad56f41067929ee9379c7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f7591d02b487b77a12b1b75aa0c28ec2ec3d0fd4f47ad7ad5bb3567fdcf291cd1a3474a924c89b545fbfd8d0171e9b339f16a7ede6e6a8a1ab612d959f1aacc89791e5e5de4210cb8945f0f3623a84d2c61c233663e69622fad620e234f9e143554d368c50b9526020e0e0b8942a76ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h446004b712ec48f87a617e1d169af53b1eec1e5faa80a03959afd5cd515c271199638f577abc693b7d1e3f106185c3ddfb36f1509b8320e458a65d36493aba9123f9051c4de2e36b8b344644ca2b0ced32de16133101e0deccba869fe4e9a54c596fae4e03163b4827b900b1707492ecf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h941054f04ab289e78dccab3248e4fb791569bd25d6cd61a19b0775631c2d5481582b652f057721ca0cb4f88949d8edad5d907bdf95fd7dec424424fa1b5f2e9974f94e6b3419b10a5cf097b15543412300a61b1b8517410d0a797dea6e8b4f610876431c3626dad1af1453c868391f277;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he136c9742d3784307d1d816682a68962c2d1fbbc8bbe0d3e4e40635c40def5ddb45a3c4de88e9ecc18031e356b6bb88a386a09500c4c19bccce780b7221ca0f1c610a197695c806d07c1ebffab77e4da5a5676bbf405d7a18f37eb2b20b549b80b75ddf5b03f69044c91e79c94b088a61;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7963484635ccfbf144d499c3bfad4eb5a926186f2386c6fe127dd6f1ea02e9a1c3b760e9f0bb4f3d43535b4d76d55ce1cba1b13c895e490c866b32b5f3a01d140cbecbda275021fa5137613c9e0310ccff376990c5a735eeb5aa9edf17fcf958f486d419d57d6a2fa2529db8bb049b686;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdbd208f80e4fd8d363ce9f61f86e498416ec886f41aa98c2aba3cea57aafe45b94854cbef39f4c340de713f3a9e0172f79674df7236ba004ebaef2f8477dea0930cf7f6b2c9b51ed86e9896045488a584139149cee2d983c401248c887ae7d1b7cbe562583244eaa0d57b98b35ac0d2df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd440e580ee5ca9aedff603e8bc8b10b081df8eb8ad0f3a27db1d92e652ae03eee790c64de74b9150dc535c95a90ce2bef5c8cc06dd7e4f2d00963dfc11167bb862fd38c2a89e9f4a1ede5de4e56f9b48218f3c46a659ada295e20351d120d9690ce119e152190d67dd1840ea41217fd5b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb63f38fd1a818433088b341293dc31f36d0654ffe0d77f36b7789290e4479384c58abc533bd76026811dc14b0479def84a8c2f905cd5e73a328706ed5a745192f68b5ac56795f3cd450454ac42448368bc1f1de988968fff2682da169c54411cff05a58d52802284f03e0f5f2083d00c5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h245ca5dd446fafc32ea8c99e764d4a1f412055ceb05d811a9f800ec5294dd192f720c3a983110cb1456a25a448dc0770dc9a03982ac6867e0930cc02cb28cb0f6e8b0e863096c75df571e7145c0d71e187fdd9582c1025165ce0f46bcd643fdee0f551cc8627e776c4a7a81dd8b36ee68;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb030f480ebff65e68b150186648444ca34051e1e1f7bfd9804873d16777bf06b0b6270606a6557f882cbb8d08a25127ca9ed2c71576daf07d3f8ea6e5badfcce14aa4e2bf7e986dea3b50af139de8ded5267beb4f692e1bb5b3e779233c578680199a4bbf860b84e2f8eb1ed4b63362a8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3bcd382a65c8251341cbc0970e43d5d54343d65c9b1cebbce34ddf6a9ec4e53d3c58fb59e1bcd4c4c398f686adb8a37c86dc390fd3c15bfd19bd84a9e1b8b1939cac72f8ff4ca4f742661d85a8998b77363fcb888b38e106f98ecc6233d4d9f84c8fcd9670cdbb0360d8345a3f5be87c5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d85a5a753db1cd7b2b62d40936d65ae3fd8ccffdbce1b1b556a652ba39266f8c42cf8d42a1bfa8889b271ffdbbffc4360a87ac8fbb74132fb469f577a6f549a9222328aec9f821c380ccb2485e5ce3772bdcb8e506ffe4f61d3041a0f55f7adbe5eeb7f8c59eb2e8459d9c7291e4495d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14a70c4dc97279daf21a90421110dd4f219d7dae6f1b7b4a548f466635e54f23437eb8b9502f0f7fedb79308c3b3d39ed99d9d647985093905420cf21a15234b23dc36f56a032227f269d84691e7ccb527638c03bdba53a7162f5f502069c1e8035afa121a78ea22c5f060160b4871596;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3902a1924714803ce0ca6d19e046ff72f8acd1dc85b2c18396539a65b8f869a96bbe61eaeeb5a4099464ae75310311dff25fdec4f4c0c4c7f7a90811281ba8193a27f3ae3cca54cfb6ce514599f8a2135bf0f484c130ac1a09516d03a63ae96900e60a2edeb77c909a7b3162197182074;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h776662fc9c691955f6d3e26676de68d5e706761235b2f42ad55d8cb91494e5d823aaec1cfb33fa8aaf6617263893d4884ab22064f8dd63650aa4a22ae630ea02868ddb88d6dd4023a5445ba0d5b49c587a1feab7b9b6f8ff3f71d0e980d280baf1aaeca00683783d0558e3ab401f949ba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb058d7c1a711dd914c78dc82acea109c7063d49ebcfce923f8cecbefe2a05c2931bf1712ab8e62ed120464a7b64e9f739ec2fa48b590e690060ab94f2f0bcb6c91d9311f2aa79a33040308ed9faa255f3377234fef1af6ef46ffbd08ab90f0cc3b290e497735ddcc0dc2fb68da544e54c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0fb83231698ccd6011a7b0c6f68e2b48ea4360d67e22f94a191117b231039e23ade4f5425dcc3fd36dbe4da103bc7dbb67aa810f2363a82afeab0dc3d77fea4351621a0e6b1f52589d856051ad0569bb29b5310563ab5941c440a19ed8bd9555d4f84954511f85914ff59f432a6c1a84;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h716e4f373bca556613134a15c206e04f55d0f149e0b6a6ba2f3c924bd612fce12430cdb72d32ef5f5326dbc0c81a0d145e222b42db2739c9bb09a0f42a66b9e6d17bf938d219842c82ab609bde2ff2813b1cf761d246d7929f965b95c36678239d3e3515a0e48d1694772bb73c94862d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb75f74b65bea87981ab0227b9dac077cafab18f2c76c5d0c28108e62050e4cfa28ccc77c5d6e1d1c8b4797aa0c7d8fc0c4d7b0c48e717d497c98fbd3e15a85c80dfa14d04d903504a4a14dfd6eb5067c008dfbae0987abccb21b2583047c764cd2218adf8ca8154ea9b2a47865bbde58b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48852365854fcaf1440ea638ecb0870214567add87d73f271dc5b53f2b8a7b17db9492b27f9ee05b01f27d0e21813729c83193214e540a8b1d7e28d6a060a559501fdb5dea3b2c857f6bb2e38a6d9523372639db7f0155846dfd7880e498b4587c339988a841f8a6262a61a3aa7d2d851;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc946b6040bbccb17a3c8ff3d5a95525643ec0bb58bc21aaa9c3e1442ac772eeb89b032c3ed1c67d29a0feb023edc811a3024fec6048df6f66922af309e2b491ded92c45af98133ac87d1dd60496ee45f7f46236413dc7b8b005d9ef1434344b0463caecbd6cd8d407cd5730c53ec1c4ec;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfcacfb4c38dab866b3002cd8c27f105b3f3d43795a99186ff982b1ddaef7609e2601df838d5cd8c11378de13c8552abff1ed56f8f6dc13a53d676c98c80da17e79f0942fb7100c086afcc1031a525d6e7c4097656567cf20e490b8c275273d881387fdd45da6344dc7315543f8adcdfb2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb697cd0f2bc85c55a38b70f63a8cdfe82bb162f40a0a0353043e7e704bb95cd054a7d4561fe1399899ae5b662fb880d3a107379c6ced34d8ca960673d2ec3bc97470c3a492a1477653583eb9253b4b837a6f0aeecd84acba93e231d2a2a811fe74d44108f7f3f0f53bc61a6b280ef7f1e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9447f66ce34aece32d8861e5a296418d7b68002a5919b96b616424996d58f7805dcb8d2ee757d1255a1ee2302d94de87e0b64eb3240a62408a8616dd2e7974ec9ab3740f8f64820751de98702dad97ab5d6ded80b091eac369c4c30c5de02db4ab0f3fd3fc4b4fa67d32055b8e5cdb471;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd2f8c5f2eb34992bff60dce4246426fd6ae96bb92b954c4062c0791203317e1adc9f8d309a224a4e23b435d06d4b3d3458ca58bcbe63a9c6c661133a661ba2aa689db694ee183f8f8338fcfd24393c1ab9a0c13a84ba4a23853c043b0d47027011b1140f319056a8b7a342157d507deb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6618fe9d19b324aa3dccac51a0b1f25fc75e91918a84d9dec082f07e061d72e81ab71d2a44ec37305d54bc4c9937fad2280b9345443dee4dacadb2825f341516b43fe3b6db1c1f169180d4b9ec3e3b565e2493b0ad570117dd801659566f63003a1263b0347b16d11a330a0874f4de08b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd3b7ad36b7ddb69cf7a499621502719515f55fd290c0386b760617339b34569c242026a841611d8a67faa4116652f6376b833620c25775e798ccf0d5495fbcd1899861c873c4937b11fbbcf18fa43b7db99cc689c8b275db66ea19af8aa5cc4c6c33d48f0eefe9c3b84a0e2361a7215a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a6083299918ccec90dd457898f9c2959a930bc2b9eb5a063cdbdb38bd968500f062b3ba631f2886abd56998ebca294f1edfb1dc59d68aad7ef387c96028bf3f0e6d8bf4c04121b505797aa0aaa50d636489ee394d6111245e07373f6e1891babb9245678bc44965f3f882feaa05365c0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h628b2b58357b8563baaeb4032ea1438813220c2cf56f61060e10af0881b3eaa0e8c89eba84164c236d841ca0827f2d286e4c8ea0e9e266f5fe7aac5c73f526ebc447a5ed651614815967c0c3c475093fd4fcd7dc8adbcec9929ab617ef7c9bc188d81ea665e6410ba272575f894067d99;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1efc81ace40064a43a9f97b5cc61fca5f1d9b1d9c5b8ca19f1b2a84b93f4ceb807d0a114d1e6a6f9a9221ef70ff525bd65db3f57726bd700b118bb31bf65b4c741292f8a92e3e5b4cddf25f7a48142ca4d93866e2679470f07fc1240c52e54f57213887a5267e89ca9e20acf4e5c6679;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5537b59becf4afad6521410ad4a58b0474e0c9a1a8662595a9c447b05b11508ebe34ad2ac0fc7c97d89c421863316f156fd8f35a77f2f8d7e75d79c98fb6619828a773175cf17116d1d14c2702ada85dc8fb1345dcd91c22e97d0a2f8d8ac1351efcb579b573858b4ef390d1e65af803;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4241cffbfa020b4dafc0b92c395d980b5f20cfd7048504d0ff7280e643638d039bd66987b438220cdf748ee50d03c756b87eeddae886d42c8682c5460820f0e2debd3f201544a1ef0ed786adbe5b1424ff213e8e5342f6d334f66ea6cde74fd3de4808a513ab081248fe0f47ba267759a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he83959a94c160e755260e90aab9175d0dbb1f5f0192775214ec73a162361ccccc03a37ea8b863643e6324379d2440c967b0b2937c99734560ef98847f47c4f3fde35248ffccb1663dea40c79b7b48ba775a0c3cfc4b389199d4b768026d21f18342bf4e0d62407f0b5a050e977645983a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef7bc36f8d24add9a1a648a2428d93cae6de4c5bc22e55120b13187884641dc44a9f2aa7b04e264473baf9024675191955605c0331a924f9290956675e0ece36f219c127f49763a7ae7a737fb402996a0dae91afe860d2b4d0b0642f619195277a032ff22f5e751ca7dfe7a018b315a71;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h688cdbcc6f7f3d4b9adda7af2ed26c5ad6905a04ea0efaaa4df8a8645209b980f8ae9ad823ece6024b68f4116dc07f769efa6a4aa8a2b03905f313ce22e4e83439f65ad3a83c2218bf96460c93e6997c55d4dff34a7af0884d80edac2f561bdc00a5fad8232365e28802254e6e96cd9a5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h507e594177073503d8626741f38d09df5a143111d77467fabe9a7f8bdb9a67f46ebd13adc19885cdf975835f2d4e096835b34f45f8d0f6408638960197b26c88a6f458a8d25dfb314d1161ce211a4f5870ea45478393ee114f9636a50c8ce46187477c87992f3d80131ffba7901fced27;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49f05f0c2951b8e8cb9f64d461c5538a23b2852be90688f3aeb97d1b2519f47c3bfe2557f2048b60795d3f1416852085b0537048496416495343ded915778f9aac419a97f994b223f8851cdff2de42e531af99e226817ac3325cfe948de44dcb7d73ebfae9e973602b879122c03b4fb51;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf651d31ba4c8a8c5f3660a607dc49a90b9f48b7bddf1f53d498dde95c2cb3a19b322bd17163f8e9b41f6549b1c81265c09ffd18cf4de71f61182365a165d1bbc65d79334207a4b1947164a42d4993602e032c7466b127674dc14b1a4a55d85d9e347804b5173701180ff5e296c398298;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbd138ae6b63a1800a0ecba6b5a439514622fac4813b48ede64303b7afd05fcf9d8f2b7663e773b7a7774abe0c3202c07ef89d8c37d0e48726b8a4f269c50844dd2816d51486b1be8c492a9cc9c2a64f09e7d88392e550a6098db8c7d755ba2e51eb804def933f598939fd31b38cd3ed6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h646b5dbe0bdbb61e80100ce36f77fbe01d4f8c8342c5fbd781ff45963b7bdc862ea3f7efb69fe4b2da948f5ef51429f29b62a24e5f0dafb5bfc8dc3a6da0052396ad2cac0decd8b0a4c26c399f396901e9f87efd51edf86ad84a151fc8380d588aa3c35aa8e0211f8ef0349c89a3da9d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3bcc0d361f5245a4638f398a9abe0f26c4b02a2e8c54e10aa00b44fbf1135f8bebc34cb30571d34946c7528ba52602dfa630583527c94d15de7e455db522721c42fcb137b71823d7d3852a6b532c4f0053e648da0a8cf62f5c6b2f0ede085ada33606843837f30283b652c659e6a70773;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbaad285a8a6df0cf5b9f0f9c8bc9633f15600fc01a3e7b7cb99dc5f5210f5d24f0810937315a812a8b1f3d68f4312413a6230ec43daec54f7587f34f5d22870945c7a6cbaefb1f04fbbf7c1fc36d55c83ba3374fca0ce5b5f46b23a11808ac7d391e727936d53a325c2a2f14f14b36e7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0de6b521677aeaa03ac8250bbc3af771e3b662d9536ce363e5d4e907afcf08c43d3e7098b084fc3ff690bd97d039d4a41d90cf99f7177fbe2dc9b4cf6205fd931acc199c7a94ef0641ac6167f68e6668f3b5ceeb1803dadddfbf7bdc60d4ee8482c38b5f46c28dd5915b33f652612966;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32cf877852eaf021dd51e3192dcf9b2c04a4149c4fbbb0dbf8a4fd63a73e8d4f13ea997c931b92add126637d80ce94547e7febc2956e32c0eee66b8f1d5cc7582a4209cb350d5f29054af4879f721024cfeac0eebf68ae142a1039627d9340ccc15eab4cfdf563c4a7b2e1103c82e04ac;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf85aa4ef7ea154cc9a0e0b224c9a867b5f6eed4e730a8c022f609402ec179a829f4efaab85d77203802b990f41a450be16ada97ffdc3ca3a68bc007a56a30a4f83f1bf77861af4a486ac0711ae290880c686b405f3d0c82ec24d04b3cfdeace2a74f1b9c19faad370184bd50d98318939;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc1649994398bda5896913f549fba19524c1903e66bd6a51ce033e1f41474dca50d099f5c5d71d8f54819ff7ef6561921728cac956982f37b06747c4fe1a7b167fcc2c3b43b648194b5d7606c6640279765d4c53df13f9729577e4962522859d314df076f2abe015fd481fa995b1ac15a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e1eb49b6db54b986ae3544c69c6ac75809b86f1c59e09dc4ae927fc898972964442966cf8c62816ae31c87a81c69c0b9134034726911d11ee823f4ed1d3b340a151dbef481f172837fe89168f164bb4ba7e5341f9b0d38cfe8195fbb1dd32b25c0ea9ea61487237ce1a82ce3c3f6fc4e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he76815df7d680c0c359f74f621f320d7cfbe10a2a8384354ffcafd07b0bffed9cb3076b63a28d46fbe115b14f95c2b1c5f7dbd894f72fae255b12950d654e14ff31d290d65dbd63207f1c00ec30e9cce28a12317550e263f2de820818f62763a67f7d43c9171abab36fe578126997cfdc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe0ef0d6cde4881848f8759c92b088f6fad2a3aa37eddec509f5312656af0c8f240f2491f4f107483dc96790470e52983f6926736507c9ca2feced927fa14d21ab176dc62e5b479861b6333afa7998a32df8d35ce5b98b1ad17214f0e193cb5412300c2fd23f7c54eea8ecad560c39a09;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h780f8b92d67c9609f1cbc408b28461cfd02d6ba260fefa4f4126988ba18c7867570a202e7518cdfb1b642cc1c5b31e8060fd1210875ac23a39b3ef47031bc1a088613437ffd909f438db5034d0c8d01fa45b028b0bbc514afebf819282704687f80a9096ed7f6663e92f10e21b295ef67;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he9c12a354c737ec13d75df178a4bc5abdab39e77dd91585015146cf1b3f943567ce66739dd4a75bc8eecf158102e21a3fc142c6b8a25fda5928e4450f7a02dbf3b698fa681f6687b1ab6a7f39a260aaadb9056eed3ba6c12b09226ac65bd1ec6008792000fb1ee99e727fbc4f5c4d3a1e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4271aca7318c96f08c34826c6066cc5b2616ee886bd7fb471cecd8539acd40b7dc940437a1791a0c56d583753301239832a10d30f678b5fd2c79fb1f3fbaf5805ee1093ae50b96eb50bd23a7eff3f1a118d14cfa939fb7cbcc905ea6796a26e46b0406bf27bc5ac97a8f953705888a67;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfea4a4a55e3a3abc278462319fcec3661a8f154b4a4153af827f2ae870e5b1b048d2a149a3a52df3fdf92de951c4501cbd365459a36dc26d69834de0bf24ef3140a24b00e3f14fe8af75d5ae975821b6c5683b96e559f627a40277eed4e85a1f5b21995033e988030a912b9e1c581524;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbe62dec23c618df47ac2da0d87b8ad036a4576f4666b24b8f941f6504e4ec1d73b8728928fbd57153640f3c3b937be902c671d665876cbc84383710ae866e7291c1a18be46f8bf728ea916f3c294b683ca837b7ae8ccd9eb777039f66ed92e85ea460fd738dc50103ccd0f77575cbeca3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc95b7b7850640c0034f761f19b582d55395aac55858d8381e7f60d53e1e41ff4c3c92182c21bba5952f10efbab50fe70add95b76967b68d641415710be84860aba5a88d9d05c37886c3366f7734f2733e20597116753a5a1bcc63340c0f9a0707b18da54d0e67dd7b8405ede9986ad59c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8828aa283c507b5f5da86a73f4961db3c3e1b279023e2e257cf7263f1d7a7a8159935563bfe7834710fe60a982752a9ba905fec25a90f7462e011a46526635badb473be494a9575b7f942fdbe540fec6af0084ae4f0dc11feb87b0332ef81db8b699768606e1f400797aa78c8858000f6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h724ea96143160220db6d29f1943c792fdb9b45de81c855c89000631d6ddc58f27560bd0ee8dcb6ddb7948af1bcf5f5daf23b171347652b7bacca5596cba67e4db9e71e38d67218f185456f09eb2c56883341b7fbdef51caea40801db5d36b7bf2ac435aa8534dec0c65cce45eef1f1f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd42e62277360f04390ea4b286be32f4812eca6861bc43cd7006381961c09162d00e10ff7688486735d69717ee7904790bec2c1e07e9422ab84fc868250cef0bd4ec9bac540d70ecee10b82713a54607e6dc1f40777a2fee58a374fbbf212d954839a23176b1602eea8c1d8ad90b60a5f8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9fdfb78f5dc280e4825494cf952df500cb17da1498ff9d290fec3d97360cb193b6820ed4eca7b5efb0b6e03686186f9c0872c43e7e280b17a2f124fa18b5e4bbb70ffdd23bdf7f8af2e9a864f9d5c7db2d2e122bd48be2148320009fee7f2b007885894e1aa21c3a9206d7a0e8bc8c121;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h467bf419739a9d574de4d5c093cfa91d92fbb5d9b021b73209caf7feeb852a4a5d2e4f38e8c5a5d834d920905ca1aec8cc41d0902c8cfe28a6a6faaa7b5757c45a5fab46fbaf1db74265c1eca160d073ade701c009ce599b80b16f24992327a049c76f3e635ee289a0d5334ad3b6caf58;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h274308253ef8c622052519063a6202f9a537129808387ce9aa53bf1e52f978d1a4113cce7f063190d040caa6ab6ceb73baf045255329f5e5e39cc2b628f97ca61f706a44d4b9ce846fb1bfa698678b4e695287faaa2d63275458989b633413acc890362f11ba073c1f985a80d11117935;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h681416bb5996853f87da373015380a00d731dc99246f07f7055b15b9ca16dd08c7b55cf2265df613f587233b7109d4d6bb1660d788653c59badcb79b663079e6adeb5b2040ce8b7f66acd9fccbfc0e3a0e5ca5bd8130319427b997b7a4bd2839ff06a9c6911e42642a2f231e836079020;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h763beffb1c6d182f85a80c5f6bff0c2012d36ba2440e5fe413aa52a29a6d078d0d661a21b376c627ee84643bca9876e035f05473382a9066d7bcac45e61883cb432cbe652ab5d746e20ceb7f2cf2e109e69157cfa170db5d6e09374239f7cb58bee5e68984d1437f1f2fbfbba21dd773d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h793e211af05c93233509f03d7870226bd3275f7c92934b434011bfaf70e63bd2f4d1b9132d2ba31ada673868d6f7c109630a8f103c963b557a686539be61374785093784750d26851fc8dbdf033802b3528738f9cc2a2f831e0101aa13c57d39b271b1065c6f3c4bc5348ecf4e3a5b290;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbcf40ab58876a50c0fcc28eb78ae5c61a0a26105e640c95103db33579610a18b9437ea56914ba7567754007c1b89f18cc811af0841643212b138108fc087823c4bdc99d6ffd4c4ac98a4289e39b0639691c3cb9a09080481bd205841c3f519a93a7e09129a7d69e723fabb87d1b91c358;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7be0dc70b290e0febf26ab425aa4441e9b730b225d4ea415ee456b0374524fe837dabb844e870f57901ca36e074df517f6c6d3db84fa9da5e9b0c6a7cd6a962e2cc53a37789c3eb5cd792100de16400648c4c9530e13b19494a2dbdd3ce5068e24dc644c1dd96c3eb370195452a2129d8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9bfb567bfd493eb1bea3c27b1eb05254d1943ad5fd66bd59c0c4ed139e7dfcab06fa87bc9e71ae8cd03ce970cac208c49684f0010246d0b77ec7026b4ff9f34fad37860e011b935fb86e34578edd950581894080795475f866bee6390489d98803234248a9ca89d869dfe605ead8dc0d3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h52ccc788b2f432f390d4f5dfa1df0f29e5003aac3d556b1bd59e655a5783e7c5ecefcbd4b1dacc125bc27c90eae4c1b7b182840b5e01feee292b4c3318fda0f025460969c1fdc99df6e05eb46fab9c5deb414919e89b5c623ced95428eda7032afdb3698effcb1f1ff56cd4f35a88f04a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6195d39cc920a4dbb6da814d66f40f690b45d9c833fa9115d851192ab46e1b170f83c0f75e4ffff60e8ca34ddf3c41edf4239da0470484e68f7ca973869f183405474a69e87912c46fb1406fb97f9f5ee145a269ce4de6a854670816af6654670e157123a8c9757554fe66f5b8d85cd7c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hceea88ecbdc3111986264313e5c4cca104134dd8ae723cbc396f03c6d5168cee7c8cc23a3d4859a239c36751b30dfc95ff9a0669f0eee986732c9a046ae48f7facf6faa5b03d24cb9b543fc3c0b032ef25ffff0f63ab0bcf414d245a3f1c1ff6f7c1d13bdd328a5a52dd75736b1741209;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a657d56dd7c3d21d22af80ce212885432352d91026dade81888e078f16de56f95ebcc8a94e419c4b10adc5b60b59f00410141c1d76b06c72c13463a08cb157b95a50c0238034fe4c928cf0cf3dbd6a04ca7d80a335645b04e6eb4177930e269db9bcd9563018ab21d6f9a8bf132c0659;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b4a6965916b1837ef9965afecd1d7e46f6a3d9fed1406745109293830b92810aea3b0c25df50d88e6de15e9cf9a6d4391bd073a00072579c23388ecd7c68d94aeeea9c02367c39aeaae4a422eabc03e28d8cfcf127968022030ff40925bec773f65dfcae1945f4bbdf07959801a119f2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c6ffb7a8a69d694ee1a6e70e947eed92d57794962305fd7690332aee4c92fd7b911544705d8a41a59de3626d2d097aa5408fce70402ec9c28cf626b6e9e812ba5d1268851304f260dfa74e2dbb7e71a8c8b5402dea81ee2a0277a9c40cf3654a7074b29f19ca506eafcdc2f05801c746;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee884ce704c855a63920ce28a6a8fcb04d1b495a5b440ac6a6f747cb1aa0d59ef3db81c3d95683a9dfc67eb0f5c5d0366489ba58b267463625493c0b8b7f8d09414d5983955f6dc90dcb2ad3d73c00179fe43be5917040a659ac009363eeb22d25a6029b75499ff48acceef751212d168;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0680ef3452f97b6313d94d7685b6b3eecea05bbb61fcf3776b6fc866406a77aa2cefee55cad2bb064df111fb24a7831f9064369a90cc22eb9b160d2f831bcbdda62145a417979158ee5b8f92aa379ad25830a8ad9c2106c2e8bb6adef921d87f6a49eb8d6479f71f341f3cea6600d4bf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c23b0f610b010b8e65de4bdf23f3bcf0c329a4fcf36524360a95969982748cf2df8fec0f6b2dbb3433959c0a96138ea6a4c26235a9a030c69952054eecc5a4f3824a18e2358f0b0bb36b224c2d713c77208b216a0e205a4d2fbfb91ca8e138c5118df9f08c89a977e3d1efe36bada0ef;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a023292cb2cf804113a146a1cf73c18ebde1ad7e5c486d12d60aafb3bbfa59323cdc56869bed9eea7244dce504747ba967edbc74add5d2983ad7a7ce7e80c489bde79e87db570d8bb6b9c69c7dffdbb909da8e5aa72f266668668e182322b6fbcedbe35435218ca775b80b820d61b3e2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc922d69b40e56085e5c340c525f174390f50acf6c35d7daa0b7243351d45239cde8dbdd4e04a08c8fbc13bdb23eb07b2941ecb453750a2a62c5a165e8c656efc90d9f51cd45abda16703c9a634bbc2659f469cd59af21a24cfd3f2f7dbe3bce984114ec12a0a4e630b2ae2fd50517bdd7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h658f22fa5d20b16c8239898294de7504543973ce81d1c15011e2ce791981ce4fafd0876c5b9987fedea331c58ed8ddef9542207e5da83120cb8c58b20e6b469225f6997ae7ce83565fe07cfe4670dedfb40c39d7694953681a12558ee9b9622a3a978a76288058994ccc3952f4fcaeecc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h121c1f81f3dc8a2020ab0a6995ffbac69f03750b80881d4e5f0e7070e25f6e8aab752dca8abb764f82df5666dd7d768c0a2d6ff83d1e8a78a74f0445563fcce234f880e87de7e689ced7fe58ed652ded6df36b4495006d0fa07f2aabda7eb96f04b15404a98437eb6b73701335d94c1a3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h751c1c5038dd61e1eb067650c534269c674c54dd366328fbb1db2e1a18bf15b095ca6f95df336e811b4044b508ba3be482584e76dff408fedbf3a29fc9d25aa416a40f1a2159c08eda3c2d11067261f4203359565b9dd6e72970f9f19520776341b57c119603a66e9eb94cedf4098ff12;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h777ee797b57aba75a46a821fda671b8060cd5b9fc4ddc0a4075edd85b2e9a72d0b4e1f7ca837db73f01dcb826d4c8c4fe36d48db9be02b0162184ab351dd47dfb87548ef3f23ec48c722329455325d1d8b69a997a7d942b7f8b6394643e1ac0a511695e4bb5cceed3b44c66654acfac29;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d701d589b1661681fb57f29512843e810c20d5c62cfa6285d1bd4641ba5f4de2243a8b09d29084936f3135fb688a9fb292354c932bb2638940647c69fe6c07f1be429827a27f4de0c54c0dacd18081dfcb368586f58da9f95b245a0224186c87a7722bb6fef566fb8db07a65062f3adc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64abf83a9a91243b68bd6fe2a3dbc62aed1cb9bbbb71ae70a9a5b1531f524056d0ff48578665574ef01137d42955735254d995fd07e625f54000876f526747d0330c60b05507b177a0f906ec900d3b5ecb9784b5544d4a01626797c19f616b39e99252f6158cdcebf3cb6015b54e0b957;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65c5fce50fbff34f1f950c25f352af880869eeeb1aad98fdd811aa986fc1b0a2baff8459834194134246f13e7d0cd1fcf0bd1e118dee1e2955d27a8326e17663577ea434fcf9d5ddb94ac2dc5fe5379fddec3ceabe1c8cdaac091da93424cf4148627d2dc78688a276a484a78bf7bb073;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5db2130488b59ee1203fe5ba118256ea2259b8f135c941436e49e68ebda50842a0a6141b492c8c8d58fd42fece39e83b443997e12bcac6563a88f88a3d53d28c8b7b1bc9d2f48b89f3ebd016056132f0a77003ed3de32cf12ec27b72be3a1ad75c0641c8ae4026d8ad0f9bd2277af3891;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc6a27a5a51a6c16558d8433a9ba904f5986a83a9822de9d2c616a1a88ee45c79ab7b7ea5f33168a34c75e382a8a2528f121f3cc09edfca3d16a7849919e1b1b7583222d9b2facb4d04f2e788cc592115f93040f0b468bf262f266d16a4324e75989d9fbb6c8a0ce6812716cbe61e2a816;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58bc562f3d5b0bfea90682e86cd6be4165a539db7439959d8ab6a0b0982a3d9f81fe43af2879d5711592817630774da5de63e3437c08171fcf1dc3d83508ba307f5a6180a4ec4ac7df4620dd747ef0c740653397a28c6d51eebd02f4532728f0e02ecd023b74bd25c1190bc050dae5f71;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2c4bf2747955798452e2d55569b6587f6c70dee0d6ec5d305fc8a20bd7f7312276f9cbe77843c49455e99a468d3b4acdde9e801a4759044e382c16b064196dc1ff95b1a1043351414acd5e63d0e3f54a1dcbc817ac19d9a6e24cc62c7eebea7b0f61db5cb9bb1e8788c179e199862c7c4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb73a51def2f8afb12d93fdee09eb07168ef39d283da5e84a5128976b0c0c17b71e18332c928056cec92abaa434664a0e8d9af74f9e14ce44787c29da3c0899a5fab9f9f32ec52b982507988124a0ed22e1b3f4a4b108806ccc83d0847ee969c28bb19f93b843bccd4d8526063ce98107;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9dbc78acba4ae8e8d53ae87447cbfe73a9c3224201ab3257b5f96317983dd8f973c7dec891284ea3cf73ab4350d36adc85928f543af7712cba462dbf33db9e09e8d174232a875673a6a7a482f9bbeedfcdeb077736d0fdc0040a91a92cfed1c58b6ae4c9687a511a363d52cb5f2996ae;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb2a9825eefeb8899f20f6d14e284285338ce41bd8e6c10d2b5ca65e94afa32de17b1546a281a4acd093e627c1fd748f07117ba41b08806182d1cb612b4d7969fd8e6277d294c5f0e44eb417c090ef498b463c412b6db25d7e13ec86463fdfd1a27437d44c0dc9c61c6cf89d373f3d4b8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3f07621a00e03a18efa1003ab55722ec7a96407f3463e1bec7809ffe88065a92447df10092484da157ec8c592edb2745833f5554c97e2cd053c6dec96dd68d95e7bacdd072b4b4896045891e01dd23166f78a97ef9dd850a5d0b7c1a0ba41e41bf72f5ea4220c9934f6e2bec93657ba8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2785ea7c2d75d6e84f04417655914c4b9fb082852d8798901e9fe7f85683fa55b253fb1b3bbe79c52b497793d1210b0e8bfcb3390349209440fda1c1c13c6ab618957988a5b34d779f33dd9f1c6a5396a0909dd507d3cdfaafa27d3943f8e54ae7168a1c9443dcdce619ee869f703b031;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h67e2a4cbb1437510f1fa20010724314ec07deb3ac8447e9ad759c992b858ca1200cc884c45c3c16652122f778206d21bb405d458ee9d78bde3b94eb8b913551372a49dd59d269e11110d622cad4ef5564d8023eba7c2f7f4b19a31aaaa94ab97b8aaaf95bd21a6ead58dbc1f5a473cc40;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9b9b65592ca88f267bf89792ad31dd3bd679e7d1686482bd32c1f714e997c87b9adfe1422332e21202483e86d7ac1a7656442f21730e96c3cce73fb1e152f5011f384e404f72669086689c0bcb939f5308f90ffd30ea5345a2b5bce94014ff458ff87f71d689b06e497402c2e97c7276;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd09620d6d036630f9e075b85242485be906415db291dcef0075a8aa856d2c6621043c643ad2b85b24d8278fe98f00f0b3279e29d0af94611f7b1e5b8516ce52ed555a304f9a803bb12777b9b1f5f689da21fd7459b41407c20efd3165dff342d577c97bfc1b9a050e9689c1e0a783985;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ef07a9b02654877ee1217216a9cd465fbb7f83f1a32b6faa1713d3c2495d17696f6921118acfa7bc4d1569a5bc37dcffcc98afd7c836f775a6bd1d548a0934b83fef42d59f37f9e64d7750bb4ff3859a075e0a7d7c9f82cc4b39334cdc555a8c7b9672845e08098da5ea087207dd7ba6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d163e5ac7890f484d7a1a7d472ad8fe7e60834d62d07960980e686c592112940caa6b738de05fa36c791fb5097b90fae8f6c4ec85e9ed9bc577c6ff9a607d5e1d71de5b66ebc5bc3ce4ad3bcc4f625ddc3cbd025ecef6ce55e76431e6dbfee8c6ba9cf5e578198721d94725d8e0bf065;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ddeca809461b2e4cfd93cfca71c6b1468a8e1705ae5d8a3ffb5401fa100c782bb3e7473da2d19134a6deb17cf81607ebbcac93f2a16bea41ec56cd9f4c5e733375152ebb81bf8ef292d40eca02cde9e52e24f08f7ad9ba0c249cfcbca8acc6344ef46589d91f5793d261a06257812874;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d3d4877ed97ef0ffc301a23913a8fa38e9ff49180b89f266453e1744ba7aecc88b7b05f1b292fe7cabb65cf719759ae5dfa3ce4c8cfd4dd86e894689215df0fdaefd980014c784553d3af2b6397c486ccc9ede41e36831cd6af7fd51a232b40bb08cb28506958349ca2ac17748f37437;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7334657c1808db04e10b8da260c26df293320b92e7469f96635691b9518c865445b09e58ddf38414c41de28fa16b80b12352158800f534ecdd67c296222cb833651dd3b111509db5d0aac50a99bae9cf6eef56ed6e2fea5f42941bacd053cbaa107f33a10cc3b7646c280713bb128cd9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he625afb24af3d8242b5b099c34c251f7f531ad559642ff9ff1a075e0e4b59d2561b9a27513f80d0bb0484e53efc20e069b4511e1099bd23b31bf375a1b1edd01d8f63afcd12cc1cee7c5555bc3e6b191c6c4e2d655414bebcd5f13872cb165d511ea593f9e951744a71815dbac9cc41e3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2c31f7d14ff7d45657518f9194e66b79861b54436d6d4bd254cfde647a2f2633bfa1a2fbb4c74d2c298878ab6b99b712d3753c6220085d746ce6f628d6b4ecea8101b41b6236e8f769cbf59c98f32e2f3b8f3042aa0ba6a5aefceacd50e3c4eaf9b3b7835b670624387e6e90745a3ba7b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce99bff007ef18edd3878379daf132375475cb033a799bbb3189a2aadcaa04fa5612e9376233b9cfc8c2b04050564c481eb609d93a913a625b6259e2ddfaa5736bbffae4b6b9880a186e15823d253c62b11d09903ff74a59126ed8b2cf70510b376cff12e64b530756ab31f4feb8ee031;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9843d94434bbbf01e274776c732583573eee0cc4a9bb7d632f4d0b6fb05fb98e9612630e2b4f66660e55107b68f5d5f5361c9a06a07a59f0f799855cbd643fc01f58b03621de45316b9f59839c497b3d3a82c99d615330c2b809b9251d9b633e93d8fc7285de7b110661a85b78b9fd6bf;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h67c2a41a833b0cbc806006a0676fc37f9a5699021a22a72f124d2bec4f04fdb5d772cd7fcb91f7b7497cfb5ec90402a56fb8d18275650340a71244b7721f5941d5c702ad5415904f99c5ca8403b92c0c1d27ba5d064ee8a099ba57af4ea14db77a2895e34ed521fa2329716399fdd1219;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h77e3c128b13da053ba684dc3e916ad32374576425c05163dfda8383376bc006544c356196f3e9ebdd77577f159656c8e71a7f64fb8f5e341c635d45551a24eb3c8757f294787c65a185a5a582cedcbaeb5d31842c8170f2343aeb49047f5db400d1c7262b669181dedc3ddf8051de8fc8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5748068ec4cbebacd1505a3d3a758fd89b1ebbbb4348f2cea25747311209e0c3bfc1b75e16a854811a73d5e64d9ec1a55d23cdd6693f9e5cb385126dd3815d84600c36f4520ad8590b12471d14f54f5b921cbed9e8f58ebd49ac989bc5771fa1e55374abe49a04622fa6ebdde1e035d1d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h33a6ac79e20d48a8c59d8ad25a38ad8d67869a467258e0ae25063b8837f3d7ca6d41d4a244f12bd76015ba74166378a5af8baad6f3531c56ce879ebf06d812766a458dcdc3ba16faba5236711db740a26c27df8f320f41eabd44f1716b48e6dbec964ab53294bc69562217365c74b9d31;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1580590f9f2d76b269a8ec19a5f3293d86cfad1b71d93da714d2e1ae5a2cdcb701fe5ace27dc96c800438ce5b2b41ea6267a1d8cfd81989f8a9719363ff8c0e551aa7a8700467cc1911d116c7dd6fec9e8879ad5942bd8824b834a8210424ad7b96503c571dfeca47b0c41a6f8a2ca294;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5fa419c15b10195394c6b27fd661258120b99f34e951dccd148f14f832fbb000ac75da245eaffd6c25ad693eb1f11803b81cb29f1f4fcf0d0af24f028516fa475cc2862f9ebd579d74ba58c615170dc758cf044ec4508c608ad2525b06f8a1910080c6f61b4d3390a27a6caebda70edf0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h965859140ab400ff3bb162272ef790a65457c05239bf52c29915d3e369ad827239965ef3d349a74ab3c499aa98f48b195f8440e8136f0e73d9b5b3c54691cb09516acc0e67ebabe8efbd52adb9c6f2aae876818f4aaced1129f9f71ff6a6ad0497595c05a0275b80329d3480719eb2abd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6e519ae02b4f811b229e438bb646893e3b41a1032e624d4b94facb8f26d54bd04b9f40e225617261c7b3424e52a8f3e0292a87a8ea52b68c959d382221b7ffade15d429ce92a3c1ff9322becb97ff3baf1e1de245eef5d05232b97c1bf0b62ff741d8cbef4cff67347c079e2aa32c9a0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ac8186b95065eba72a1c605bac04bed478cbba901f43406c031199c499975e98a50402d6a0ec1dc41fc174aa39ead67fd048469255cfefa728c729cb38bc8cc5a45cedd524ec66805aea9d3131ea9c3f2640835b550fb7cc62b2704c3f6cd8d2d698b4f78a183371747839d4a4f04dce;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ad9c6f178a75405f07bc5de768272522fffa39fb5b737ef3b722463b2fe04e761b98c8df7550f4e63776ed0fe7de85cf5d5182c002ea8453eca7438a176f37361575cbdad44f624c604e4895c8e56534ea3f4d6464be829bcf92a54577fc552eaeb66904a0ba281816b543520520a44d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d35eeb41ac8de78771686b520571cdb8e38c69b33545c276c50de79b6351565d9d19e88353df7e55d8b4ff316b3f34f5862dbdd9b354a78141cfec4dc2d803fe5c2fbf6fb6f0501ffcdb124822d007dbfb4a7fd370c19a4d3b13ca723611920d327f674ed8dc03e60dca55aabec4f2a2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h15509eea81056196903773057cfe12892981bf6b7cbd54ed4ed779fe5f08383ba9f6ac60a40839dbfbd59041c617d0b9252c7dd3e374607cdabd55c197d051c58127eaf7d99253252d283c0b7be4f56df0cd63e88c07768486f38772c2dbde38b373d5e2f057eb195338ea37d7e660c67;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74e68ba614d8c8eded7fe467c259b359583a5e2516d664b6ee8fe8f97f1d60cf815e0e399ccef9c9ee4095522341a6548fa7bb3bd14427d3d97fd766e9832682445352e02f7edd275bf19bec46f8661d1b45bcfa08bccfaca373daf6f177c3c98043070a4f31bdca0e221b997f1de9796;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b2843041f0b560b2a15cf1cdbfb4479a81d4930e38097f0f0abac22144af24bce4791093f493c35b2ca1725889fbf525ee27a9e30e038d9935a479cf05d68d54eefb065b854315150d1ea6c380989aa365c4f56d9803f5e0da8613cdf3d92f8df8f0a609df2c3e27ae08b637bd2cccd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5362a2ab8b45dfd068cdf88923d97d683f129c717a0eaa475996d3fd74a8d245940a0943f99909db63dbbbbdca8daa6d3522eb647de0d45fd4298cfe50756bb33714d4e2d7ebd85bb51585ecc13eeb4218cb677c3b2390c83d129b95af0b58d5b6fcc89291d1ef7e91a63ae65401505c2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd3df23a83c9a65493fb94dfdfa73c6cefdeefd258d934a78982c6a07b086ca5439dac60c18955aa3510fb809b7759e4f5abadcc2c748e319197d306f6be8b6d18b2f11ab7bd51490d895becb004fbfa794fdecd10ca0c8ec0d7cac15aad35cfefedbbb1a6f20f0f3a51d3d80251d908cc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75c3ae282cae6dc77bd50b1f8ec51cfa1431bacb4f6e68806d34d02e734aa81789045e071f18ed01b004046d9424fe03d573e71054df313bf7272da248fc57203e1bb189ecd2c74273fad0c9fb98bc735f4f089579c977f1ecc169b0a0e583d06bce15385f0611565579216e06e40e589;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h554f2b9c85eeeb9efdd8ca8dd2cd5cc2474a8844120b4a36b258969e982f97df6142589b89d5fc0e17ab6429f63805aeb5c621e6ab78705b1e83b59dc43f7e272e69f7d9895328aef888305e266d9f04034d583b9d09c274e232fe04b3678f566637732fc8db532cefa71f93241a64b34;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8951ccb2eab37f3c9407787d81c3159fe02a5b2f9dde943983b28b6b933e9997483abeed62d000643079c6c6ddc07e40521fb8438ddb890c00cbf01d148440c04666e1cbbbfe7befff9907f9fc5c6670c5532000e68186b55cd5530acc495182cc25ecce6ca04c60b575680c063da9609;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0dc4f6f30548f1a5b84ab52fe9db293298d4c044600e8393718daf58c25482fc23a49b19cdca57df04a8d144f42c0e1bb83dc313bb541a442d69a5177ebaa3aa84bf931bad7da15f77b8a1c964e1a64f46d2f83c21a9bad608f07d5e9e0ce51175152e8fd6864d37b3dd4f3ab98aa7e5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd7dc73158ec929bad4983cf72214eda6a80b141afe267514c97827dae6d7ab439f1645c3431b8f1f45b71649b76ac9b14cc1819215755e8d92c335282beb0bc1884069f3829d8d3191c03b6948649b8e2267b549dc9bed6696ca448c9a818556ffcf221c9dc7f7f3904e36361e6ba0ee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7615b0e086d3322ede3d3115ec2631f9fe40ee9a6f37824faac8c884a6a69cd849b2d3b7e0a0129836e2f84a2f3eae724a644a9b7b66aca155af6e330a1572739a261d4da930e67121c7039b6a7bbfb0bfcecd825d6a28db98ce70e3de8b8e5e2ef73cc3327281485256ff533bf175f47;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72a289f0bb1a71128c67f8c22daddb9c936667fe536e614a234147dae20571e4dbfb24405443ac6e8e7be78e61230d7fcfe267c02af12ed880c232b310ede18cda6d01667c9ebfbaadfaffadb6a61543bdb5ff7d344a37d72ae68eb3ef5a146d0c4b6de8338022baef9dc0db2e945959a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91059fe60a3fd72e4833fbc6382ab66e6c24f54364016b2b6ce21e55beec7a7751e0dceb96d799d6c6b89d5e2640ce5344e2df17b477b7e68e81aa649626fff969f206dc242ade2a088156926eb9ce0575d062a668fde78983d5180d6ae9dbe356bf9a81b96ec15b7dd5a9ad9f819dbc9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2af40727ee41813940111df35c770f900418187d08db7deaf432c8376445e23e0fe560604259f9913421b6430e5bc54420295cf0d03776ce00cee96c6714920d1d56534133e0ec23e4f1285b67d58b29eb541d6d7c6c10c5881dc2b7a540f9f0d224f5d4ea980cab243ed7c89883a9828;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f5b507d1ade0f9b253e311e7e95b1d4a53bf23c25b34a0365ce51eeaeee305d65bd8750b63b772676fb576ae578d177a6e84d6446aaf5abadab71bbb2da406362d420a3a27f2b5c7d4ecb8243ece8546cc43d0d7efdab7519983b7540851a2a2bd332199ca8fcbe6b8fbd7371a68c93d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc29f3332184bf353564806eebc760cd9f420fe5b8072e4e1be44149a3f9c678207369dcf30ad161c092a94e59d2f1288d5a480baf85744273c56723d35762df5dde6c189c1904ebb6f639d67b18c8a7ba3fefe2128cd992f9136837c36b9993c5c832019fe4533543dcdede53162356bc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb72eff720691d4fdefbe4f5f6b516fc037326f30695a1b08f632e6484fd355b33ad3fc09eca83a92e6265553ed6d0ef4470d88fc2a3d0dcd95eb0dc3876aeaa65dbb74ad266c6b6057c7dcd2100910e5d1dc8dc175f5d0f32da613cde5a92bb4a62ea8a60c0cd82e0dda411528000ef37;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11b34a9de76aacd7de0325a7592bb220388eb900e2432923d9dc15e0c1f3553ce6fc22e86c2cd7f449b19344d8ff818b318e3161e6677e0d2f730efb6cb5d79f4a3cc7f4c5aba1f647f863810e1e1f012716bbf436640ab9399caaeb2b9899b85326534cfc6dd98ca43a69dea4518c092;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9050afb17d88fea4f887aacb4448d8399b67e40c4869c481b5bc9a4cfba526b0b140238dd641002ec587eb8d272f416dd9a3683ad2834c5a8ed7d6ce2ebfe13b20b7a2f53ab575268b282bd54d5a085d16ff1b0cd839b6a0ab94c70698180d5ee2b6ee2765b9b9c3266d095e307b52e9d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7b5c997122a7b1cc6da28b831786376df96fe891a824453e6a1905ea80e51ed029ba45a9009526d5eb314486803aab9525f6a3a6ddf13f1fe0ffb473d451286fa1cffaba83d464eecea9d8727f89302d8b8e6126cb7705700717179f66b4d45b538362b3dd63cb822bcf12127ac5bf59b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3f72028418835fde09984d8a817f426047d613cb154a551235d9c363575fca194b623b59c27d837e518318dbc3e41ddc19e65de0c3cdf63c35b9d8a45d331176210699644f64f6a5d256a71ed5d7cc1ebe632041bdfac097d8d21b22a866e30b16b6009480c37fc146b72657b98ea1779;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h16600e321731b2b3aebcbb29dc7171ec67ee5bcfb38c479e987ea3ed5d103b7869daa58e1f1ef56ee745b51eda078c641eb7aeab7c694925ca0254412c79322f99019092ec41aa3075961fc27a64491d1e3bf61c9fdcab2672af930666a30ef636f5198f1c8bd71d293d457735cf1064e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8b9e0ceca80d99868a0dfe88300cdee750bbb61122da2d7a4832ef2f88f54d87464eb74b387575c1c7ba4f2363e5f049d48cc4e09d0de373906c3ba642459204e08232a4a74daa0de15f453fdb7b9635eb44ff93f65f6eb687e7f9c168036579fa8323f0a21cc90c6d9df6b2ff8238f4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31794d261b8551957a92c376f29e5b6e5b9fc5f269728418692a0342f7aae21fc3db0a148a14fb337583b4dddaf82de65f7cb70dc7722aa7ad6881ff5dfe5ee414575627fb1ae3d41659473ede35c7429357f3e752cb805a5a7e7391ba3530551bee5756c9e9a91a26b1dae745e4340d5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b7c81a0072191e7cd4e4607a008ce066ec1bd793f08d3b62836d7e2348da7e737c5ee79d41610d3d927ec5c1cdc15e858ea23766f888fd079d50d6d6c6122dd43aa620f746e9b95d74d002a52001518b4aca9e42b27bc1b62596c277e3c9be962aabff14953e9811bb39fc9ad791f467;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1ec8b3275c369284026f4e4429c8f314a9beac6c0574cb38d976af15f671e99d75bf4fa0ea533587a03902dfd48b4cafdfdf998324269218dff91e557b76ad987bc68669833bd2d5dd216447650afd449b5722a392142d6e7be461f9371fafbec53d95c7ad293fb9416cf3e66f4a2e83;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfaba5cd5c953d6d33f00da90d02d654fbd5c3b7b975a03674b54d24be78df3d3390d183e5817aecf83d9be2953964272ec459f17808abb2333a54f62e0a5ece35fd10add5e2ccc6e8857c3e027bb3ea2d19eedfaf4ecced1c1e48d7f9beb26a98f603827d09cfbc283951aab53a0de040;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc6e23f6151f44beb7de21dfd5e84ce4880d22b1ee216d0da9855c80642b5eb0118269776459106ab21f598dc5a84414b82bc05f0fbd0d9dbf4d131c308d1ccb56a9cbc1f7e37f2db351bdf08f88922cf64d43960bbe38a29e36656bf1c63a1b962510de72d698fb4e6947ffa83fc82bfd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7692997f14fb337faef50788c1e6f909cf30c07577352b7bed0f140dcfde8d5a9eaf5a2f1a2446bd9481ba5cb1c523fd45e35ab73b2c54b8c37d45beb1134eff9de07c8a25af1d83aca380ad9b9f98685717ff5e4f177f0357785583dd10faac2b309b3e74e35f6831641882d95753c5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd191ec71260c44cebfe15892ea846cb5cc6ee48a60c5471030d8f6d7052def6c73e7b2ea6cd1d87c3b78967f7c531227513717eb5d26725ca84f9a2ab12651174fdf383823e8fc749af99329cb3d84e9f9794bbc54a53c52ebabfd991f81e2299be73bcdbae6cbd769300a2f1c164d28;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a514fe18c5d455b97274c4b93bf60bffd22d98ee6efa2445501dade74e90a7099fd874fed3b72bfb4e4e12a3dcb85a1bc4ebcf3fa5336912d439ab76f48ecc3665f36c4fedca4913a0f8526b79e8a1980ab240aaf3f1a6e4572a50069a54d0edea7545ba910de8eec8904ae8ea91b292;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29201c5ae0e9e17915af9667bbc4a04b5dabb0e501cad9ad44800502ef89a9ef4807375e63bbd26390696ba46cc25a9d08cb1aee5317305f066749dcea56b9c6828ce72a2cb9c9257c8a369848cdc7e3293b6815c20617c27c2e6a61a5dd914fe6adb8edb0bd3954389630bc031c141b6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd490e6e0e81d867fc86542baa9adda1120719d8bfe72ed234e5d150023d5e68c69238b8c6f6ac3d27ee64942ad74a0b4812f94969deb43ba0cd351721b6b4603fda38009e0a3606af8885416175e03ea0c346812061ba1e61962be76503c72eae6c95f653aa44ec76853ae3bfebb2e5a2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f1fc01a0dc8587da9845122aa60923ba26a3d24c22c442dc4a132099d054caecdbed4f7ab33a08f530708280eaeb4ff6a71c41f3db0f91a5485eb0619027c90798b5091774a5f73716c59dcee41988e73b6dc71b770886945a5d2f635f5f1c811d148cb09b266ddfdb8aa9aadabe5405;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb181ed34715eeba82e07254e5cd76fc50bd608c7333491fab696a417e132f50d160f3fe27cf33ab09bf8c34b757faff100e06fa73e9afffe45c476c972d244c632da61832dd35a630fa547587d2b5c8782da3551010e626757c6081fd719522a9e1311ad8c40d68812df51984f49d1543;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1be542abd6e4238d481196a9c10f1b4871ca39b406ead5661e6661f6ace1a3af435bb6e036beb34eeedbc47787646dbd466c25a7164ef24c83be1c4f125e9b1c7e55925852e83331aad936f360c44b5345735d8a3b110324fa32b5ee41fc991a6ab3878589155e6cfe12f41e2d3d3af29;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd44a81e97a28ff3fe00e32f7133b7f199841b1e1520173bd40534c942c280dfda15afb0b36856f3c250f0ae36312ab22e41b55a6aa5f1c4876bc9df3d683efad6b6adf0d4710a7a82ec0c24cbc4002a976519d0bbdf4ac2f68c5753be85ccaaf0bc572a281bfbd69c087bf2bba67270;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hddb68cdb2b45cfd99f10eee031621f986e86e4b64f64fabfe4d3798643e6973325e91c0f46cd5add6503fa8074c5f44c519697eb277fbb35e43b750899b9642b994707c2e47ef85ac1776a2736a608dc035638f968f598730e0214e3b643b5b07931c926cbd8da122e12d99f35512a5be;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f904d7021fc7e3a731b0179443cec02dce508fad38c9f88889fab0ac0bc692b162b209c3213480d4fba7811fd45d3e5ac8a1ab1a05c0f199d4c8cbc1c816ddc1aeb0b213606aea125a8c0bb9c9ce9c504cf48b223c30fb6b8491a49bdd48459f8059fa54d2d67b147f338073e0e31cfc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e077b9796cf448e97e9b97a121907383593c088fe1eb0ebb731789ec45bc8c74f744f31789a77a444e587847852058cf74ba6fa9f50e6de947bae26d8b2e92e1c15d24b89f8b7f8a509d10bc0436d070cf882cae6489413deed3e8a2668f71d11b9b138f9955686eb06dfbf40c70bf73;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h971b718a528978e847709a582ac53b48ae07629df101b6997a38946d43f0b4e079010b340879d47d039b1e6f5088d0f4f77210263d9b0f6ff6266e1ca9a442fcc4e2c27c937453c37dfefe2ef21ed232accd5ccbcc495ddf0188ae9f4a1ff25fcef9620b0cc2a87f5e35325531fff9bee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff60a9477bd6e63161309dc02495629f13e31640707d642431b139d5568e90944f79e6dcb4a8199b9e08ba0f9e6aabb9defac074c1c0702f82d9f061b424cfd0589fcaf9d45199092ecfe848e938d9ca2e2946fc28a2dcd0ec78180de1580d229c7489eb9eb4519e662bb5fb84744eca2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95f8f5514ae5e1bb021216dd799a7cd545a220d4b67b350301d766f37f10c0891409df1aab354b30e2e54da7c5118ebf0c49d44f0c795a48670d07c0422dd9e202cd4876b5bb3c635a6e0fa6d0be7df6027185bf4b965a56af81d5777a118db1bd7cb2a33499d69997c99489ca886b4f6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24af3ca39a0a51a3833988bc2ea332c5b9be5e2f71eb8e75202d9d55dd64179c6efba3a05a6a03e0795be83e09d5d6d9ffb489983e6a12209a730423bedd84e34e0523820d95e78c393aca441ac8b9187f5694b9f9f0e1bc119124cc00aec83958fa7d05cabd5ec2b7e39847801dc4b5e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbba5d9189646ecbd7c266d3d72a45bb8986a61743f871b0014dd97afaff98d4a8c3096cbc048f72e6f0e19c398f7b928285185106bb269a49a16d33e6b976eb4a69e218cf1a0c048136463783ded1efa1f8dab1ab0a411669a2b87940eefa26c3a4dbff2a6c8287c696bb5e7d1d8bac2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d4f77c33e258379390ebf848ecf78350a6773595482309893eb7411829a6ae4e90a8445665087765d68dfd49b2efd005c0ff22ac7b8a38010cdcc02dca9f807ed9ee11bf79a09ee6b52562e15216d03dcd902055d247b6da5a569e700cd946c87bcda4fc2a321953837c9a7b9384333f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha800d10d98d601220959b5d50bcdd7cf30fe22c72ed45a51298c8bc0b6c7c3480b67724dbedaacb6c3ac790563a3a33ea6b9b7ea64f0486affb75845bc4f211d8308efc1dc96f3f2f1cc69dbac314751a325c9854aee89666135fda97fae5c23b314b7ec24285f1b87e2ac99055e6dfe4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3cc0aa0c2e0404ec51985eaaa64751b205f04172815e0afafcadb6ad9ad4a83b3a47f8d5fb0b3e341f7d6048b5837062bf7fb50756adc83f2160daecbe001a42fb62c64ff9bc7ab9cdf2effe5c6f8631c0d6083e6b77c4979421df09ea8397d69aa0e984d3e3ff4a99aa7831578df54ca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f14053408b4eed92b374b106bfd08831f32c61b7afe3297e5902bf4bbe87a2c3e760fa4d702ac4983adfb1ad66cd6268b08b375e53c6e3f23b618110854f974f69ebaf526e5a4612acb2dd4e1c79d4edeabc58fb090171b5cc989ac6029c51e8ac85c74f00d6aac89946ffe6e69ac0fc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73ff963c75e8e729f4cd6b3f3e199c2c040777f4bb0df41caab71d07e194240c41623584cb763f5e70d819f99f8bc5901b221e89b3f40aae0d69f016a5a16c96d843dabd661e3c259fc1e8e912d3dc3efdb2190bfc9b3a57af2eeb4762ae330326c5246a319f812df8251c2c83cb27498;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ba37dbf1a2b643fdfc875e394f88ae1cdaa3fcf05150faec8119b1df865e927ad554802795ceb185e2588f2abea4bb1e3ce94a3dc26977e63135b23dca936555439a5c49a04f8e2882398ee3ca1e395bc9a063112c5853a571c30a7bc164d923f8d12f37e14eb8919256d759657f3662;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27f305df7ea3a46389e29a7421e461febbec1121a27a12d5f2e63b60ce514eda4c3cda9481307924a9f3bb2bf3621f734c5debb2e79dfdb65e68af2a2844a8ae3d4a7523df6269d3a4742a7ae8f4e6390741978cd900748a7b8cfac1f5d83f2ea9b88ad9af7b126414380ab5078946c0d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81534d43ababfd36b452f60a13fc5e9412875b770a77a79f9468500ec8e4786f94ce1b7b991c4789d450b9077835f19157085fb875a5c08fa1921e2fd210cad898e34d128c06afaa79b3a0fa9793b54200d641a78ea8344530c41d68b4b91890b455723573a1e1ffaa7cbcd48f2beca4d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7817bc0d44c809f5f13b745459462bc60e429f0050e2350ff9110d97ebd8e4a674976692280025d190d228e22fda0399371b2d3f34ca305d6b0d78dcefb3e03d0eabe186b951d393091fee0d5d584393c212943b838053a9c7b131ec0f939525e3ffbc819466c335e98d6633cbbb49ba4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd47c720bfc8743c47fb10edd2d8412e396164cd0864f61e11e110afbfdd8367f8726cf333a54938cf3b78da9db0b9114c4d87140d5a6e7f9481238c4a70df6b55d0716835492fa420f48276807dac06b98fe7e60bcd5cfb9d6ce991de3cd36d2a0c9ac8b3caca538b323207f89175493a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5050bcda2dfc2d272be26e4f0153d0f1799a794cb688f68358ae3210a662b526eee246e52e75d5ccbb0ea39ca949b24d886057acc6a04f5edb0e1bb6a02bf03d2506b88af0ba3e3b5fa79feca0aadf835e6386455defcd81df669bffce9bdf663a6596f842ed57aadadb4fbc79f5a5c1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45e78d160c93cda9fe4fc74103991ab4363ac5113b605add8281ae8005d4cd45ead3444f44b08b339199691a4e7863f181cc2a7afad78a1aa36e364a38dbe7b7d353eefbb952949d7b9bbe4e806d3e51bd8afd59c1a0d61168d024d8666a71955f5c8c879a117bfdd52333f987e528a1b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he763ae5dc8df2b87cdf5b97b54132c35d7660f812128fb5be5a425cc7d177bd1ebdf7d971866a1f645d5b20c8a2feb2b5e64ecceb73a6c9b7febd91d01d0d1131bf752e6a6fd8fa7162024f1821efdd11977d4f5f31ea127c88fc8807b1196a1f028b885e9e746ea8513fec017bd75a3a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc53f822f4db9a9223d9bb558d3e03aaab38b6ad744d6ee77c76ac099081558a8506aab816112b124cfd1665670eb644dbc01d33910e2f2e6409480328426a1b9d7652b8f0430ca2cbb315f367d951004c13ed82e4cafb52a4f52260d30c661cf2fefa2f4fd8058285699b508e70f0e51c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf3138d2f622576ea9a692a0fa7cd49f5a1b1502fc830746d268d8811b0ec018a195ce15ef8cbe0ebe2f7a2d9c0e1e6467162234d4b089d64b3663aaf34d83c728c11aded0c0cf6d6833179fc019a22605df378d731022f3a289a12d72fc36d6e566b129b69e3037f7773d38035eddf5f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he124f420e432a460cacd0c7f29d2e362f93669f95c37c7e2393bab2a8207a689597b2c9b6dc552ea2067adf69588762fbdfb48694d8f2b13bd83213b3401a9df73c7ccacd5f778628b59f79f2eb017f5fa46611c180c9f231eb1cf63cef2b771a73647fe1faa04c5179de9f8cd35ed1ca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4e33fade837bb4c5bcb9c3e24e209248ffdd9597310d395be78ff43f128fe8759b39f16070adbc25b6bdbecb61d0cadcc44522e82601196df02de5ef1690932132e609704ba3e6b8d06a83c19fb1557d6c606ad7ba0e532c417fbb79538b090558f66812db462a9571fc1a3fbc56a74e6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b49b088042ffce1f3e2b81b94fb911c74a0f341d2cd0e70980b26bec3e40ff12e663c92c4a99df912b76b2143999549d6b3461fc810591fb0d6e4ac3b40383ad9d53da4e904bdd9b05bfb3ebbf143993b981764d61d554ac19b368f5821e06cda1c9a601be6d6d4d5f2417db9aa73180;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb727a2109e900271fe1a8012abcc79ac7e4f19392fe171e87a103233deea76e7cd01c568afb918800a9029960548fd31eeb5c3ff66fcdca46cd18c4942d6163345d2826b1a6d5052b2fcb5167e8b6777e2c62a24bc9b6e3ee2b2ea9306a26d237e3f551ebf273fe80ee4f8ebf7d49a06;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87c82be1c114ab6650d6cf44d1d9a7466af295c9612e73a4db91de6f82ba367829cd61f6a7c4dc5991e39bcb1dd5bfdcc6e7bf6e607d4f795c07c2f499907287332b003894a50be70286d9da01c4da7eb47599d15741d3f81fa29dcfd487cd3bcd38e2bb0368afe062775c4638f85185c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he690b638f121641145d8a7d6776056ad7c116974af5a67734853c5c76c828c11bfad9ad9280cd8568569e834729cced5bfccfa75b30b7fa878e365bdff622578f317ed34bd20dd2206e69c136832d7d931998c5f5067e9f537f50fcb4b0ba80351ea1d172251d47251a7acaa6c68e0907;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a843e950179902e28dfe8237951ff73129d85aef0c3eea0873a67e41df5c918a3fd401450d5c3daffd4f90880ff713e63c55706cc35ac925a7056cd7cb9ebb724e864a227e9231f7a03c29cde7eb8bfc9ca5b004fcf86dece6c33784467b3b5b958cba80efb5a86117bc05cf6c684863;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h508eab01cc3206a3883f12304beaa68dd4cca38947686ac1e05414c72f02186232ae6bcc8a325c95acf4aeee644a0e19d5ea588edbf8622e56b49bd4f3a0fa95deeec026b763974f45e7f554bad86203c6cc1ed0dd7b548766d53ded602e730eedcd980f6d3e8cc4c97da32ba72856c50;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h554fa275bb22ea6016a5790073637eed0f0ae482fb29c3aed27d255cb8c8bfacdce485c8f3430db95a2c414dedd37116192d4fdcbf0182c526af198e2670d29455fd50202a15ada3f38c5358cb3abdecc44e1352ff8f5fe0ffbff77fa043aed0cf9b385eebab44d113436a55ad4758699;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6d048776c6c43435f5c6b2bb622764f5d95f9799109c9b4d9e74b8c4329580b097256831343b535e379fe335da7c01b281bb3febf0ea2e57f05489fb867596f071bbfc7f76bf6675c158e666b0642f4fc35290bae65811c940cf17e0d179f2c302ba4e3db6b23bdfd578c8c112807510;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89806b3f29f7f24ea22971f5975ae55945a590a2926d68c05dcf8d12e381118d45e4871f0aa803b9fe4857e63f993267eb55644e1abf32f38707f5951dcecbf498d5514c0587cfc362ff7d06fb4158a9b4bd458a18f503a8cbb42af979536f82eee592eb26ec5e35bdd30abdff147e402;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c4d0da0142caa97ae4307d65d717d245aacd50debffeb13d3b04b6751986a5a5b24af4303f253aae9e9fc52f3f5057d1a4941340bfd3ab1e1a3ccded65d37fc1c9396ca2432ed49ff415d0d205544bc81babf68998bb593711a5d2d2bc5fae2c046336b1d9a6c4371519597a99a841a0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29838874ede27046d7a04a0a6c2a701d12ccfea8a980096eabc23a27175b8b65576d0ad0196bc67bff84f36e7178738bb8a1cc84a834929ca87eb0fafdacf48a2c620a21dd14f9756c60b34441a61157f39bff6cd948741a2aba463901c585774333b23ad882046854ca339a0d273bb64;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69b3670fb5c4eb71ee9313eebfae14a8e0e180a011f112fc566ea12b73862a3d1fcf7444539480754ed1335b3da7b7a5311ac6bb685dfbbb792a9371799f7149a5ff7fcf14a6611c869240e5a8d990d6db5da312801836eeaef13b179216048625fd51de555284e3523359804aa53324a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha0f34d8db88a73f05f7277a5ba23fe5bb8fe10b32c2351c437aed1167818b18dccacfb7ab77616a798399181c2589c1b62455d4739d147ec5c824a4c774dcc6cd61d4015538178c07172d6d86c28ec8359eaf0a1d2571cfe3e6d10144e52d50d05bef79bab972e21942e12f83bd365775;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2342f3622b5ae32296f7155c624bd8c59e13bf4d8f1ebef682a68298afac8c8b9aff6ef9be1bc737f69124eedf0cad28ab0770b4e98a80f345fe1e3066bb4da25931601f11958f20ae8b9545e3731dba422a531d3dc4882e3f3d71fee2ce40853624f909e916bc8104c7d5fb48f5375df;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6852262e40c76a720c5d77e30dbe72d87e77882a9b9fc4a2bc58e014eef7e812f2a0a3fbcb35d4eb8645532e4a382f95809fbe45692ebd55ac209a13fe0f3e2444f64e8db1c47f0fd0586dbdcba8dc71420221fa93a5ddaeda84896690470c97848046895d45d155f001b6e0a2f1941b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h884199d9b0bee851146a2bc41575411be0ff7480e2458661c8a63acc671db1bf0ef60b5e27408465ef91c5257fcf0584f6138538c3ce6d76be527f46dafdc8b8d141c86cb2075d65b711b8ab7c407f891ed9c6876e286404055ac9001488480db40497b7d4252b094773b57a9c2eec1aa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f7f97fb800aa9682b1a5d46f535ec014c3683a1c52776b2819e6495e76a358371158d3780355cecb490e5e7241a47a00a7cde895e7715a01112a15b5b317def8d08077e267950397dd2e569063768befa9ae55b0cf9bb99efbe7af31aa4ce96f5425fe065fd68c495600c51bd0598f4d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3973568cd7dbc07e12bc1c249e105dffc6191d1097f01d726ab6423225af057f6ded48fedca3e4d364a74756629bde5158f17bc18da5264d0626ff7c36b7be23f527fdae09e5cd63a3c80693a4beb557ff3014b86b2f9c33d9b8f16cfbf2a8320cd2b5ee94b716191b7ce8aed6ad36175;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb8cf4aacd1f65876924eba85a224e5dbb823de99d7dd92e86d43338d06c4d720e6f50e079dae9252f918c045e4704a34c2029d3b5a990e0cb742f0550884cbd740a57f405576da2324dcf9984455734b17e5e8df7db66c377221382b76111d30c9409fcb4c128521be71c96165b8fad7a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c2d0b56f1bb21ef29d71163412f108574a21acf26dfc1e0af4e91ba1ac82657adcd306b067ebf3e3653e0b5ea1107ea07f4e8cb11699ea051b114a323ea7c026a2098db0e42286a89db53aaf4eeea1559c770f1535607d0c40f4d0fd9c152cce7e69c634209781b451f09c322b050d7c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5dbd73fc72e8d6e38467cb7f8ee5a4e42a61823303f433c92e7920e35f4514ed75f2ad29ec4d9676cf0b23b85ad07cb721dd0dfbd9b89be84ff7a3e5179b82d23e2bac9dcde56bb13111015a622150fd63aae9778c5e95b39355a18b7a54a870ecb77fb667bd45172d5ab25dcfe5c7c2a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8bb9a1e4cea717a1ebbba3031272daf0096a3ae90b8d5ddab1da7b078148a54560832b91bc4a4e5dbd83adb13c81066b2f96c8051b01c251cc1aaa8913f689fd480de826681d9705f702f4e108e9d3202c8fac5b85aab4ea61a586d8943f3af195be2c1043bc4fa646bf11f930f7dbe4d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd1321bb82a4826f4d8ad38618dcf8c615e86d560ae0a2ce3f549885ae9d76b066ed935d8a78e618c07e434f6f9f8cb1f2e82e85bd1532bb7af8305f12ee093c2d330f3160ea01442bffce67a5ec2016a0645d81d90c17d13f98bf3facac4d5e533a5491dfaf503a81891bb1f71bec749;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h342f6cf5d8be54a9deec378adc6ac6868fabf8ad5c3730bb3b6445c4a750309a0109c9189ca2937ff895a597ba54f1d0b1a4edb9640161955f828b80111d2a5b8f9a8083d4af055e98a3d4bac2c31a7684789e0f40db5c84a349c2eb4abc1bd9a0aa06638a62ee7345464112f04dca1d6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbfa0fa20742655e096f148f5bbd47281c4d5248b0191d667b53b5d5cb1a97640ffaf92020c68dbd76f64356be3b58db351ddb3198b4a692eb18596f4a4f6e9932784b991baa0542469e0dc652e28bc9874c9472235dcdbf80c868ea5579ab0b00e3a9cb30e76c0f2c7bb6d6fb0c19f836;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98f56163d2876fa691d863d10ceaee0caa8010338dd9f005ece029bc72446a46005b3e8564f53d4c1133bcb187c6823aed55e7c9f3ae5b0bb3b8b6480bfee190c92e8f0694b0a483a35482fa937e0ac226c67d8a9dc95e4ec7ca4ae8e52e8e7fd888758c665762d4732c8bd7829062cb0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbcb6b468a5deb07dff3be363684d57878328012e47a361b866e08313eeb18836fccd8937f4107e5b6dd4fac93592baf9c40dd5c88ad43d2cebecd2aa7c8fe55e398f1fc9e98b88e8ac0e76a5248515f78afc41234cca6ba56cd9fb174fc73f58c894a60f0520d973bd7e360660dae4566;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8ce6e865becd664c45230998be31778f57c34304776c5873e8d47e60683876c5ecaafa95add31a459d2ff39a7838925a96e4ada66a946ccbad079e3bb21d14de17c5ecf4d717d96da23854750bd37cd429852c010e091299851ec6a278e039b54a23f0c0601b4ad73c00aa57722ed25c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd52009ea468c212768f4692551fe693e8848a725bd460cd22504f7458ad499662a6b42372f5295c0b4ff00b9402146849351c751c57eeba76ab759c405981d8492c9079b96d5c47181c5eef35f022c60c3be130fdc779328562d7b5cec1f28b06aa8e26825b8b989f678a9fdf11c51461;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h16816ab9bae3f8238f020972a7d3472baa715d42b3fbdef2748b8a197c6e20a55ef090c13db6c596cea5585893c97c9d3fb86099c020c7bdc578655385bd605e7387417dbe96c00f8a218769649d8a1f207f94828c447abdbd2f6d4545b75d4c9c15b856014678d33a385daac9a453593;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f3bbf7fc55dda23ce32d8f4753f7224287952f4951f54dcd990b041afef7025bcaa69dda64f89038a66a26ea4739aedc0863b9210555145aff8883f94505335eaefbce7f35ea10237416b85cd0b12f7e72901d957cf7467f7d2a0cf0cc29b8fc886cb5429e99afa73a401a487b47fb7a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44dadca32d21ac470ec83f0a742256154f8e74e926ef84ea1fbcf5a8379bcdc7db3dcaff625f620296a7f7db8d258c91094dddde1e4141ea1bc99a3acd714517720f7d1569324a6ca66ad7f9e69cd63643858a6ac7a5ba6fbf476cf9166d5f40a7a7dc2d7372776ec3e4f413530f9481e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfafa7984a2344dd5e3b04635b2438e8cf9d8dbb82285a98b5978bac23dc6bde58ee54e15b8eb426a8b314dcd12968e9834d4e513eee615137b9d8800769f442d96aa27fb885fa783cee515cbf23241b29851d3961d57ead396eb055ec843782a489956b0ce450f8d06a9054e037474bba;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8c4dbb7c3cd13ce62623ab8c80aa82b0b3676b134c27fa7563c39c6fda0a7efa30a3d3d2d1c120aa6309f577254d2b05a88f367a1f2e7fa322f22360877fe1715a74a0a140aa3a9a1fb93e3d83b7200b92261b2431996859b61e54ded4ccd1bbb12a5ef8fca1729f179857c30641a621;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac3eb7c5409d74d520418e013f78b39e4a95941dccb91c5a1238a616f9bab61a675c1eb6fa9ee4d532add527b94b100765041327185fccfe503c5a2eb52d5c4c479268088c753237c126ee4fcab06b487ca7fe0deebfd07ca9b9b46c14b7ecd57a78db90330107995b68927697225cdd6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h33cf15680836dc730ef9c10293715c9b145a8830f87dc2b778d618e50e474f6decc0b80bbc7efb9e543815faea76ba1c13056ca8459d1d607128b1c496ca0bd38581399d07d468b3c78dcb31e6bcaabe857551ecff9a6af30f74c3b36a69b8b6058043bdfee44e379b644e8a3d638294a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9fb5a7c6e08d58a141179d6e29fe1751eab57b39cebd596db32d4d2696d803e86561b07ac1c2db4eaff5e79c0df7b6622233ebd2b39817b253e1170792d5a60e730861852d703c6ca1c2cc712df9db213333f431b90f9da9e1fccfc60b4b5cac7a4ce434a8e2914ce2a9525511aaa963;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc9a4a2bb64cd283a9bf71252a9de28704502138aca73da73859528ce20590d919ee6ede8c6eeab4331ae3ec6eea927b72110234f503f53652e3cd81156a8ec73e10d7d1ddd960e9909e0be67e77b373fb04e18f4ef01216d1d351171c6dd5937d184a81cb08291f2412daacd8f6a8779d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a0f68b192707a8f82a6d778eaf32a2527c0b5ec5bbe63a8d429a165f76a4c7d09f61f0c60cc31aa40946ecc3935c294da5c06a1ab4fc8ac8d82b21cd0e9d0150a8ce5e64f1c79aaef91cb4c983678abe15ec78cb44df0e18f99658495a2d50dec661371d07dcc24dacf2a87b3f0ad46c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7923b3b5d54a020bd73d11f4616872e10f069919d3b4766128a60e067004258a170980933e44c5afa71b69ad2f76a9f93679f76ce34eef41c7c10fda45e522d1abfdf89fed71cea4d0a6922f045313063576d1c47e8cd446bb602069eac46513884c24adb100b3277e759594cdb55c59a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he4cf82c233e9e91a115e1d0d2477f7049bd8a477b1de801b2b8a5f8ffcbc9e99835bb93a8ad157aa5696f123a73640eaeda764ec5d73132b38c2e75e15928f7535fe17d1161db1a93c87c7a1f0de806e8d3dac86064d41626f570eb0ae6352eb4d1fa6850ad78e6813e04ebcb858a2399;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h357413e39d4f29782d90c19403e273375d1ae996c956d53dbdc34b8b5de91acde907561f5c745fb9b9fa8a292bccc5b473b0abd8f5881dd9f79b647a9f61fadaeaecda797b6c2854f437525e2e923a6c8a930441208ff548c86b1a5115bfd91f7c7be1453ff49ef0dcec7ffc3a03b593d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda31e1a6ea56472a3a42c026601dece4840c8259ad5e49ea7169011050f6bda9768d37012b3a63a1d8c5013d26e70df1aa4d12492162243bf7487fd656edbc0a38ae419cece6e2f41674fc792f9b38bd22f582ebb260d31b6ce1c3b87c11ebcd9fdb8d545e0528fc59cbe5e81772932dc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21de4bd9275091b0d7902bb36b3ff9a8c68df6fc8b60d3e52fc4da71262d82b3b36357e7a7a54080d0f4b953569700c71f1193f6d566b7fd6b4a033f1870ad33d6dfc125310870487ed6f81aaace167ceba11019b76de3e923603e030cbc439e2842e0527bbde7cd31ea837b2f21a730d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc99d18e6471b9afc6692154f22f72da872a0a3f171ecd9c1704c4cfed65b5997493aaa7150511f0c96228c2b6328ccb9799051e40a4d02c073af83f3a70978ca860339ac9777b14ccd216de54d23207bac9199c105b0d075b0879657222a2616829944e5d8b2c040e4e2cd69293c6ee05;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h402c2921e04ce850215533faa470b8220547e9fde7b33c80e3fadb0c838a1d4e0017870d952192c6078340eb429faa9fd92ffc2ee6dbee31888ef9e21d53e29664c769a22b75ebf6574d22051d0bfb78f3645ad66fb70a375277faf0a9cd1664626836cab0f4b6fc4aa176dea66795458;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h592970bcdd69c8c2e7236336c8a288c9c8aeb95654c907e7a181630983692afd73a28d205df1e886a7791cf2b201623654fd9479fc28cf83ea008c601ce3464206213856dde708c6d38bb37e90f386c182497459a863db0a049ea2633e29c206358ab1f24b40be56da849d128ef8cd2c3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d6de85611e84af5e6a7707780f099b6a2e2d81c72f79b84c445208348a63e9d01abfdcbbb17b454962eebd7985782a4576be844b9eb194e5976aa01e47d17bac32cfd32fa067e53c6b2edf7fa0dec87f07ad8555cb05a979b82ac07614c205be3f4b14b19d824a22cf19cdde742cbe7b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32aae6e8e024d67300a269f231f4ece517b5ae55322d408d05fd1497ec062df858f9b51e033b64228a0053c26a36d85a6e12faf3429637204d544a5f9ce5cd50016a6e9abfbbe990587fd3077905f31a1e7d3a7336f259476686c16680362ed7b6e4f6f32ba69132c81b3ebada18d93b0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h19e81d4ebe0b773f3953d63540cd183589386d8d43157034a8e44b7c09f029f8a60ec25d544222aa14ff3f4c54deb34cbb85155e5cbef36cb9727927e5a019a462af9ec75545c9b3cc9abe477c956773e2320bc4d786ed42aea247b2d400b44306e28fc706c4a0afb65aaea6c31e72826;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e3e973a85d3f726ec56eadd08af9a71086cc58eaff4029029adb18ae1d151bba687a8e1e8467d5e551162e50adbc10af181a9416c766e9019a222491de3469ccf83c1dee64c7ede8542497b0ea368a95ae49353c9c991a06a2861b5402847cd0a297a8314fe63aa86dbe7d63bc5b989a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3eef3fed3b2f41921aaf6c8c6a569096221874b15f9d5a89e676290d6612d1169861ea25e03dec08ae6f4657fe06e9e778366b49f94041869181a105c95b11df08e1504d95e65389df0d463d194e29b24fa3264f453b1bef7411f2b9426c7c81f4d5268203353a96f859feb85064437fb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9e255296ea47699dc74529575ae1833c9cef4d91f400120a85a93b267b55e27b9b48bf41afc739bbafaa480667c54cbf73c8da4aae1ac4c2211bf7271a392d8f3effb04bab1fd421bef968f0157e7592a90e8124e75418247546a1276b9e24cd16cf56986e102cc97be0601b690a13ad;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc60be8aff29e3a4e624fdbe75974a68e028f80b920054d9dd35987be5c8b047a28c6715f4a3f1cb1a2569d4bdd2eb96cf371849213b01b788abe28e0cdb6c652cfb70ae843d784de0fc5962beb00a29919d6bed75def12a2acf525af385c53e5ce912cae07a90f84b9b2c1c03c55d5140;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he40630a0555636e2f9eabd6a5899c0d86ef4ff9a770406c95e0bc4a32a9c9912edc7c92be997709a917abeef6c2b01ecc63307b0c3143f45f3c10ae7c5fe1e98bd368eee9e9155fd7a6ac2c6af280f216711c0e7052ba91d64bc4dbc504a9ceb63f7897f3b6862135558ec25866a52083;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd7443cda73300f2223cdeb46f41f38bca2b24dca3cddd554ab29b0e31fc17ae529243478e400a4cd48f9d7a6f24f400318fda097399d049183dc8f30de33095889b2d524d30965260700e2d8d756d427032f8993e984429bdaa62980d82d47d44ed82308390f7e3ec93497c0c5830a279;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf73e37c318beeb49aef971a8125055a354b4a6fa2e52ded900eaf4def76986f449a30c1d343b98ec97df2ae198786b2a14901cb440e785f03ee13f0ba237563e9ab481df618fbc30033c9b4b698b765bd6a4195953f8949aab69594947ec0994dbc7621e53a317c96ddc5cefeba36ec99;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfeeb4c017d1e0b7c5196c031fc708c9bcfd62a96ac9249ccf9b62c08324749464d4351289a839cb3ed898d1ff30cf0383f9d7979fed32fa88d1dd3d488d16c72f2b7d54e14cce964fdb15053aea7aee41361239e3661be76db4d6bcfae8dfb838d069751eb8cbe19d54ba14e1adc1eeb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ae590e5df83a01a7c7e4b033b21c71b7247bb57c7a20944ab8998bc678d8397fad572c781bfd760c6312a4cdd181930af63b94da586dd2ea30698c4079d489e6e2351fd93b1302145a22a8ecfdf6ff80ad4bbf641c382904aa384645af1aa2cbde9a8be69d34c457805a510d8897f386;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8a63af5ebfb3925312917ff6f193aea6c21f0872bf835f599bb0925fa952a0926c94684d30c880343565829347100b00586cdf380e19e5e57f3dc8019c3d5973fddb0c59d40087f5a0277c636455d8a6ae0cb3909f52c95ee3a1dfb6a869639a74846c0fa0c0741d1a79948817b4e876;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8eb30e9fbd8bbe3326d194105daf3041bf41bb5d8a862f8e7989ac38095baf8ec7768c0f557063332493949a0c01d66db66ebb40a5fc229bf64bcbe2b095a0425c126ae936c81987e80ac86c87dd6a9e28176598b1b5ef27a59325e0578ea3bd9148b8f605b2da07b3c575ba731eed6c7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f14202261736b19a419f2b9a8eae9d31428d3ca1ee80c3ca1e2b3f9e37d98f274c458ef2596eec395fb1602d48dc912345132bc88bb735665cdc4c5a23e77be8cc74533b11a98ec076a8ef249393bda931854d24859c7454f925cfc24bf66e3b57ac49132953afc79b3631914b7e6f60;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h617c85a2a718ccf2a4cdc0ece5eeb22802c8208453fbd46dc2313e8b55f499c11ee59af5162551c6b1fd7c5e04e059f8ee4b9d4e98902bac8f53e899d3b8a299c24ced197a7accd42ab42a77459376aad33e19d97656f3b08d55820de21a9a3a232bc912c7ecc402d4631a0f90af5e09c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h946c02232c70735208535bf74c6af40cb761acd41c3d1a5ca2872c69e59897223e80e80be7975a51c6ef54d59668396b10d1ef3a1d8837ec43aeb0a7700f151d4ed30505ff9adeb5190a3b1a549b6fdf5218f8c5cb566faec76ff9c7f6a46b47b8e62d9e38d9dc70e3872d4df77d21ae1;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69ee8a5d4038e9dcb1188d75a36bdd8cfc1beab7a6dcd9c32b3e851d8dfa4a4f8b24bc6a2fbe97b55478e63859eb7f667b02bb0f6a27d2f3b67c0b7c4ee5cc596c6dbf891d9a638667c46463e99908dde658832a5ec04c17a4072da50aa5a758b4223c361c62f16e7e5ca6de6ed8d18e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8138959f9f7ef40f8ac8d923bbfeb21e51c409ee8e688fbd45112b3be16fbab68d0923365e3991d8da8b1e690c8810176c7bbd6e693ac73453ba71b01dda5cd1ea31aec3cb1d8c9b095d73ca52eaae7da61ba5f714992c6d396e8bc63b423af4da51dbf6245705d566d93c1929212c00;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6a5b0241b429cebd37c0c50e071933cb565e8adb797db0b792804ae54c8874155742db10eedc1233107a15f4c453a219695e2d5f7a00e34c5f02aa8d99e5d8fc603d3af2834bebcd3fa9f74b70aebe8cec914d3de2ca96c2df4619fcd2fc65282f40812150ec8059c8b9a414c7b0aaa81;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h16f9946dcac3b6b812c69f1d93becc51dd3c8d2332c991880815a3acb3518601479cb01c7bde53865fa8c872dd9b73afbb6d50b87864d523acfefedecf2d60645eaaf3fc915af6b1f75f44134e69ae031af18895191ad8a2c62700facad647463ef8c843466729b2b7a21fea635ada8a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e2adefc9294ac8f890cca3652f299193a7906b2d70943a5909704f4109b505de4129ac6da9507973064edb9d69e3dbfe971d50de3205f83a92d3ab5744fad5bf2f7973b2119a60a337f20250f84f8ed55678b9a24ee931b5f9a407ed547051040e94954890d2931dbb311c57318518f6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbfdf8d2c9155145819f4ae7e3da466a0b0c54fc61c7b564c084613293ff54019b081e98e9f2640c4ec8f6f90bb97f49691e1e7981be678c0a3fd007906eed50547e270def6a8dfb815cce5fcf87a276150b36836f0e2f6fff93dc42b69b7476ec219499b84d4a821a82911ca559147e21;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc842c9c69c1d94d00e9cf8558a6f240d3101eceff5b7a95e99a7918b1df6be2bee661d0da9fdf6cea8c232caed73697e766f588e32287a92842687abde866e96bd92facc38a7cf87a40c1150013d2832f61931bb9e3b0794585d367f67266097ee92ef1396f3e92449687d1f28f336cee;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4fc73d026df1c7121d85a261fd353966be27ce3219c91bd4e3a9f9e8b009155f56077a8ce4fa01679a1011ca75ff120d0e86dd012c92ab419c061bb14cf796a4e0da6883bfb33197c6ecf9a5c1e60aa6c0e211f5dc88048770c8944bef4c9e266e53e6211e0ef51c80e802b6bee0dff6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc17b08d3fe3f177a0b29eeef29f57a1b33edda3615c596331d3e4a74451f0d913b736ab33b8618b5c15c85aea86f857f4294960e4ea3e71ce527d5b9dc97a7b96bd129d415a48d6787789b6f5f1f56e1f3e17d2355118c423bfc2fde81aa5a66f2cfe90bb72278356e301d4f2944cd325;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb175b6e138835ad21b16b25334d1bebe95c82ed15f480dc340080828fb6f032863ade4317b363bd94df98eac8200a338fa9e12abf07308f0cdce6bc589d59fc74612131bf9e47c7a60e2ffaaa7c9a8609f50c0670936b08232b77fe0b50d3533056efb415786f9e425a9ebec30e4e452;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd33e300a67456d330a9992c0eaa2ec566e8ddde7c89ea0a9f861a35b9bfeac67bf0f57467835df33632777c068c9a92a9064ccbb124afc2b789f74c5e920e2fddd124c607cea7fd4ee8cb4d54748ddf959576328557421727ce57b9dbd92b6f91202d1f71f904078613deb83c196b5a7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h386884e0aae281e9cee0ffbbfe0bf9d54cf346ec5dd9e72b17a4b0b042603c3daa8c5379b919baaadaf66813e10ea88652b902f3f360d49fdad863360daed918348eb121a438b225d91d737ad45544b9525a2596bd25f8f3214f28b923c9cf2d0773a0d71c824fbe34bd50f698aaebdd3;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hceaab67e8ee52d2691114c1a6b206065f33102add75b2a90c31cf9a7d2cfeacb0a238ced41ff04388c7bb62931f591601c75f5d5c3f5558758f4adf7c99315ef9ff1b74a8a3d6dc25529a23b8dc8b214cf06c4ba0d85e6c384b57b2ad558f38d791de5a635f41b257aadcf86a2318d360;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f2c3373ffe7f3aba9a5f2392716c46a0565015895cc695fe2d01c4b6b2de96e5162682d044d82cb6a5b88b464c3e5d3a09fcdf8235de52a86bf38af7a9480e3637d97444e8ba2901a3183e8b4819569a47d735b783d3410ea565d555e8ef0a7b055d90a85a6c53340888269b6d56ca02;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0723725ab46f7e5f5cc808069ff027412080f49446e890ede659563ec8d0509db29c87c9d17884eca195c293c92696aba1aac4a0e52c7d5a2a5d397baaed5786b9ba1971c0b06b0df95b53e260ec5f945ec79bd305b445b6b0ef7bc05c31cde25e64ab6238598c65516d0e474a57aaa;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb92c12c3efdc4e3ef30935eddcd86072d5bddd22c6e3638863293c3cac61915dfe21a4f3a3483967397ccce14de45412e4299d4a2795580db23d6870f2b1c74b445c670ebf762eddeb239a2a953ff2578879c8e35079d7a9827c600e00b60844f8324d84a8487c248d00ab208abe2a7d0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd9e885b64ed961921b778593b27950c91039bb46a399ef284b8fc103d612a6150c5618fb5f1082ad2b4c5544b1b1dbfe3de7b177e4b77e10cc25408cfc3c1709b0b7c809ebbcfc1cd138e7c6422072499c3fc93d56b3ece1f4002d6a66bfd9f34be66dbe369ffc4e97e886f0e0e0348e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc41be9ca21461bc80be529b9ea160411e712e7a4a370c076c52fdb1ded1358af09545ed423489aa6412e7906735bcaee606fdf8ba2038f31f09f17e2cee26061da9146487f310bff4f7735ea08f8c099e3e1ef632be21c70f853766d1a212d45ccfaf74fe9b5f523fe958006ce5ed096c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb306a69406d571e2e81312e12f8818534113bffcee79f275b11bfdcd48bf7fbe276dd0e1bc15a962283064b393c33a4ad6e6944b1cf2ba3defe3c06ae41ba035223426db04f59098778c9db84be6a048c40c03f8ac164efb00531d9cbccc4d898ed1bfca475b1d8fca2e7823482e05cd;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd44828966161775c179471050508440628bc880ee38324a49c34322ae7b0f3f82138f97b7985a5f37d5420209bbc59986dcf954978dab286c60255c183a3e6d61c8b83ac4cdf8dd960fd7cbced1d80d0137b20f53e29bd73df4b5d32beec3138500f861811cc51bf717188cfc48ab0962;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25a6813bb6fca73627b27216463e4c4561436f0136a580d1387b2b9980d25c8a0e3345935f82ec4326ad0a4f77cef9b99f018aa1da9d1a826ddc8677e0545db266e561ea9439a2fcb4a6a5a5ded837e479c599cc341d7258657b8192368e16206d4a60103da6a462daa002d2185547cad;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb4abef40234785c1d9c4f5d23c34b8b6d87bdb8748904c1c831868dd4013466cb4325c226f87cfa07b7ea5564bd1f34e76f09a1e282c70aa04b34dc88b9236c646eb7be3773e983a6d173c5ce47cb1fd3c8477d03b8987b848d5b6b68dd3f5800b64ff975909ae8ab00fd991d429846;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75a80a69eee9e7d2b804437e0f406be5886d0ac5887a1650c2eef6fab39f62ee5935df60ff5a8ad19d974396d19adbf7fab7faae583232e2e1048c9be20d98fca537635a54dd03bc2a03350abe18eb611242f891190c101da45e6264cdad03d8347e3969af60713f04bf6b2bf2dd8c572;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he63d4ccc0db3a4355d7acdc86299b9e90f1fd02b91cff0f74296cba776703b8bc63b0fa112eaabad13fcbcf11ec6c0f825a7bc50f1b5c2781f24b627d42c9a15a7a9436c7c166bc3d1b4807541b0ae0ad87e1d421ca052775a3f5ad178e87cfd00c727d3f8764c81737b5e0bb0bf06285;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c90bd8bf3d962f45bb9038bfa0893c1639299abc8107c51b7e79be1b89afe1b9932b0aac2fe7f312486bb098e88a0d686acfc8a355d51fd1bec31050645a375d8ec5d17f6655b921f517ad9b54cc112e4507262e9c95a84a00b823bb6a63a85db2e582210f525b9cc400a5d01d8b3413;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h628ddb9cb64de3a212ea1fa4fa76b55e617fe32a34fcdb1e0a882d9b69999e213e42b3ed36eff60b24f550a8abe920250b611da2d0053e7802a7ad76fb961a5c95afb30cc924869dd0b152ff15bd8dae841cedb4207d5dc11432e6f8380e0d4750f204b44a5cfa4341dd6ea9a19b6687;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9351c6e03311ded51b85075b2bbefdfb462f48e2016465499c4d3702ecece0f58c191199aecc532cb0cad937d2b0638d86e2bac1a7baefe0a38c8db444bda515afacc9ad277a9c40ca621f733a8ac27aa4e649cdb39dedc0b4dc9d7b32f0e8fb25221ac57d19c705ff85d1e8acec91a6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he9399c0f02e9cf37b66cc37a84e84dd65bfe67b52c3702d6670ab3e3bd9113f6a3789538470bdc6514d75afd417fbf116f12fddee6e19394f07cb55b923a34e1d2ec319bb5bac90e4e7a596a0f6e36b35e60aace5b7b70722efdb043f16f1401ef243c5a6e6130ea6322cae4044e0477b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d11c8ee705f092629d354e72383f4d76ac20fe98cd50f85bfa7c338cb359b10c343b91d42af8c1692a5c9b5ff6df62a4ebd4e070ced2fed0db9768bcd8b78270353fbedfe81b6ef4e3ddd557b6874f97c0f1a24ec8268bed3f4750696154812ffc2332af12a6af0c9487ccf762e72812;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf28009e29ff28ef09b998509d498d98c8c1d8071f4b56d09a0a0dc6b41c8582dd232d982ef87035986ee94578e256b32ca6ce6e145c947f9e2a9b7b4988581b0cc28e4ca064e03e7ca467c50d95d29cbcb55dc7014088f7197079a3b8d21e9b41c19d69f454ec83c948c5b159d28374c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7af20fbb5bac3a312e30be56d90f863d3b441574611aa303ad7036253722d9fc1e1590df54e807b22eed6bec205e1a7133dd5074725ecf3a3ca3f0e3ad852fbae51b372ab87bc6eda964bd94f1789febb405434bd650dd7ceb4782c116c5f58b9e04551766878c87b8d18fb68e9279e96;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98d0982d47761f28fb3e4f7d2a4617f122666480d5f315dae20ab19f86a98268371618db78a8574bd336f22db6d8bffca20223c8c81b674b18d1d4a2d8bd672f4845dbe041cb50ccf3313ff364bd0bbfb12589157132400d2a3788c24f2448ea71310cea293589229958f5537bdea852d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ee63792a6acfa9f6210a34c001b96fb1879bf29e704a9a36520e8f89b1cf633e1914bf0b955bf0cf77cb7cffdd0c3eb8d155b63a33156100d3565d4888f8b0eb76b9ab659811173cacf0d893ca05b0cea33635bcf482f23fc211c4c1bf8e21c38fca9bbd1d8b7dd9cd02be05e9747d5b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h877f3a2a983972d7f2b9359741f3bdc16ad79b2026674e5a0a7a4669ab3177069988dc2477cf3382ae618fb5fb9ad4b880b65897dcc98db0246a2e2df12a05c13eb458c943a621029004d89ff48b902c71175adeab24f055d6b6ff48918d5ab8321b28b5b723ebaafa24154f227cd73ca;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7937ef5338bce903fe5849e158b8a7557fd2283ceee96d0c3f132d799ee8ef2b961aff28a642e615b865ea0dfbd42cdedc7b6186d1e3a02caabe8a781a848d73f48c36c492c241a4d3b0ffd4e5c722faa8ad22ecbd68840caa6a4e7930c739a6df285ff0ff90cae58ea5a134dffc4643;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ee69a0df82422468cdbf8be2dd47bcc1020a192fe67cf71fba76eb062801c7623b8e0795a06d4a8253a89cad43cb8cdd652dcde33d3355a31241d12c3a7771a86c9568991e3774703d9e2aaaed011e7e8a8192217dc6550075c246942f42b968d31b67d9fe5f0cca4281c1929c6285c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h305ef23d100efc4bac9b316ecbc4cdf9b5f4cd6365b5ec80e900a2d6fc34bba17332695675f769c1889efd902bb62ec1ba1c655f19951ac5abf35adf5761cf1ba177c46a6348ac2257cd494d71f9c02e6206a4e680f67f778d596b4c042d1cc2ace594947469cbbf0875d65938f6b86a7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h830f4388b707d49818e6bf094932899257c61dcf94861a1164b57e599b1bb75304b8532328f10f6678d1df3cb508b19b19b6d37d2d58ae7eefdca0d1ae272ae1a894d62c601f26497d85c0db0a2cab6f335a928ab7cefc9f1ac4d0275d2f8a4ebd5b392d50a8ec1d668f7175693176912;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d5af1fef9343b2cfdc35fb13e027a98db5a2350cc5e9819cb2969fddc14bb53187d4d7373c83e6b43c42185dde727f52582f13c12f01e1457516d2b6a730b497523220a2ab7bf45db727c8109398169c98f7614c623a26e77d2ae637b1d8577b6a3497901be59ebed13d6484c5fba1b4;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h435fbf08445960a2cd939b4101de49692634f3a87f927fd8a05bf22110fe77caba55abfd633bf5b75928f011e7accf7275204d4ef7c8f79fa7048df4de36a8914f1e0b03cca79b3574fab483c2779452bb263c687537ce74f4f9e8d6e8607237c92b7a08eda85fd985db78ce0366e546e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2f6df88dede1f45ed539df521982346c35fa519ce65ee1c675d7f6a9372d12f53922dfb607f539ec04a26b6a26123876c7ff4afaa948e4c39ebb4a7febf7e4ccbb1093c0cdf41a0d70f5105dd0e7a632bb460609be7dac76014bb75e27b335a801ac2b1bbf56c436fc931533e38d8b37;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5edca7885dd923379014385a1e1aca9994e8b16c0bfd1ee7dafe75f8fd112cc61ab2b18fca18c0ab5b5a01f90a7043602504f4e68af931481c1c4248f23413b581a68a2380dec13e6ac53c2112df386dbf58f6f282909fd3854deee5e25d5b05663b7e6877b85492ff3dc82c111227fe5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h67fabf388c1b1652e8b77c24bc62313d7991d0425eb6c888f254eb1efbed98eafaca903871556774af7f77bc3a27e552c4826143f95fbc98f011f0b1a921dbe2aa3d130e1a3e8b1c4778491b858a1a87b4d3924daf1eae34713cea4be3321d5218ebf0db2144f03240414aa1b3b988474;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfcb5302589750c0181796f3dedafefb9073ac29dc4c548acb5430d45c7da78fd34e749f51dcc9f44ef8327cf7f6c3c57eee415c61cbc0c023f757c9b072bd7a3c5a7937b4ac537a5a8ecbc93d54e3b576c20eac9e3de2864e79adc077e245884281784e26b744f960992a54e6ccdc6c4e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28cde31415dba846c89f459fcfd2ee3b852410f53b2b43b10dcdb819d1505e29194902070fa24c3cf419ddc18e4e8aadc4eb94013981b3463e4f01ed63f27545bdd8a3c49093be116e4096e5cd64605d4201d0ea842ea0ab3318444b76c0996825c73f03246fe6ad194ac3f5501f4cb97;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4ecb7e41b7e3c2cf767e0a6a7c425d2b65aff860d28f4e1943f3e58e5a3bcfddb0ef7f70333c987acaa8f2c18bc2995e1945a9b1db74208cd63dc25242ee8d8fcb47aa5a37c7e248585ff64a4ed2e71158abb83b9ff4de57c62be00c52e3d4a1b5bad7b24077831469d0334201ff560a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2aef4ecab3dee50f5f91bfe70610a9e9e564fde39a5b202ecdcbddae675bf8dbd3b5ff269ae9bbf937a2b860571ccba93a8996af016f61865b32158b91579ee2e7e6b0a912ea807c877d495922594420d80a09f447dab3b0efcd821d4a9b4b1d40c176c926c4e7eb496f372ae510b96eb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h636321f40e3dcc971cab8bc49c733e2be7ecfe3fb3a2668d066976f40cdedb4c5e812b5dd2b59d5edd6584cb1934b34705e20d84f40579569e0c5dceeb5ee7f81c54479b052489ef5846c60b2255a5862291451354a569f17f7bb1a21833d8db4f8a41d8072bad9e5a8dbd25120e11d5a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h498e184bdb1ea667dac1eb8039c9f4e0e5b0d34c95a52eb1da3fa8dd8b84dd803e1ac0abc78bd215a030974c8af4725086cf84f8a1da7de7b6846fb59593a56504156d40daeace03c3deb339585db9d4cf95931805c6e372c7f11aa3d38410530daed33df2873d2099074cfe0ff7f6c68;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb6712f771d293aab14969b7c1c9472170b99bb55a78b56eb29990931ad9afd1047c40905e1dffd25355a897c2ff8cb2c1079ff75e4f5f4097ae2fd29b153d3b3ade017916af0cf4d595702d86a25b9ba49f261ffe8fd395713c4ecd837672a19e7719579ae4a01ee5a442d7218d2ab937;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc4ce78d26e8e9808a38752162c23e663f4b6b652447aa9fb4f2820ecec0f6e0121561614098e83412d73f29926eab6ec3cdba3b471f1b5c7fbbc321f1857c6e73e3b286598de8ef94271cda448ed1a1f43d73923e5da0c61fc66615c2c246ff7e66a7c0c32d20371f5a814006365b49f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c49187473576fc38bf1655902b6e525514a59fa42851de6cb5a0c3eb44a20b80368e6492811921779311aea92924282a5554d2d80340c714abdb8c534dc2f439c509afb7be58d0790b7ec37fead86ee9a5f26891e5fb71375bdea8f568e5fbb368fcc2a5b05237144ef0d9570a9133;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h467cac980fefe321cff1b6a2af8aea2fd293a28d3a1f27fb1358c3f5f832ff5ccd83b068076cc4cfd833dab5710578266ef1e123e7900a7deba1957b82a080e850c464a9ae3a0d4b6472e1f61c4aabf94663af58bea0b1420f862f1ff8c4261309ed484756dfb1cdf99dcebc2147522e6;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc92d087ab849c03111719b423f26622457b03ffacfeadcdbad5cced45aed8a42adf0355b62f50b458cda5ccfcefce7fdf648ffc089a4eda04d2e4f36b10fb0ec27b6e5d8e5d08e5e9e30e815ee12ac893bf49bb58cb93c49fe72132390af32950802cd915d0c7f85234d0dc813cfa3e70;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2cd77aba5b92ecee77b9cf3cf9fca206388219da69bdfd8d60f1175e239e2ba0d6ae5e68d092587eb5ff65cd7fb25e14c5f865644f5bcc573211002dfd166d2f70ad89222e73b0348dbd5a005510a3142a57d698e9eecd5beda4c9943486fb6aa428bfaa2e3ef4874940f3f77d5cdf22;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcdebdceebd080924df376a606c0731fda80f9cd7fe8a31b7f80703631ec8c1b56e2005500e94282739f82b5926f3916d119aabae3545d9897a9c81d4649c07649ca2bb481ffea9325d59690201ac13903a4ad77e06999dd70025938e081b5be0be3aa42277e06067d9f17b402800a563e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27127b666b94d4b88fa35057dd87bcca86ee9020cd089fe70b0a797d15d5b6e07f013da4cb3fca9f93750b571317b2524df5659229250d8f88c9e33363c92b00d17fd8a5392118b055db1611fb608fba9edfca7ca835ef36d323fe515ea5822e75b5d733ddc8f77a0e50049a1becd89cb;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3c88ab64a82dc0fe75d0c0e3f394552aeb030dc05e770451149f83e0687f58f2fe5ae36d19eb4d6bb8df85b2adee346147c18ed68da446675fd3d0fa83352c1afa45e1b30aff0a0f89c17dc0769e8269bb9851da0cb53395469ccaac5df9a875084dc0d9a800a64432659192859f6a34;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hceca4385bc5ca9be9d7f13ac13c5342a4f82dc03ac130cdce655b85f655c8966552a5938ada946291d538f962adf008aa32688787011de70fe350e2388bc0876d3715557ec370ef3c163e6f37ccccd1be8c1ea348425727ae2ed01e433da5b0e3de45d7d5d0a7683ea6bb7e5fd17825c9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he0ce27533a0c9f6f534722d24fc316d49603ac906c2f8d07fcbf98eb97d6467cf4514ab28ddb3e78916cb3a265082f9a3af1cd704d0b58a4817862b7979d0caf21bdee92a418bcff557875f23424a2968a3a43a12061bf1a0a0ec9a5cb27c130284373eddb1017f75ca5b40c11126510e;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha956837feea9fce9029be9f06c87732495f776aaafed58d9af695aaaf82dddd859b96abccb2d78cb2ae2ba169ce8c23dfae8c127c3580492dab279194bc7a18c38790ae97c3c85b0e77d19b36d660e78f1cc5d9e12618688d33feafc45890f9a86e59befb3b2318132c7f812da20a939f;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9daa9f59e0ae02acc9b23206f2508d93bedacba0694ac9bad0258cf470f27574961c7777945ac0cec74f02bc636f1fcb7db6f269d36dad28fab1660e0a44b14ca108183a18d073b32aad10ed2b067967dbe9623ff7d7d5490e92bbb666cb07407c8440bc7433e426bc467df16d769ef4a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdfdade557454091be0c4e9fd7605bb92f15991b46ccfd1a6b95aefbbcfde09da4fdbb9d8a47ebfc4c1da753ee205dd872cc7ee88e5f830cb87924c9ef3c560bc3c118c51630a6d04b589f92f9d92ea492331abd9ed5e8ed672c565c9b8f826a776047f1007acbdd93e986d18189cf0e64;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb49a1cb6b5fc68617bcccab0b8cabf47b92f71b2da7dc2c4fa53247977839beb7309420e3d58baf43e12f7c8c07cdd43e6b2f93b9a3acf1f05e0b7a764beda267ae77015e1bc3f81f61e67144f4fcdfacea7eda307ec8171ac4a704c8e698b9376debf1e6ad3406a066c524a185f01703;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a9ca2452fb62535d700744c48b27a751c3237286b86032cc887fab9adc8da8ca3bdb62801a142bd46c8ada03233baa50439543e955d5b56c2c345360df747db2f48bda3080129933baa9f4aad7cfa2cface3f6d4dcd77c9f47e063cb542e30bd8abf109caa307b9b6552a38ac112c989;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he33322db8d1a408c5b5fd63f12bba130d7a0bf6c629a0a5701414c7b4939930f51529d9c2f0f984ec955a7796da4ef2fa59c5b222f4ecce5ddf6966927171c778768cac2223930c1a6d382f46b1b59a61b18e52c11438891fc3d3da5515e032eb5f1f7dde3e8eed71428e16b368f044e0;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h29331440fb9ce5d749475806baf9876ed47b4ff23405a075ed3715398c9ea62afc51b0f67086a492ca27c344a22716a6ca819b8772f5a45eb3a2609a4c86e5b27e0540c93992d6ed4fd2e886eb8648f52fcaa0bfb1a92a53a28c0fa6f13f05fcea6eb1ee8415a28255f2a0cdc3ae73733;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94c2bef0b4bf50ced4877795882514ca6b0e7be04aa68556563a2fc748b63f9053bfd9502eb7bfadb83f23fcc911c291e089b87c9a9cd2c47363d38f7c109edbaac6c8cd85096bf1d356438831ebdacc910225d22af167728dd4dabddd442305f255306756c9542745c6180643028819b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcab3951c41864a730d317922ccac4c923ffdfac835a6127acae8a9c1530c3b58f9962ac3561297cc77c6630cb3a86c30474e7eccaf2026290e0a9c7da232869b8803d50dd2e171137f81e91437f568a7fadcc173dd49272f142f1c544081c70ce1b5582be3251379ba4b6abefc8fff39;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91e1ff8a14083b51e4531fa80e6a09089de7382ac7ee23dd0beab4ac19da1db4cafd9ecef8f6e3877583186d54202e527774aca3ba8c66a22e72192e37fc3e6de7c130b89becb840f16bbbd74c39909d98fda89f1c997d06850f6b040beed92a967f530ca16166a8f89bd9edf86513ade;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51e9f07aa589eb9057e530668bb1b8d479a08897d497dcda91899cee66c0037ff71fa13356aa5256e87d8a60c9728708b3d5b3a76875f9a57f7bea979b296628c569661d698f8b5311b5090a55609c4b71452982eb1d24eff6bddc95c11d34b6f9e90a2c4d06256b0d4bbe25d5601ef00;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87e7e94f836555427e6f3eab30446c84ed6959fa41ed45c759f4db277dbb0d3d333d8eb293082961388cf7e21f10885d434f76d610f74cda6d207f9a4679363218f1cfc6d1ee0f9ea9b4701b4d0e6dbdfb5aeb46effab6a1aa44967ac836f6cdf02a575940a0019f72b3d3e81d221ab31;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d17f93906b9ad85076d7b1b09d7c377927d2ab84bc6c0313913d596986ae01d18c93437243f7e8f5824f9c2d530cec2a0d3b9a023aa90845df5f56dbd40bf9c7f0a40d04b5f728af502db1ed2ff51158d3295c6361f8e90288eca775e09685266807af6a52070cdefb22c7dedda64835;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h222e818b899251ad3490831f0453bdb2f30f7d4b904bb391d21efd18fc9b2ad0e9365c17d3cfdc257d0a2f7f57f032e479a24feda79d099886e77e23a0f773cbf07290e01cc63514a28e44c6e81de033de61214abf14e1095798e07429b153dcbde2f6d2ea46278ca845568c607f30114;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc93d373c6ab13992abf2dc7c97fa1bcb6c4bf58a2d64bac9c908433d1c5d0ed2fc4fa871f426d60f0d649a861c5629808ecacc60cea5609233a3cb12fffcf46fcab45b8270e4d97e5d157ee98692b2d63568c31b0966626e9672f4f8a7ce2d3fd8f1fd1402793076ea3372e0078be474d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h884b9df0383c878135f0585d93c67b7ab0b681fb67ca0e5b43faf59551b75e0b46c6e2ee5655c582255b44fff97253762854d0338df3145e868e62900781e02f6f6383282d7f52502da60c53173dc3ff76dfaa8df421b4d8b437396a32aa90b68d8bec8679025611747592884c8b484d2;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he6fb49016936ae9ba235628034c706ddc5a59fdd8c73e0d1aaa769cd99d1566953fc199ff500e5c9129751fe1537f8a69f768e5a624b4aad9e53f452689a87168b10ae256bcd8270106e4bc472a4777138c03b7e6ada87142353bb1e1c175bc83bbfaa3f089dc66ebcd74472bf7929bdc;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfff234fa428fa9f9551f221f4f6dcf190fea07d0444704b42e3230b3f111f4650fb560ee36809046229832c8fa1ab9240eca2023b7f38a30593e1b948d4b799844ef88a3839f14640a7e23dc16706be34a5e7324d60601c3fce5574a096a2d95f773d1a52d038b870c0515b690931b842;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb324f3a3fa18949e217916138e1d1053efe32b0c7413d7008f080889862a60703f4038a16cfc49fb72bab5d1c1f379286971823641ad3ae835fc4f041ac54743ea739c5a444be3fd82113fc1cbb28f017251c91838e026473374fb24172ab4ee134a97581963762a31b15760d1d6e1c8;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb362c9efcac02862a0880773b071eb4c850937dd2a38d14bf58284bef6c785cea57a347e7e4c229a19ccd6390f79ca229470e65d66d798ba94be019bd83d8a2488978ed87e37d4deed09afa85acea253f3e2640fdc881c10e437a82ddb964208e703495d14eed7546491c516f573f6d52;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcbffe36aa6bd99444a6042c9adbf77716e39c81a9a2b23546e8dfc5ac076839c1f742a30a9b47d7324d45802d87249d478131da455d68894c0d140ff6edc6e4028115a110d08421fc07f27d4d4a27b61deefe9dc7e3d6f45950fd5dacfa4e6a26b77e1a14193ef866d0a3531381a1d45b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h784e86a884156c635869d83b9c8e858d74d7fc57a58162f3492324719c923537068bd8e4389dd5d3560ee717842b725d8f2c77ea6052a60d3f76381f476890265b67d251e2529c261aaf1935dc0174e3a3750888266244a50cb5974c0282e4c7acf06e1cd1c553cca7d7210b3194f6971;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d8c86caddf5622c335434a4137edb618c78c1373c78aca765afe32a4f957f1c795ebb17e8d6b1f666ec83d4f3824815b654ad1527c4b4518d55c763312c2cf4c228b1d1c4d4fda842cca125febf9a2c968e32b0571c9506141fea0e6321521c5d9538a943a7cd9e148383aca8cb704b5;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5adde1ffed9ffe595e4b4f103a2ddc8b49a2b09bd0461d00499259463ad5f1d0df7e1b7c71001ea92439a989d9335fde25db63ba9488783ffb9ac4aec7ed16c9dbadd22b61748ee414e4c2a335e7a3db41550be54d71e4ff5b1d104992d5b4f020cb4ddc2d7f2a8088a7c1cd54bb57a1d;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd25eb8433d7f7c480d2b3802738a4d25d49988d65d392f70094c58a06330e9d143e3fcedc80235ffac2e51655ebb97e5fc45634d1f3a1b3a78cb7aff057a632103e380f5fc195c096b113806360ea50ae11be5aac997af6bb4e0144eae25a71f9b27993044f3280948151e0693dd07b8a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25ddd7643e8da0b59f456a4a24414cf3c1ee1cc0cdfd1f59b51bdb71f8be22452252b1737a4b03760a37a37a38680ae4092bf971316c3cdbf27b72e717a04f9f23d1e7991ee38e5307a6d110d4cc0c0f50fa09ba9865b74a34c7cd834bb4af04f3389b31cc64ea8966add59b28e4f6dd9;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc16bb0c7d8d05330ecb51187c96cd72cb2336c9ab8c50fcca588cbf14c256602116b50b909d21e8234b2d5aa138e731c5f577ac4c20fc2427a2676e6b540f2b2e4b20be2f2f806bfc2242bdd34eb137f1f7bd342c3e2f255020b2cfbaba6d32d1ae5ea9acc137938d3227ee2d1ff80907;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc2539ba749cc48f6e9fc97fad0bd1c29e753427915ba4c58bc8da4422358d19b4062611309930dc0f36f6ab8f3adaa57022a6390ddcabb7639942c55e9f13ec6f388edde77fe9366becdb7694f9a8113331ccb4ab9fca73c906e38ba55c258e46e8f4d6ad438cf4f4d6e1ec881b7575b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45370834e6c91cb3c5e8c6a3fad330f7cadcf52d635752d9629e3237657de30befe8975d688740157bdbccff926e660cb7c4b44be3d77c0ea69dc46e7091e27660f22f10aff0327ed91eb08eed4f4e6277d9c6eeda0e88152575a2d44300051afc3cbccfa98ff47c2e3b372c3a95ac76a;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57e2fea210a71aa018a9f3809871786222876f087f6a1c5d12328d1e435c78dd2ee676c08ad1d8d0aa201e1e66749a97e9e07fd6609a127d593b401d9641fccb0d3ab227b23c6728cf460090e0f0155d06a706843b7c85bd97d9c1912628774ddaecaaf0d9a9ff99ec393ca7cca4e62f7;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34c0f287ddb21ef22814157a31fe1da7689f3cf20f97ee57303249b40b9e1f86603f4a570c60ae176e425cf92687ec2d8d60a5cf93254f07f39bc3ce7e125d115f1c5d4d1f636d658256ebfd9608983cffe60391ac8545ac98c55128b7eb36a3d0f2865ee74959e511a8f2ca4fb358112;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h288f3d55e9689b33cb1c4124e9d0586af16cd7e1a758448e0c856718c55b44ed9ba90003e77ad0abb7dec156d0de5c6f4cd34fc94ba241801d087a054e65ca6a5b065d58076f90df1331e9d816c58e1b8a7b47cc756918ba980c4cde15f945190a3333e6da10c77c57723de83a7c4f915;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc232cd491836a5dc951e308726312515ee13dbd08d6d2c1fb36072445e68f1ecae6c47cfb640e8b68897a2d548d8ebd80d11eafef960dc861b3b3d848a992d044524df9eb961411ed96d1194da8e499feb24604c942524686d56d39172b1d102d84f76774ee9e5137c3b910be4668ec39;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb87de2bdbfbcf2beb600651d547c6eb63920aec7da8bc2f6277c30f8a85aa215ab2557b671cc3b4a4c04778dcc2aed18ac7844a9fdafc83daec252e4152c89810bb7ad8a609455ea75469dfaafaabf655c05d3f894dcbd8d7bca69bee6ac7bf8019f30b24e824dd8964c60f38c2955e77;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he141922566943e003bf8a2f6c32c6eb75105ed071c1471a93ed5b472be2b1e6e9c45ba8270073db7917ca5859fcda848ed6dcb934dd00263f5749ca77181ae7ef87b00b02a22a35a5b41d8d8b97d9e0c3ac55e668260829ded33c18b290a30e75d133f14260a6b181fb238e8388834055;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd648b54f18dead493bc598c1a31653e42c2d6820013be278e6c3b67785d7f8d1b835d720c35b4fefab8711599c2636ead9039b2e4b31505a0f603aa5fdd3cf214dbd2620c968a52a5242aef43b64543bffbced906b49705298c0d69a8a6068551af1602a2888f0ff46e6000c27ea4d51b;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5306710f1c6fb7bbe444c2e3b5339230868b02f48d4c66b851941cfc3e6453470e8b050889a78e39abd901b93f83379b276cfe8304407ebadbabac0ac2a2845f26e650727ecb166e9cbbf3c67049740a464c6b79f9530ca6a3f3ddc9d047173b17c52dc322e4f81239d8d3a9f0759f9c;
        #1
        {src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47631440fcdcffae4811e92eeb069616b87c342854ad41154fc9e92cebeaf15a4932b7c3434c76d1ea0d38958a489097086a60a90a6ecc79e2d92d1cef61e1a5ece3acc1a8df2b9cf6321b6767753b4e3891b009119b766ad501d0bba08d38cb30e287b2265f396933a0867609e384a55;
        #1
        $finish();
    end
endmodule
