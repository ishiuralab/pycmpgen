module testbench();
    reg [0:0] src0;
    reg [1:0] src1;
    reg [2:0] src2;
    reg [3:0] src3;
    reg [4:0] src4;
    reg [5:0] src5;
    reg [6:0] src6;
    reg [7:0] src7;
    reg [6:0] src8;
    reg [5:0] src9;
    reg [4:0] src10;
    reg [3:0] src11;
    reg [2:0] src12;
    reg [1:0] src13;
    reg [0:0] src14;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [15:0] srcsum;
    wire [15:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15));
    assign srcsum = ((src0[0])<<0) + ((src1[0] + src1[1])<<1) + ((src2[0] + src2[1] + src2[2])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3])<<11) + ((src12[0] + src12[1] + src12[2])<<12) + ((src13[0] + src13[1])<<13) + ((src14[0])<<14);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffffffffffffffff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd1a8cbacb4d9884;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa844873ec6a3e46;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66912c9b5b2a5ebe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3eab07482d360c55;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6cab8351ae321207;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea4cc910fabaadc0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20d952857d73bd50;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d550b4f087c9a79;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h741aac82f0f4c70b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6eceb965c9563762;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h604cae877e7cad08;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a8b3e178dc723a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c7dd3e4d697be7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ac945eca525279c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e2e741e1df90f1b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9990d801c1dd534e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6810fabd4c14029;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6440fba65b986b33;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a856bc8420fc03a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h325320b07a69069d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h60ff85ace930c7fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4d2a977be38da7c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9e68c3152713d1b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ccbd069b3055709;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9190b856a338cc83;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57a91c955c908299;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7e797cd926d6cbb3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9fc911e1fede22ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9f518d6e63e8639;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8980b69603f5562d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2514bc6b156c5fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b1d5fa944b6b3d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8109d527a854912a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d8ae83754d1c706;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ae8b90ab6cbbf9e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfaaf6557f278accb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9801b36e7b3562da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a5f78600341eaf3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h919aa97442be4e52;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1008ed632c3624d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6f8930a3b71f013;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce63d8afeb16510b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfde28b61ae79999a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha375221178a7bfa2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56024e1841a59755;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ee03f551dbb74b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h26f3810a68dc843;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c72736489cafde9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h88aa5c75d1b2c527;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc466377f33ef7557;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4725d0d73b0cb89a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4504f010a0277535;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73e36325f4d55b5a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e6cd233ed7e83b7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9271f57ab11a04a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ffa2fb9ff1d5708;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc21711e7f9fc41ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e80a7c683367479;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha11038c790cc2942;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5b52f63a620155e1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d1c0cb04bf222bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h90fb2854da86c7b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h88639e5f90556f26;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h327ad82f710094a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc69263ab32feff7f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2151437826db5356;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d501249c7344f5f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h391a953ee76e6664;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8228b59f422c385b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a47a88120e5592b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc401ae826e1f006c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6399bd88a814a544;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b0064da20df1277;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h35dbaefb511292fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd15046c029c6892b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4fda454fc7f5a4b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb083894ae501793f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd1de030674e96b62;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h87e50e5c8047354a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he387e0c81e8c5414;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ae5d2b8e171e8b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h54f39bf30269ce4a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h631f315efe026407;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc02943e988d83fd9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h76f9a2d3325fd9fc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5101bb47795c18cb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcae03562e00c09f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdedd943dd897ffff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h845330d09d418bc4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28056623a842a43c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9644d42b157d368d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29a37d08ec50ab7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55159c6c9ede6070;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h680ed65dc8df5528;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had76f21f78094e9f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99fd6d63800654b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde5ebc16df4da619;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78605c4870842cc9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25d56ff333cc3c77;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha72d82c0a67e21ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he703cc212776f2b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a18cae0ff8f3752;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec620eec7e56ba66;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea7dd648e9ad1b90;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6be899e371a72495;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b5db5ab4aa013a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa8acdb2076f32f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc25b170caf78c05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h557b7842ffc07457;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdeb930c821e84d96;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9eebfec6e4d7d613;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h871f8334550dc897;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b68479ed0cca2db;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h750c331a9e3ef131;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfca13ec35135a88f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16c747e721dea23c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7882f419056cc5ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c440a432db5547e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h430583f0f60ca500;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ae554cdc25da37b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf69d42f77b90c4b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he75ee94acb141d02;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6bf3417fc6f9bf68;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99dccdd440a33f14;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c1fd0bfb66455d9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7efd4ed41f8cb5d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e4ebddef82f3ae5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25fdb81fe289e219;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he57f05c2ea4cfe9e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6551c93505874252;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h562afd1c53147dd1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b28c355db303fab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h39635da0064a6a93;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ec78f8189e91fe2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f9b8e59f7f67f24;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h486de09d0e4a3ccf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdca1fbf7f7eb658e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f0eb77a33fb29e1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d4b44fdbb79518f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40f505c04f0fb6cf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h984d6848b782a969;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h533d6d8812ce8b5a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h232b814de476711e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf67e5d6740beaf1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he2171e62d57f74e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ad65488763e0edf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hadd1f23e8ed1950c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he568be4b1c7fdc06;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he547887adb6a41ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h47a1544c57ec902d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2c78071e4993c2d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33b00dc97af6773a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33d9c8c9e3e7b604;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h611b3ea4c500568b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha32cbf7ecfebdc22;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53e316d5fdf6ac8a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3aa0f8d7f1de362f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9eeb950b3f55f872;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92bf22c60db9c421;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5397920b0839cf26;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1da65ec22b5fa397;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91e1c5094addb510;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb4fc7846e4e890d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfadbb29cbae9c7e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee60aebb6fd87af;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he582442b1fc90ead;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb90346e3714903a6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2416c48b9deada3e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf51961cdf46737;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68090bff5102bc6a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92bb5738b3a4a01c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6830806ef74d08e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5fc9b3eb0743e6af;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73b2ce6cb316c479;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7cad2513dec6781f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h814f55f9e97a5a13;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27558de4a2165832;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41c55cb9422b9a12;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1eeca9398c05f81;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc81d7d8569e03063;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf7c4070d8f0673f3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70553e43c96528d9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61693b623159dd4f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca31ac17cb9017ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h499e588ff150450c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc54a5c24132d5f39;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbac2156d289cf955;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0e03c75e213b25f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c597bf0c746ff2a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6fb62dcdcb06389a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h594fc4b0c76a031e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef9e4cf1f6fdb54;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he90f7e2b202e74d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e15cb8f51ffe38;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h702abd646728623d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d2438ab89bb67dd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9cdf596ddabdafa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbb6262c7947517a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf8fc724f70a1a3a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h74567b585f20a78c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h350dcc25a3ef11ee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29ce72f053d06834;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a6dc0dad3677236;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hecda5ee5894f986e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf92b9d7a9785380b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9743b761429aa0ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcfaf97dfa7be13eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd8648b6df397e4ee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd27f5a65c856763c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4487df3f22fac033;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8bb4415ea994d392;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80ff2877f12048c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h351fc39ad8ddc3d9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40fd9724da43d398;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85cade712c5c16f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f45bd58e5774ee2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b11ac02a677ccf1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2121ffe7ace4ca29;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28d6f3e3f001a0db;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78059eabe03bf22b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a8bedc4b5f657bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h26b772feadd29dd2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7e5582e3ba7be6d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b09b2942366bbd8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91c6940106a842d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7b5fe21799004051;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9382ba69f5bae330;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe64b6729379b2b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd79b285c2899707;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2316d40afd71c5a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec331a1aac098607;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hff71c6e32354eb02;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ac37cc0ab1f1973;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h212338bf9490b992;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d5c7d623f8eed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4fee87b0c63dd454;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44ea3a5d51b8a3b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2d098b72230a70c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd57debe863095c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55df49438f049714;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha876624fd848d048;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3a325b5a3566e6e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c819a7429317df0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6afe5703ead8e276;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha2118f817bf148ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a1fc54d8c783eca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41e279975c3cc05e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb7a158618d0d4a7e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9a4890010ca389ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he948eaa1afaf3ac7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5a27ecc91dbb4ce4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha27ef1a3e24549ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h593bee5254d55a78;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2db15698acd5db3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2afe5d0c155b939f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h64608a2d34b6f013;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc747de0390f112c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b8249ae3569355a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he61c1f326fe716a6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h71cd87d4d74a3db8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hadee5ea71b0c620c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h21edd40bbf5e3da6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2153812625b42144;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4904e7515e61d838;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27e5d518e70d376;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f8d6b6377bfe39d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc26e910350a0cfe4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61106a550ccf5a1c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf87ad908bf4d0b0e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heccd1d1c3b8a5ec7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc3c3bb5b204800b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d515b1a7eb26ebf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6af7be79fffc375d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h680ff74d9419e53b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0c048faec9229e3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h565aa0a484e88311;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he386f787023cfa29;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ee5d52991e256bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d45ba42e4f8e4fd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c625b5efb54174f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h922fd4fbb954b88f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h833a841b63d9b392;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb58507dbfea1a073;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f4b4a86e250b7cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ab477987ed12e15;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcc07bbd86913de0d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha58fcb297c76ad28;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4716c434294da92b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ac5a9482f6a23dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58a58a63d863812e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25df4813b1ffa3cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93774fe424b68fa9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd03d9da42d95931e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe11edbb73145309;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78a8e4a7f78de7d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h524a3c3b331891ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0549746d02cc75e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f5a5f32b2cf2012;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b08ec2ab36a3830;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7829e25dcadd66a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h438d103434fac4c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9df8afffec324ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1651d6dc615f827;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h13e14297c228cfa6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5fd10e3784612791;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48ba944c36338957;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ad34da4d244b3f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha50e7309ace0a365;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d045b2b27c1896e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd977e33789802fa6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb278f7abef21e3f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf60a972a72629ab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h55584c4df81e809f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85b9ac232da3cc52;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5c1bfc2521d8dfc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3e0233a17995b39;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha1c3536a41cc4c02;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8901e2cf332c296;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ec5b5d267ef8ba4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5d7731b0d66cfb3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h66abc3aea2ebb530;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h986506376b6b6285;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ba06a345117b198;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d82b91bafab37ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'headaf4bee64a1e17;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha93d8d4ea8572c72;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he056bed06d98d114;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h220edcb58bab9cd8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3ca578bf23f5f2d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61876f1d93e09a63;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f885623c4bdb38c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h86ee423ffcadb547;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha8b1e27c1c204ebf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h636896a2b83d8436;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbca157461f158ded;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h856224191d4e8cd3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdda85f477fb63e75;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc90952b6feddb3a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b27985658e9fb6f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c7ab01e5345e20a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h71e684effc2bf1d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd685adda2d556655;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd96dc9233eb95b84;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd5ea43fe8a06bd34;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf111d457a165d44e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94d1dd7f1248643f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd46473995ede1c00;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda82aa90b3c8af3d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbcf18b3035e22b24;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4cd72f472b93b371;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h732ba94b469f1dcd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62cf6862c737c926;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h406d1dd7e14095a6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7946b20ffe157562;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ec75b42e9ae2908;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdab431e8ccfcf2a3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59ed1411f0ae434;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ad5db368286a995;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca10c4fe25c656b1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h63f1707cebd2b1c9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc21968848c114cc2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4e9d4811bb2ae237;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h381947f9301143f3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h60be92a320fdaadb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3aef70d5e2130432;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h304e537f7de436a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he2c1bca977b632fd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ff3ad0f57dbd9b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b0727c23d471ecc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5fe64ddbd9f56f61;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h22428b78a04d760b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hedcff1988258605b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c9f086f8f909d43;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd95bea73935285db;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c60b3ad26236085;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9db83c14f5aeb8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2cd4fff84ace0a96;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h443df24a26b6ed52;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hedf93900f97f18c2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcbd625075827524b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1cae7dc2b19fdab2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81f4789b1462222f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48b4156ab75487dc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb248b90371246819;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2986b83eeb7e4838;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he12bdb2ae7987c38;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hddac6d626b23ae74;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee2bfc144868fc07;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h65c10254eb881caa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f3fecf45249d81a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6bf75ed5f36b7e51;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h603985c630ec0f41;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1915a1c2ff108166;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8e6d41a0fa39adb2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6018013ff81cb2d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha53a2ac6e9489e5e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he396669c1519436d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d13d82689387458;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b44dced3f35bd4b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf519043e84496de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h58b33b7685a110eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hda10b060d53e5bb3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4bca875413ec3078;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99e809524e98b152;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b3e4cc9f4165e31;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a23cd8a88c1d37d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd40bf52342f3a4c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha255f566ad061c0b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b7af400d7a1c6b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5d630c946b1b50b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf5bf113352f09754;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8501607858756ab1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5c43d322347d1bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h104f137cab4318a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77514ed5358278e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef37a794cfa96065;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb8195ddd8a2d8498;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3ed9e9e9102536b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99519901659c4526;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2fcf77f4873ccea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ddf063de56e5389;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h341361f8d8b17062;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2234a299983bcc9c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8201b84e747c5f43;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf39d29702b81fdbf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9090b1e624bb5405;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43a19e789c476f7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2a012352f4dba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2556b7b05fe6329;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha35c341a7aaa12bb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc723573c2359a6be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he588958815ba251e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43fd7fdc95878419;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he61567333e721610;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4517903b02ddcbc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he2236666ca2b5b5f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h30cc4c98c33df3b8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h431248cd02e2bd8a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3e819b7f20aeb0d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc24757bc5fba2bbe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb6a9592b598e3011;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd29dd8779c05a597;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f2d2cafdc03da6d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h385a01095cf113f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9081da3bac7d0aa3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9be7bdcbe36efdd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2e0d3e22c9cfb4bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf26bb9fc14c0fbbf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33de64ddb14a5d10;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6293582b93fad50;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3cdd8f52ff200c10;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe4986d5b4dbca6d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8061f85384b556c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h282d713b2b8bef14;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h767210fbcdfca2e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h672225e476927d92;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53185cc800477b53;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h175f89cde05f86e1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ae6061e8247562f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1db0381ae817e9be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h79292404be4bfad2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb76b2fe89df5a7b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h73d99aed0c8715f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h29ea52598acd28cb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbbb663f8aa96d3d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25df3a11d2b4116e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbefd6ca52d5e98da;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2123bd0de43c90f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h841856aa91b46631;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd4f4b4d3c01cf4d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h89bcfc766098fda6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b0db1d57c81d365;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4926d243a427c20d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hadef83e59d97073a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h154725366697f719;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h381624f05f8d34d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h32e756b711b02a46;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h995297a009956e7d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9ad4182a4947b4e0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9fd8d7111ddb5f17;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48a2d847cc23db8d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc376b4e6b370a890;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e7ae79cdca5fe24;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7ab53c5e782872d7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92ddb839892b37a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb2d79e7a7f3068d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf518625f5fa6bffa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc073ca835f31ce7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6a9cb6690f5b6f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h13c3a9cdf72fc334;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h351e98034059c9ce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2dcad89f42e32653;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc31cd35116695a7b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd58a05f0a401621a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1af63cfc61f7df3d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc5adde6066c1b64;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h26a729d76b1102f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf2fbbf798c36607c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'habe2da374e40ccc5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5df24fffc983b7ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfbc8201ad735d473;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27b3b49b6bf79ca8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5bbe64712c838a7e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h751e86368959632b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2f827563fac2c06c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae2c87d2ce3d2cae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h48cbbe43fa9743ca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ea5d10b7485e804;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ce54cfadb79a7e5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5fc225e10d1e934c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc352583d729458ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdec12808866483cd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57a832838b218ccf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb04d7b14699582f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa0c39e1b26a3dff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc9baf7458b20b0ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8817a841eedbb07b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f4a62d73f92cdb9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9368bfef2c50f905;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf70daf5b3f359253;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f22963301064e7a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h82a022fea1509d01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5ab2d553d262e2f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h906c2313c14b6e01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40af6d99c71bf3eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d01b78d01db0192;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h85ef6e9caec8ee90;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbe9b2facfc35ac9f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h909a840066f46033;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd820ffd86580316e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb28973953d4a8895;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc52ae698ac5fe371;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9723b537edfa86f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha10c98433b52d35a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb01cd0ee0aebb43;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b9b043fd9e0e9ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31c4ac189e24e029;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h237f74df32a9f0fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e6e14d6550003e9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4998af184eb94c05;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h33984873818a8a86;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h54e8c9b2c14620a1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha758b18674797fef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb04036d500a00c6c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd57f8841779d576;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he38874adef92638d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hddcc0428ac07c635;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1272f6b665a98268;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca13cd0cd5c667bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd517739f2d7808e7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hceacddfcdc5d164;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b9d330dd036bacc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h996681bca3248b29;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa99ebf6d23acc3b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfbd043b319de015c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h25454ea355688c37;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7409c12fbb29a81c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b011788b115fbfb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd73bea348f156fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2835afdb24d2cbb3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h132a824c0b285c68;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8cba16a15b6d59e2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a012977bc439f06;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd25867f255621ec0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefa18865a6514a50;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heee6b9797ca7c774;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h704157e05fa6e686;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5ffbb1c8851fcc77;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf363e39aa234c3a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb53fb25825ac1c93;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc52e60cad3879c3f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f33eb7ca7d3e7ae;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfd7d55fde2db394d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7d92a504076834de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca0e1b46aaf76f90;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf62bc29e05376e30;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h411a1cd458405a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h225d02fc4c723d58;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70b861620818ab0a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd97ca5b1d4f359d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e2ab660c163fbcc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb370530e7747f215;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha80be3fe81a1eafd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he623d6449a3df6fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e416e7c13adc1f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9544d1acb812d8fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1c7124c8135527dd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffb21ba0c2af3bb7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffe0f1482304b5bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h421c314150d25e4e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc109b49e74330c1e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h42ee653a96d3e52a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4cb1feddad86ad8e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b496e9a9bcedf66;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72b646593346170e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc571b0d4fb609acb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd560c1c51ec2f118;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h49e349e36379b3aa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h643eeb1f252316e7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7124c34d9368ff96;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hedbe217335b7cefd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdd84658e3894ead7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1197c765da926147;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb31c9d3b9af2d3ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h372dfe30fc84124e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdc80d828dcd4b9f0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6441c2f80680ee5c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h641de19e669a82ca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa28d5e507526610;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h408e23d9c64eb46b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h81bb7f68a83abaad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h352c7bed985716ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h98ee6e2b3fae1bf4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h50eb70968495adc2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd4c6f1047307033;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a70a198c7a2c60;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27cb1a199e56ddb5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0e5c533d4f15be9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5c256626e633f19;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h45ace227bf135252;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h46c8e4524fb2c709;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a1c9583710b9908;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c7988cd4c12cf52;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c29ac681f6f5e25;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h198eb4f007fe29b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc08984acecf901b1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h53228f6c5e8d5bce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ea35a5a973aba8d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h444fa880253fb00e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heb5da06418776399;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h61c54ac6f836ccea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf95f7b5aeecf2c26;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he2ada855daa42c86;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8261d468b19e85a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h34fb536c3a23ca9d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h553db1bc691f6337;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92662d3ebbc402bb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he0c6f63c38d701ba;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd6637c771f8747f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f141293b10fe5ad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h62f78e8a8a846cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f06af1117b1b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd8ae3db492e82360;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd8c6ce70d7c77d37;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec138445d8576b2b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h903b55a73a70b39a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haa252113c28a9740;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a1309d023b08c75;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2c3b45076eed8d4d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha55e2433d9bdf07c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5cbf20bd22a2afef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc5ce39b8210ba3f3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h93765ad28cda088e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb05caf2bbb6c5d90;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc2ec5d4611e9ec46;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h70258d82564623c0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d679da3dd2806a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h888ba907cc46d019;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h65894cb2b4507cbc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6352ed9c88c4c7a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5d49fab95346a9df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hedbc1a8c5ef5104c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3181f0f9bc27a9dd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1cb78e9d170b607;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb80f9cb1bcbc3ac7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha041a049721b90a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e81e0d4e9231638;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hcf6f0094e88fc45a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h23234e401f7292d6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h576316f8a74a81d0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e3e16c539f6e806;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbaa1720f6fc9f7e6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he4f482114efef25a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8856bed3d97ede81;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h44e54ad9fa2c5028;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hebb585ec0d1b5cd4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc41467294d85410;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc618c03f603174cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ab6a08fad0188e6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h373a643b63b955f6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h339a45ccc4f2873d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8d0bfa63374f4873;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a77d1ffef1ddd7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6c38611490eb2f1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f94e5a0126a38b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2613d0aae023d20c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h63e28b957b233903;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h22a1df0093c16322;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h88eac8e0698147b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9e4cdec0b3e2486;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc4fccf9053071de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9b0bc76952ed61d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3d4a92c334f75f3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5445eaf2da4ff95f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc213eb738fecadd1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b60e1c273c8b54c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h694fbebe11aa8d9e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he7dbce88466bc9c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h643a04321ed69ee0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3d82f30c271ebe87;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbf9070b40009f11f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab9ce5459e50c09c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h805926abc467c28e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4d1e52f765fc8d08;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h465897ffa4318303;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he2faa2eef3426ef9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h15c58c865c116979;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h95bed239e27a146c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdcd6c359235c97de;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc6d69539099df053;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb816d836d3fed5a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9116cddc2c9555;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6475a71e17559d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56a1cec3dc6fecca;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4acddf8236ead015;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h40832c25aa58345b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4da90c6fe7e6d421;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h166416a78c271592;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha059e989c5612bcb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc4ee2d51ecdc2310;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha93daaa36ac185c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h28d72f552ba71ff7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h625720d8aaf26b9b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8aae6c9e39cdd96d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6cf09cf3fc6aca48;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb8bbed33f0ac5ef5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf96031358740e4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1821f8165028652b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h229ea438ed9d2984;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h88b420c594eeebbe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c9232612830949;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfac59e1cd3ce9a73;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b8523e65b7edcb3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb21acb2b2931d551;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7cb830636a579793;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hefb1ddec184f722f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec3fdd529d246694;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e2281bcdf1d5a8d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8802c54f67ea2d46;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf15d1ab2818722b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7349d4a8b7ce3275;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc47567aa23098cd7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3a2ecd6ad0fc18f4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9d9ac55d1c64cc92;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c8aa258f38d52b4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77d325291906b50f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b85fe4e68314980;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c707a764c001ae4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdfd8293f2125debb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91529ea7ebf00c15;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b7e5d8222976d7e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hab3fa874b32d5fb2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h559b1e4c84c6a0c8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h515a7b9ee874e3c6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b258784bead252b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5739d3df04e7762b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h755bc76238b3eddf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f0af9fe664a7ec9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfe78152677604a0c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha07b5b4e82c888f9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbee1fe4ab264f977;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfbe2aa3343cb8d5e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd007611ca478f114;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd92a6569a371499b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfbf22298f7dcc5d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd9b53dd2b2236312;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9b1d8b2cf3ee053a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'had86a43f6aee2489;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h51cd3798c5bb4e6f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h92f1dcb381394081;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9790ec3496a49799;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h906c3546500ca1c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5dd066e0094f28ed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h936a5e12bbd79817;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc6730c991d9ee7a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb0b4590742926b2c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h584ad9bb22a69302;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4bee28e66face07d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7f028b0e864a05ff;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha0461c0db475a92;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4b5de4b405572402;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h43acbbcdebf3e442;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf19d81e5bd8f1a93;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd80d18c7ac5340a6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h56dc0b253d9e4e25;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he82ce1614655676;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6f7cf28311c82e27;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h20f989697dee29c2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h131c4d4d6dd7d5f5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd22f97c4ddc537bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8675629c6bcdae72;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hffa34ba71326b310;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h60223ef4890426b6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c58236111f830c3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc58b3bb4303ea18b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h548810fd71b45bb9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2356038c340a45c9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4631a7c8f9163d4b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd56c583246ff411;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef23c74e9b60bcd7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb5d9545a4cfd607f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc1502bcee2244ee0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h439cd17f8bbb3cad;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc12ecf2d0d5d7ca1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ca3a67f5c9060c0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf39ce593bfee4247;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d0deac618b6112b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf362fdb51616ab94;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77886340fe711870;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he4c482defff4287f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5c4feaae62a6e61c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41c5c5943d5c0c7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he3cdcf3f61242da0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6cdecb2d2e5f30d2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h78357753d0a3ccce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1cee9d03726dc6d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h82449d92e2e926;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3efccd2e5090b5f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h17cfc7fc9565a566;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3f4b9481d5fc5646;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h690bc65365cf78a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h91a7bb32cfe7fd2e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde7856f0557007b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b86a8afc8e2a53e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5f9e5a4d2782b6d5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd0ac9a5cc644d585;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94e01ea87833e9ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb025e9e689421eaf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1e7de2dfd44df782;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h452a32ca099fe01b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9cc6c48be223b28;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7aa33fefe4d77af6;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h36abf6235cf83a86;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9e787163de2c08d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6e20a2b665ca6726;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1f5833216b2e26c5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf6243686a761047d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6ccddb91aee25b9b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb587930b8aa5be60;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4c17336ecf1701a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d5fbbc50b28ef2d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf0e5ef7184ee17bc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc56532d0bc87a714;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha4d59117cb770806;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb200444efdbd7348;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e764eaa0ba29e9d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h475d7d982b14c2f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc36ef71ee470420c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha872baf3c999b138;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a2a82bb05e3eb5a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68f1b253de7b8029;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h708f1618476450ec;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4a64573627754811;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6fbf7e0664437c0e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc59fa33a9f6f719e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h52df2f36c5ad67d7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h169c680c1816c254;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2686f510fcb51c0c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6d7e23e7e2665d2d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc43153c916ab1836;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he278762458297550;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9e13b98c599ed95;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'heeb9148e4a6439ab;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf82022ed7ff4a681;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfc92c543b2498cfc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3b93016ee019df24;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h67b1d65d78e9222e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h682f66c603507e5d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4ef870cff25e3e16;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h87e13f71ec64c225;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'haf22637bcf086427;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8188a789e6a6a581;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h84bfbf663c96bdfe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb9880f678488a745;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h76babe2c149315a0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef1c1969bcedcbcf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdcd85904a515dd4b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h417de2e21c379a26;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h211cd57250efb566;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h39ce10605c9539c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9ca88f6010a63cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8ea4630d240c48a5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb3b244a346c16713;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7850e1babf112470;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8dffd5245db543a3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6a0d44b3fcf33a9d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h59a3ad809c8fa94;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h57ad4487428ff20f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc764772e344c038c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hef4ad14252b0e946;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae0ac6804fcd3330;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h673923bf19b08e39;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbc9a01a941fe6f6a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf3f339c03d068031;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c2e61bc1d0e7a6c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8b4707e512449ef5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha54ee2ed39499d84;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h401669575de6b8df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4da1c7ba09dace52;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h77441d09f28e7987;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha55d77b78b544664;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4226f083154140c4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4215d093481b08e3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ed6b51e5e659931;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8036e407549bc2a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea0deed1b703b7a8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb53f8c4ea66e54ef;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc3ca59489a6b35ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hecde37f1ee313b2b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8de6ca56b3d1eca3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb71c5b1f1b202103;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h671580ab937ca324;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h742cd49ce7ccc173;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfda435d0eac3e459;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99f857d41a1598ea;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h653aef7873d2b236;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hd112cd65e2da4be5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha65366682d356fd9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h75ccd762b7ce22b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h140e71c0aa187da2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72b7792592e81144;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5786e7e0c46625b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf09e9b88b36f47a7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h76ed06c267246005;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h970ade90e4342136;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h31fa558971ce3958;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfa7dff79d8bdc9b5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1467190a305bb7bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfc10170d2b082a2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9f3718263c40afc7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hbd3e6c539bb9c229;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha10c1c83e0bd67b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3cd2a2338b327e4d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha9b82ff1ef231002;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72dabdd1ca3b0589;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hccd81493e36c87bd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h586cfa2b418f8d1c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h258b24950cd2601c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hde75ebdf507ab9d3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hca1fe1d9a5d55e44;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a292f03c88330b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h72306ac12f2c4e78;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4fe1cca199a1985c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf4b4add5aff4ba01;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7712b93267688ff8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6b6051ae859b9444;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hce2fe94d9f8b953d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h18b0e9e2fa1fc7af;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3027cdc73edb44b3;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8cbdf1a73e3c645d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e9d6ae56b6639fd;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfc8471252344a569;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2a6423249adb2c52;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6c23d3dd62e96dfc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb1f42a703ae63ed5;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hea51962cae1c94be;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7284b30c6a258eaf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h27baf7f2929cff33;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha3401b271d1dea15;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7a501c03fdc2a93d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdeee23c6b9d1a4eb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b9865c23450c6bf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfb5810bc0a2c4abb;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h38c7517247e1a0ee;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h16494b08af779454;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5e87a37093cc8512;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfac5163eb60b7fed;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h9102aeac56433a11;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h63d4b31a6c3517fe;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2606ea7496943be2;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h676daeed97d3dc21;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hf9e77c54c2bd01b9;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6efef77560b2b47c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h68e571318e39de1c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1ae0106bc16caee8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he9abbd4b5eb2025;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41c355ea16e55050;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h302f5a641dfad525;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hec133834949a3924;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b918b2db2be550a;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2ee57a7cdbe970d8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hfc7f3407dce53198;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h94e4dd5fe4fb5931;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hdb34394066ee9932;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b7c2e34b6a81d29;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h41457ac8b498b446;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he49e915f39dd875e;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7c6f4be06cbdb126;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h6db3a124f4fb066f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3df1a5c07d2dbe4b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h39b05a2ecc1bc897;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb37493eb4344030b;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h5eebbe9c7b764e06;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h820b5a903cc9a7f8;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h926e651fe4719845;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8bb88d717ae26ccf;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4f61020cae52931d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8c628a870b08c7d1;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hee5b751c19888821;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8f1e7d7c7ca60a4;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'ha35c366939a5579d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hae0e50ba8c86d414;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h4cef1057b4f6d5df;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he4d3f31a6a754292;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he838059a803a02fa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8bb2a3fd69c77222;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7e57c5d4dc36890f;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7cc7b5b9908fb1cc;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he37481c77273969c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1b1f658e39668487;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h99a1df1bd486ac09;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hc93b084cd796e067;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1d2a924aaa67383c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'he968a3d110e1fce;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3dee294aca7ba665;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h80f3eff0e7d4abfa;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h2b93491c15202257;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7fc2b37732d1b87c;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h535787e0155c48d;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h1fdc0c241ecb0ce7;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h3c2bbfc2b6db921;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h8758718ed11390ac;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'h7724e36bfcc822b0;
        #1
        {src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 64'hb2342ba18c913a3;
        #1
        $finish();
    end
endmodule
