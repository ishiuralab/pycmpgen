module shift_register(
        input wire clk,
        input wire src0_,
        input wire src1_,
        input wire src2_,
        input wire src3_,
        input wire src4_,
        input wire src5_,
        input wire src6_,
        input wire src7_,
        input wire src8_,
        input wire src9_,
        input wire src10_,
        input wire src11_,
        input wire src12_,
        input wire src13_,
        input wire src14_,
        input wire src15_,
        input wire src16_,
        input wire src17_,
        input wire src18_,
        input wire src19_,
        input wire src20_,
        input wire src21_,
        input wire src22_,
        input wire src23_,
        input wire src24_,
        input wire src25_,
        input wire src26_,
        input wire src27_,
        input wire src28_,
        input wire src29_,
        input wire src30_,
        input wire src31_,
        input wire src32_,
        input wire src33_,
        input wire src34_,
        input wire src35_,
        input wire src36_,
        input wire src37_,
        input wire src38_,
        input wire src39_,
        input wire src40_,
        input wire src41_,
        input wire src42_,
        input wire src43_,
        input wire src44_,
        input wire src45_,
        input wire src46_,
        input wire src47_,
        input wire src48_,
        input wire src49_,
        input wire src50_,
        input wire src51_,
        input wire src52_,
        input wire src53_,
        input wire src54_,
        input wire src55_,
        input wire src56_,
        input wire src57_,
        input wire src58_,
        input wire src59_,
        input wire src60_,
        input wire src61_,
        input wire src62_,
        input wire src63_,
        output wire [0:0] dst0,
        output wire [0:0] dst1,
        output wire [0:0] dst2,
        output wire [0:0] dst3,
        output wire [0:0] dst4,
        output wire [0:0] dst5,
        output wire [0:0] dst6,
        output wire [0:0] dst7,
        output wire [0:0] dst8,
        output wire [0:0] dst9,
        output wire [0:0] dst10,
        output wire [0:0] dst11,
        output wire [0:0] dst12,
        output wire [0:0] dst13,
        output wire [0:0] dst14,
        output wire [0:0] dst15,
        output wire [0:0] dst16,
        output wire [0:0] dst17,
        output wire [0:0] dst18,
        output wire [0:0] dst19,
        output wire [0:0] dst20,
        output wire [0:0] dst21,
        output wire [0:0] dst22,
        output wire [0:0] dst23,
        output wire [0:0] dst24,
        output wire [0:0] dst25,
        output wire [0:0] dst26,
        output wire [0:0] dst27,
        output wire [0:0] dst28,
        output wire [0:0] dst29,
        output wire [0:0] dst30,
        output wire [0:0] dst31,
        output wire [0:0] dst32,
        output wire [0:0] dst33,
        output wire [0:0] dst34,
        output wire [0:0] dst35,
        output wire [0:0] dst36,
        output wire [0:0] dst37,
        output wire [0:0] dst38,
        output wire [0:0] dst39,
        output wire [0:0] dst40,
        output wire [0:0] dst41,
        output wire [0:0] dst42,
        output wire [0:0] dst43,
        output wire [0:0] dst44,
        output wire [0:0] dst45,
        output wire [0:0] dst46,
        output wire [0:0] dst47,
        output wire [0:0] dst48,
        output wire [0:0] dst49,
        output wire [0:0] dst50,
        output wire [0:0] dst51,
        output wire [0:0] dst52,
        output wire [0:0] dst53,
        output wire [0:0] dst54,
        output wire [0:0] dst55,
        output wire [0:0] dst56,
        output wire [0:0] dst57,
        output wire [0:0] dst58,
        output wire [0:0] dst59,
        output wire [0:0] dst60,
        output wire [0:0] dst61,
        output wire [0:0] dst62,
        output wire [0:0] dst63,
        output wire [0:0] dst64,
        output wire [0:0] dst65,
        output wire [0:0] dst66,
        output wire [0:0] dst67,
        output wire [0:0] dst68);
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    reg [31:0] src16;
    reg [31:0] src17;
    reg [31:0] src18;
    reg [31:0] src19;
    reg [31:0] src20;
    reg [31:0] src21;
    reg [31:0] src22;
    reg [31:0] src23;
    reg [31:0] src24;
    reg [31:0] src25;
    reg [31:0] src26;
    reg [31:0] src27;
    reg [31:0] src28;
    reg [31:0] src29;
    reg [31:0] src30;
    reg [31:0] src31;
    reg [31:0] src32;
    reg [31:0] src33;
    reg [31:0] src34;
    reg [31:0] src35;
    reg [31:0] src36;
    reg [31:0] src37;
    reg [31:0] src38;
    reg [31:0] src39;
    reg [31:0] src40;
    reg [31:0] src41;
    reg [31:0] src42;
    reg [31:0] src43;
    reg [31:0] src44;
    reg [31:0] src45;
    reg [31:0] src46;
    reg [31:0] src47;
    reg [31:0] src48;
    reg [31:0] src49;
    reg [31:0] src50;
    reg [31:0] src51;
    reg [31:0] src52;
    reg [31:0] src53;
    reg [31:0] src54;
    reg [31:0] src55;
    reg [31:0] src56;
    reg [31:0] src57;
    reg [31:0] src58;
    reg [31:0] src59;
    reg [31:0] src60;
    reg [31:0] src61;
    reg [31:0] src62;
    reg [31:0] src63;
    compressor_CLA32_64 compressor_CLA32_64(
            .src0(src0),
            .src1(src1),
            .src2(src2),
            .src3(src3),
            .src4(src4),
            .src5(src5),
            .src6(src6),
            .src7(src7),
            .src8(src8),
            .src9(src9),
            .src10(src10),
            .src11(src11),
            .src12(src12),
            .src13(src13),
            .src14(src14),
            .src15(src15),
            .src16(src16),
            .src17(src17),
            .src18(src18),
            .src19(src19),
            .src20(src20),
            .src21(src21),
            .src22(src22),
            .src23(src23),
            .src24(src24),
            .src25(src25),
            .src26(src26),
            .src27(src27),
            .src28(src28),
            .src29(src29),
            .src30(src30),
            .src31(src31),
            .src32(src32),
            .src33(src33),
            .src34(src34),
            .src35(src35),
            .src36(src36),
            .src37(src37),
            .src38(src38),
            .src39(src39),
            .src40(src40),
            .src41(src41),
            .src42(src42),
            .src43(src43),
            .src44(src44),
            .src45(src45),
            .src46(src46),
            .src47(src47),
            .src48(src48),
            .src49(src49),
            .src50(src50),
            .src51(src51),
            .src52(src52),
            .src53(src53),
            .src54(src54),
            .src55(src55),
            .src56(src56),
            .src57(src57),
            .src58(src58),
            .src59(src59),
            .src60(src60),
            .src61(src61),
            .src62(src62),
            .src63(src63),
            .dst0(dst0),
            .dst1(dst1),
            .dst2(dst2),
            .dst3(dst3),
            .dst4(dst4),
            .dst5(dst5),
            .dst6(dst6),
            .dst7(dst7),
            .dst8(dst8),
            .dst9(dst9),
            .dst10(dst10),
            .dst11(dst11),
            .dst12(dst12),
            .dst13(dst13),
            .dst14(dst14),
            .dst15(dst15),
            .dst16(dst16),
            .dst17(dst17),
            .dst18(dst18),
            .dst19(dst19),
            .dst20(dst20),
            .dst21(dst21),
            .dst22(dst22),
            .dst23(dst23),
            .dst24(dst24),
            .dst25(dst25),
            .dst26(dst26),
            .dst27(dst27),
            .dst28(dst28),
            .dst29(dst29),
            .dst30(dst30),
            .dst31(dst31),
            .dst32(dst32),
            .dst33(dst33),
            .dst34(dst34),
            .dst35(dst35),
            .dst36(dst36),
            .dst37(dst37),
            .dst38(dst38),
            .dst39(dst39),
            .dst40(dst40),
            .dst41(dst41),
            .dst42(dst42),
            .dst43(dst43),
            .dst44(dst44),
            .dst45(dst45),
            .dst46(dst46),
            .dst47(dst47),
            .dst48(dst48),
            .dst49(dst49),
            .dst50(dst50),
            .dst51(dst51),
            .dst52(dst52),
            .dst53(dst53),
            .dst54(dst54),
            .dst55(dst55),
            .dst56(dst56),
            .dst57(dst57),
            .dst58(dst58),
            .dst59(dst59),
            .dst60(dst60),
            .dst61(dst61),
            .dst62(dst62),
            .dst63(dst63),
            .dst64(dst64),
            .dst65(dst65),
            .dst66(dst66),
            .dst67(dst67),
            .dst68(dst68));
    initial begin
        src0 <= 32'h0;
        src1 <= 32'h0;
        src2 <= 32'h0;
        src3 <= 32'h0;
        src4 <= 32'h0;
        src5 <= 32'h0;
        src6 <= 32'h0;
        src7 <= 32'h0;
        src8 <= 32'h0;
        src9 <= 32'h0;
        src10 <= 32'h0;
        src11 <= 32'h0;
        src12 <= 32'h0;
        src13 <= 32'h0;
        src14 <= 32'h0;
        src15 <= 32'h0;
        src16 <= 32'h0;
        src17 <= 32'h0;
        src18 <= 32'h0;
        src19 <= 32'h0;
        src20 <= 32'h0;
        src21 <= 32'h0;
        src22 <= 32'h0;
        src23 <= 32'h0;
        src24 <= 32'h0;
        src25 <= 32'h0;
        src26 <= 32'h0;
        src27 <= 32'h0;
        src28 <= 32'h0;
        src29 <= 32'h0;
        src30 <= 32'h0;
        src31 <= 32'h0;
        src32 <= 32'h0;
        src33 <= 32'h0;
        src34 <= 32'h0;
        src35 <= 32'h0;
        src36 <= 32'h0;
        src37 <= 32'h0;
        src38 <= 32'h0;
        src39 <= 32'h0;
        src40 <= 32'h0;
        src41 <= 32'h0;
        src42 <= 32'h0;
        src43 <= 32'h0;
        src44 <= 32'h0;
        src45 <= 32'h0;
        src46 <= 32'h0;
        src47 <= 32'h0;
        src48 <= 32'h0;
        src49 <= 32'h0;
        src50 <= 32'h0;
        src51 <= 32'h0;
        src52 <= 32'h0;
        src53 <= 32'h0;
        src54 <= 32'h0;
        src55 <= 32'h0;
        src56 <= 32'h0;
        src57 <= 32'h0;
        src58 <= 32'h0;
        src59 <= 32'h0;
        src60 <= 32'h0;
        src61 <= 32'h0;
        src62 <= 32'h0;
        src63 <= 32'h0;
    end
    always @(posedge clk) begin
        src0 <= {src0, src0_};
        src1 <= {src1, src1_};
        src2 <= {src2, src2_};
        src3 <= {src3, src3_};
        src4 <= {src4, src4_};
        src5 <= {src5, src5_};
        src6 <= {src6, src6_};
        src7 <= {src7, src7_};
        src8 <= {src8, src8_};
        src9 <= {src9, src9_};
        src10 <= {src10, src10_};
        src11 <= {src11, src11_};
        src12 <= {src12, src12_};
        src13 <= {src13, src13_};
        src14 <= {src14, src14_};
        src15 <= {src15, src15_};
        src16 <= {src16, src16_};
        src17 <= {src17, src17_};
        src18 <= {src18, src18_};
        src19 <= {src19, src19_};
        src20 <= {src20, src20_};
        src21 <= {src21, src21_};
        src22 <= {src22, src22_};
        src23 <= {src23, src23_};
        src24 <= {src24, src24_};
        src25 <= {src25, src25_};
        src26 <= {src26, src26_};
        src27 <= {src27, src27_};
        src28 <= {src28, src28_};
        src29 <= {src29, src29_};
        src30 <= {src30, src30_};
        src31 <= {src31, src31_};
        src32 <= {src32, src32_};
        src33 <= {src33, src33_};
        src34 <= {src34, src34_};
        src35 <= {src35, src35_};
        src36 <= {src36, src36_};
        src37 <= {src37, src37_};
        src38 <= {src38, src38_};
        src39 <= {src39, src39_};
        src40 <= {src40, src40_};
        src41 <= {src41, src41_};
        src42 <= {src42, src42_};
        src43 <= {src43, src43_};
        src44 <= {src44, src44_};
        src45 <= {src45, src45_};
        src46 <= {src46, src46_};
        src47 <= {src47, src47_};
        src48 <= {src48, src48_};
        src49 <= {src49, src49_};
        src50 <= {src50, src50_};
        src51 <= {src51, src51_};
        src52 <= {src52, src52_};
        src53 <= {src53, src53_};
        src54 <= {src54, src54_};
        src55 <= {src55, src55_};
        src56 <= {src56, src56_};
        src57 <= {src57, src57_};
        src58 <= {src58, src58_};
        src59 <= {src59, src59_};
        src60 <= {src60, src60_};
        src61 <= {src61, src61_};
        src62 <= {src62, src62_};
        src63 <= {src63, src63_};
    end
endmodule
module compressor_CLA32_64(
    input [31:0]src0,
    input [31:0]src1,
    input [31:0]src2,
    input [31:0]src3,
    input [31:0]src4,
    input [31:0]src5,
    input [31:0]src6,
    input [31:0]src7,
    input [31:0]src8,
    input [31:0]src9,
    input [31:0]src10,
    input [31:0]src11,
    input [31:0]src12,
    input [31:0]src13,
    input [31:0]src14,
    input [31:0]src15,
    input [31:0]src16,
    input [31:0]src17,
    input [31:0]src18,
    input [31:0]src19,
    input [31:0]src20,
    input [31:0]src21,
    input [31:0]src22,
    input [31:0]src23,
    input [31:0]src24,
    input [31:0]src25,
    input [31:0]src26,
    input [31:0]src27,
    input [31:0]src28,
    input [31:0]src29,
    input [31:0]src30,
    input [31:0]src31,
    input [31:0]src32,
    input [31:0]src33,
    input [31:0]src34,
    input [31:0]src35,
    input [31:0]src36,
    input [31:0]src37,
    input [31:0]src38,
    input [31:0]src39,
    input [31:0]src40,
    input [31:0]src41,
    input [31:0]src42,
    input [31:0]src43,
    input [31:0]src44,
    input [31:0]src45,
    input [31:0]src46,
    input [31:0]src47,
    input [31:0]src48,
    input [31:0]src49,
    input [31:0]src50,
    input [31:0]src51,
    input [31:0]src52,
    input [31:0]src53,
    input [31:0]src54,
    input [31:0]src55,
    input [31:0]src56,
    input [31:0]src57,
    input [31:0]src58,
    input [31:0]src59,
    input [31:0]src60,
    input [31:0]src61,
    input [31:0]src62,
    input [31:0]src63,
    output dst0,
    output dst1,
    output dst2,
    output dst3,
    output dst4,
    output dst5,
    output dst6,
    output dst7,
    output dst8,
    output dst9,
    output dst10,
    output dst11,
    output dst12,
    output dst13,
    output dst14,
    output dst15,
    output dst16,
    output dst17,
    output dst18,
    output dst19,
    output dst20,
    output dst21,
    output dst22,
    output dst23,
    output dst24,
    output dst25,
    output dst26,
    output dst27,
    output dst28,
    output dst29,
    output dst30,
    output dst31,
    output dst32,
    output dst33,
    output dst34,
    output dst35,
    output dst36,
    output dst37,
    output dst38,
    output dst39,
    output dst40,
    output dst41,
    output dst42,
    output dst43,
    output dst44,
    output dst45,
    output dst46,
    output dst47,
    output dst48,
    output dst49,
    output dst50,
    output dst51,
    output dst52,
    output dst53,
    output dst54,
    output dst55,
    output dst56,
    output dst57,
    output dst58,
    output dst59,
    output dst60,
    output dst61,
    output dst62,
    output dst63,
    output dst64,
    output dst65,
    output dst66,
    output dst67,
    output dst68);

    wire [1:0] comp_out0;
    wire [1:0] comp_out1;
    wire [1:0] comp_out2;
    wire [1:0] comp_out3;
    wire [1:0] comp_out4;
    wire [1:0] comp_out5;
    wire [1:0] comp_out6;
    wire [1:0] comp_out7;
    wire [1:0] comp_out8;
    wire [1:0] comp_out9;
    wire [1:0] comp_out10;
    wire [1:0] comp_out11;
    wire [1:0] comp_out12;
    wire [1:0] comp_out13;
    wire [1:0] comp_out14;
    wire [1:0] comp_out15;
    wire [1:0] comp_out16;
    wire [1:0] comp_out17;
    wire [1:0] comp_out18;
    wire [1:0] comp_out19;
    wire [1:0] comp_out20;
    wire [1:0] comp_out21;
    wire [1:0] comp_out22;
    wire [1:0] comp_out23;
    wire [1:0] comp_out24;
    wire [1:0] comp_out25;
    wire [1:0] comp_out26;
    wire [1:0] comp_out27;
    wire [1:0] comp_out28;
    wire [1:0] comp_out29;
    wire [1:0] comp_out30;
    wire [1:0] comp_out31;
    wire [1:0] comp_out32;
    wire [1:0] comp_out33;
    wire [1:0] comp_out34;
    wire [1:0] comp_out35;
    wire [1:0] comp_out36;
    wire [1:0] comp_out37;
    wire [1:0] comp_out38;
    wire [1:0] comp_out39;
    wire [1:0] comp_out40;
    wire [1:0] comp_out41;
    wire [1:0] comp_out42;
    wire [1:0] comp_out43;
    wire [1:0] comp_out44;
    wire [1:0] comp_out45;
    wire [1:0] comp_out46;
    wire [1:0] comp_out47;
    wire [1:0] comp_out48;
    wire [1:0] comp_out49;
    wire [1:0] comp_out50;
    wire [1:0] comp_out51;
    wire [1:0] comp_out52;
    wire [1:0] comp_out53;
    wire [1:0] comp_out54;
    wire [1:0] comp_out55;
    wire [1:0] comp_out56;
    wire [1:0] comp_out57;
    wire [1:0] comp_out58;
    wire [1:0] comp_out59;
    wire [1:0] comp_out60;
    wire [1:0] comp_out61;
    wire [1:0] comp_out62;
    wire [1:0] comp_out63;
    wire [1:0] comp_out64;
    wire [1:0] comp_out65;
    wire [1:0] comp_out66;
    wire [1:0] comp_out67;
    wire [0:0] comp_out68;
    compressor compressor_inst(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(comp_out0),
        .dst1(comp_out1),
        .dst2(comp_out2),
        .dst3(comp_out3),
        .dst4(comp_out4),
        .dst5(comp_out5),
        .dst6(comp_out6),
        .dst7(comp_out7),
        .dst8(comp_out8),
        .dst9(comp_out9),
        .dst10(comp_out10),
        .dst11(comp_out11),
        .dst12(comp_out12),
        .dst13(comp_out13),
        .dst14(comp_out14),
        .dst15(comp_out15),
        .dst16(comp_out16),
        .dst17(comp_out17),
        .dst18(comp_out18),
        .dst19(comp_out19),
        .dst20(comp_out20),
        .dst21(comp_out21),
        .dst22(comp_out22),
        .dst23(comp_out23),
        .dst24(comp_out24),
        .dst25(comp_out25),
        .dst26(comp_out26),
        .dst27(comp_out27),
        .dst28(comp_out28),
        .dst29(comp_out29),
        .dst30(comp_out30),
        .dst31(comp_out31),
        .dst32(comp_out32),
        .dst33(comp_out33),
        .dst34(comp_out34),
        .dst35(comp_out35),
        .dst36(comp_out36),
        .dst37(comp_out37),
        .dst38(comp_out38),
        .dst39(comp_out39),
        .dst40(comp_out40),
        .dst41(comp_out41),
        .dst42(comp_out42),
        .dst43(comp_out43),
        .dst44(comp_out44),
        .dst45(comp_out45),
        .dst46(comp_out46),
        .dst47(comp_out47),
        .dst48(comp_out48),
        .dst49(comp_out49),
        .dst50(comp_out50),
        .dst51(comp_out51),
        .dst52(comp_out52),
        .dst53(comp_out53),
        .dst54(comp_out54),
        .dst55(comp_out55),
        .dst56(comp_out56),
        .dst57(comp_out57),
        .dst58(comp_out58),
        .dst59(comp_out59),
        .dst60(comp_out60),
        .dst61(comp_out61),
        .dst62(comp_out62),
        .dst63(comp_out63),
        .dst64(comp_out64),
        .dst65(comp_out65),
        .dst66(comp_out66),
        .dst67(comp_out67),
        .dst68(comp_out68)
    );
    LookAheadCarryUnit256 LCU256(
        .src0({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out68[0], comp_out67[0], comp_out66[0], comp_out65[0], comp_out64[0], comp_out63[0], comp_out62[0], comp_out61[0], comp_out60[0], comp_out59[0], comp_out58[0], comp_out57[0], comp_out56[0], comp_out55[0], comp_out54[0], comp_out53[0], comp_out52[0], comp_out51[0], comp_out50[0], comp_out49[0], comp_out48[0], comp_out47[0], comp_out46[0], comp_out45[0], comp_out44[0], comp_out43[0], comp_out42[0], comp_out41[0], comp_out40[0], comp_out39[0], comp_out38[0], comp_out37[0], comp_out36[0], comp_out35[0], comp_out34[0], comp_out33[0], comp_out32[0], comp_out31[0], comp_out30[0], comp_out29[0], comp_out28[0], comp_out27[0], comp_out26[0], comp_out25[0], comp_out24[0], comp_out23[0], comp_out22[0], comp_out21[0], comp_out20[0], comp_out19[0], comp_out18[0], comp_out17[0], comp_out16[0], comp_out15[0], comp_out14[0], comp_out13[0], comp_out12[0], comp_out11[0], comp_out10[0], comp_out9[0], comp_out8[0], comp_out7[0], comp_out6[0], comp_out5[0], comp_out4[0], comp_out3[0], comp_out2[0], comp_out1[0], comp_out0[0]}),
        .src1({1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, 1'h0, comp_out67[1], comp_out66[1], comp_out65[1], comp_out64[1], comp_out63[1], comp_out62[1], comp_out61[1], comp_out60[1], comp_out59[1], comp_out58[1], comp_out57[1], comp_out56[1], comp_out55[1], comp_out54[1], comp_out53[1], comp_out52[1], comp_out51[1], comp_out50[1], comp_out49[1], comp_out48[1], comp_out47[1], comp_out46[1], comp_out45[1], comp_out44[1], comp_out43[1], comp_out42[1], comp_out41[1], comp_out40[1], comp_out39[1], comp_out38[1], comp_out37[1], comp_out36[1], comp_out35[1], comp_out34[1], comp_out33[1], comp_out32[1], comp_out31[1], comp_out30[1], comp_out29[1], comp_out28[1], comp_out27[1], comp_out26[1], comp_out25[1], comp_out24[1], comp_out23[1], comp_out22[1], comp_out21[1], comp_out20[1], comp_out19[1], comp_out18[1], comp_out17[1], comp_out16[1], comp_out15[1], comp_out14[1], comp_out13[1], comp_out12[1], comp_out11[1], comp_out10[1], comp_out9[1], comp_out8[1], comp_out7[1], comp_out6[1], comp_out5[1], comp_out4[1], comp_out3[1], comp_out2[1], comp_out1[1], comp_out0[1]}),
        .dst({dst68, dst67, dst66, dst65, dst64, dst63, dst62, dst61, dst60, dst59, dst58, dst57, dst56, dst55, dst54, dst53, dst52, dst51, dst50, dst49, dst48, dst47, dst46, dst45, dst44, dst43, dst42, dst41, dst40, dst39, dst38, dst37, dst36, dst35, dst34, dst33, dst32, dst31, dst30, dst29, dst28, dst27, dst26, dst25, dst24, dst23, dst22, dst21, dst20, dst19, dst18, dst17, dst16, dst15, dst14, dst13, dst12, dst11, dst10, dst9, dst8, dst7, dst6, dst5, dst4, dst3, dst2, dst1, dst0})
    );
endmodule
module compressor (
      input wire [31:0] src0,
      input wire [31:0] src1,
      input wire [31:0] src2,
      input wire [31:0] src3,
      input wire [31:0] src4,
      input wire [31:0] src5,
      input wire [31:0] src6,
      input wire [31:0] src7,
      input wire [31:0] src8,
      input wire [31:0] src9,
      input wire [31:0] src10,
      input wire [31:0] src11,
      input wire [31:0] src12,
      input wire [31:0] src13,
      input wire [31:0] src14,
      input wire [31:0] src15,
      input wire [31:0] src16,
      input wire [31:0] src17,
      input wire [31:0] src18,
      input wire [31:0] src19,
      input wire [31:0] src20,
      input wire [31:0] src21,
      input wire [31:0] src22,
      input wire [31:0] src23,
      input wire [31:0] src24,
      input wire [31:0] src25,
      input wire [31:0] src26,
      input wire [31:0] src27,
      input wire [31:0] src28,
      input wire [31:0] src29,
      input wire [31:0] src30,
      input wire [31:0] src31,
      input wire [31:0] src32,
      input wire [31:0] src33,
      input wire [31:0] src34,
      input wire [31:0] src35,
      input wire [31:0] src36,
      input wire [31:0] src37,
      input wire [31:0] src38,
      input wire [31:0] src39,
      input wire [31:0] src40,
      input wire [31:0] src41,
      input wire [31:0] src42,
      input wire [31:0] src43,
      input wire [31:0] src44,
      input wire [31:0] src45,
      input wire [31:0] src46,
      input wire [31:0] src47,
      input wire [31:0] src48,
      input wire [31:0] src49,
      input wire [31:0] src50,
      input wire [31:0] src51,
      input wire [31:0] src52,
      input wire [31:0] src53,
      input wire [31:0] src54,
      input wire [31:0] src55,
      input wire [31:0] src56,
      input wire [31:0] src57,
      input wire [31:0] src58,
      input wire [31:0] src59,
      input wire [31:0] src60,
      input wire [31:0] src61,
      input wire [31:0] src62,
      input wire [31:0] src63,
      output wire [1:0] dst0,
      output wire [1:0] dst1,
      output wire [1:0] dst2,
      output wire [1:0] dst3,
      output wire [1:0] dst4,
      output wire [1:0] dst5,
      output wire [1:0] dst6,
      output wire [1:0] dst7,
      output wire [1:0] dst8,
      output wire [1:0] dst9,
      output wire [1:0] dst10,
      output wire [1:0] dst11,
      output wire [1:0] dst12,
      output wire [1:0] dst13,
      output wire [1:0] dst14,
      output wire [1:0] dst15,
      output wire [1:0] dst16,
      output wire [1:0] dst17,
      output wire [1:0] dst18,
      output wire [1:0] dst19,
      output wire [1:0] dst20,
      output wire [1:0] dst21,
      output wire [1:0] dst22,
      output wire [1:0] dst23,
      output wire [1:0] dst24,
      output wire [1:0] dst25,
      output wire [1:0] dst26,
      output wire [1:0] dst27,
      output wire [1:0] dst28,
      output wire [1:0] dst29,
      output wire [1:0] dst30,
      output wire [1:0] dst31,
      output wire [1:0] dst32,
      output wire [1:0] dst33,
      output wire [1:0] dst34,
      output wire [1:0] dst35,
      output wire [1:0] dst36,
      output wire [1:0] dst37,
      output wire [1:0] dst38,
      output wire [1:0] dst39,
      output wire [1:0] dst40,
      output wire [1:0] dst41,
      output wire [1:0] dst42,
      output wire [1:0] dst43,
      output wire [1:0] dst44,
      output wire [1:0] dst45,
      output wire [1:0] dst46,
      output wire [1:0] dst47,
      output wire [1:0] dst48,
      output wire [1:0] dst49,
      output wire [1:0] dst50,
      output wire [1:0] dst51,
      output wire [1:0] dst52,
      output wire [1:0] dst53,
      output wire [1:0] dst54,
      output wire [1:0] dst55,
      output wire [1:0] dst56,
      output wire [1:0] dst57,
      output wire [1:0] dst58,
      output wire [1:0] dst59,
      output wire [1:0] dst60,
      output wire [1:0] dst61,
      output wire [1:0] dst62,
      output wire [1:0] dst63,
      output wire [1:0] dst64,
      output wire [1:0] dst65,
      output wire [1:0] dst66,
      output wire [1:0] dst67,
      output wire [0:0] dst68);

   wire [31:0] stage0_0;
   wire [31:0] stage0_1;
   wire [31:0] stage0_2;
   wire [31:0] stage0_3;
   wire [31:0] stage0_4;
   wire [31:0] stage0_5;
   wire [31:0] stage0_6;
   wire [31:0] stage0_7;
   wire [31:0] stage0_8;
   wire [31:0] stage0_9;
   wire [31:0] stage0_10;
   wire [31:0] stage0_11;
   wire [31:0] stage0_12;
   wire [31:0] stage0_13;
   wire [31:0] stage0_14;
   wire [31:0] stage0_15;
   wire [31:0] stage0_16;
   wire [31:0] stage0_17;
   wire [31:0] stage0_18;
   wire [31:0] stage0_19;
   wire [31:0] stage0_20;
   wire [31:0] stage0_21;
   wire [31:0] stage0_22;
   wire [31:0] stage0_23;
   wire [31:0] stage0_24;
   wire [31:0] stage0_25;
   wire [31:0] stage0_26;
   wire [31:0] stage0_27;
   wire [31:0] stage0_28;
   wire [31:0] stage0_29;
   wire [31:0] stage0_30;
   wire [31:0] stage0_31;
   wire [31:0] stage0_32;
   wire [31:0] stage0_33;
   wire [31:0] stage0_34;
   wire [31:0] stage0_35;
   wire [31:0] stage0_36;
   wire [31:0] stage0_37;
   wire [31:0] stage0_38;
   wire [31:0] stage0_39;
   wire [31:0] stage0_40;
   wire [31:0] stage0_41;
   wire [31:0] stage0_42;
   wire [31:0] stage0_43;
   wire [31:0] stage0_44;
   wire [31:0] stage0_45;
   wire [31:0] stage0_46;
   wire [31:0] stage0_47;
   wire [31:0] stage0_48;
   wire [31:0] stage0_49;
   wire [31:0] stage0_50;
   wire [31:0] stage0_51;
   wire [31:0] stage0_52;
   wire [31:0] stage0_53;
   wire [31:0] stage0_54;
   wire [31:0] stage0_55;
   wire [31:0] stage0_56;
   wire [31:0] stage0_57;
   wire [31:0] stage0_58;
   wire [31:0] stage0_59;
   wire [31:0] stage0_60;
   wire [31:0] stage0_61;
   wire [31:0] stage0_62;
   wire [31:0] stage0_63;
   wire [10:0] stage1_0;
   wire [7:0] stage1_1;
   wire [24:0] stage1_2;
   wire [16:0] stage1_3;
   wire [29:0] stage1_4;
   wire [13:0] stage1_5;
   wire [28:0] stage1_6;
   wire [8:0] stage1_7;
   wire [18:0] stage1_8;
   wire [15:0] stage1_9;
   wire [17:0] stage1_10;
   wire [16:0] stage1_11;
   wire [18:0] stage1_12;
   wire [13:0] stage1_13;
   wire [16:0] stage1_14;
   wire [12:0] stage1_15;
   wire [30:0] stage1_16;
   wire [21:0] stage1_17;
   wire [10:0] stage1_18;
   wire [18:0] stage1_19;
   wire [11:0] stage1_20;
   wire [17:0] stage1_21;
   wire [13:0] stage1_22;
   wire [17:0] stage1_23;
   wire [11:0] stage1_24;
   wire [17:0] stage1_25;
   wire [16:0] stage1_26;
   wire [10:0] stage1_27;
   wire [15:0] stage1_28;
   wire [17:0] stage1_29;
   wire [10:0] stage1_30;
   wire [16:0] stage1_31;
   wire [24:0] stage1_32;
   wire [18:0] stage1_33;
   wire [20:0] stage1_34;
   wire [12:0] stage1_35;
   wire [12:0] stage1_36;
   wire [13:0] stage1_37;
   wire [17:0] stage1_38;
   wire [14:0] stage1_39;
   wire [15:0] stage1_40;
   wire [19:0] stage1_41;
   wire [12:0] stage1_42;
   wire [13:0] stage1_43;
   wire [13:0] stage1_44;
   wire [24:0] stage1_45;
   wire [11:0] stage1_46;
   wire [17:0] stage1_47;
   wire [19:0] stage1_48;
   wire [19:0] stage1_49;
   wire [11:0] stage1_50;
   wire [20:0] stage1_51;
   wire [11:0] stage1_52;
   wire [22:0] stage1_53;
   wire [9:0] stage1_54;
   wire [29:0] stage1_55;
   wire [14:0] stage1_56;
   wire [16:0] stage1_57;
   wire [13:0] stage1_58;
   wire [23:0] stage1_59;
   wire [12:0] stage1_60;
   wire [12:0] stage1_61;
   wire [16:0] stage1_62;
   wire [10:0] stage1_63;
   wire [8:0] stage1_64;
   wire [4:0] stage1_65;
   wire [10:0] stage2_0;
   wire [2:0] stage2_1;
   wire [8:0] stage2_2;
   wire [8:0] stage2_3;
   wire [6:0] stage2_4;
   wire [9:0] stage2_5;
   wire [17:0] stage2_6;
   wire [5:0] stage2_7;
   wire [5:0] stage2_8;
   wire [9:0] stage2_9;
   wire [7:0] stage2_10;
   wire [5:0] stage2_11;
   wire [5:0] stage2_12;
   wire [8:0] stage2_13;
   wire [11:0] stage2_14;
   wire [4:0] stage2_15;
   wire [11:0] stage2_16;
   wire [11:0] stage2_17;
   wire [7:0] stage2_18;
   wire [5:0] stage2_19;
   wire [7:0] stage2_20;
   wire [6:0] stage2_21;
   wire [9:0] stage2_22;
   wire [5:0] stage2_23;
   wire [7:0] stage2_24;
   wire [5:0] stage2_25;
   wire [5:0] stage2_26;
   wire [6:0] stage2_27;
   wire [8:0] stage2_28;
   wire [5:0] stage2_29;
   wire [5:0] stage2_30;
   wire [8:0] stage2_31;
   wire [7:0] stage2_32;
   wire [16:0] stage2_33;
   wire [6:0] stage2_34;
   wire [5:0] stage2_35;
   wire [7:0] stage2_36;
   wire [13:0] stage2_37;
   wire [4:0] stage2_38;
   wire [6:0] stage2_39;
   wire [5:0] stage2_40;
   wire [6:0] stage2_41;
   wire [10:0] stage2_42;
   wire [6:0] stage2_43;
   wire [17:0] stage2_44;
   wire [4:0] stage2_45;
   wire [7:0] stage2_46;
   wire [9:0] stage2_47;
   wire [6:0] stage2_48;
   wire [11:0] stage2_49;
   wire [6:0] stage2_50;
   wire [5:0] stage2_51;
   wire [5:0] stage2_52;
   wire [10:0] stage2_53;
   wire [6:0] stage2_54;
   wire [6:0] stage2_55;
   wire [9:0] stage2_56;
   wire [8:0] stage2_57;
   wire [5:0] stage2_58;
   wire [11:0] stage2_59;
   wire [6:0] stage2_60;
   wire [6:0] stage2_61;
   wire [5:0] stage2_62;
   wire [9:0] stage2_63;
   wire [4:0] stage2_64;
   wire [7:0] stage2_65;
   wire [0:0] stage2_66;
   wire [1:0] stage3_0;
   wire [1:0] stage3_1;
   wire [3:0] stage3_2;
   wire [4:0] stage3_3;
   wire [4:0] stage3_4;
   wire [2:0] stage3_5;
   wire [5:0] stage3_6;
   wire [4:0] stage3_7;
   wire [2:0] stage3_8;
   wire [3:0] stage3_9;
   wire [5:0] stage3_10;
   wire [1:0] stage3_11;
   wire [1:0] stage3_12;
   wire [4:0] stage3_13;
   wire [3:0] stage3_14;
   wire [3:0] stage3_15;
   wire [2:0] stage3_16;
   wire [3:0] stage3_17;
   wire [5:0] stage3_18;
   wire [2:0] stage3_19;
   wire [4:0] stage3_20;
   wire [2:0] stage3_21;
   wire [4:0] stage3_22;
   wire [2:0] stage3_23;
   wire [4:0] stage3_24;
   wire [1:0] stage3_25;
   wire [1:0] stage3_26;
   wire [4:0] stage3_27;
   wire [4:0] stage3_28;
   wire [1:0] stage3_29;
   wire [1:0] stage3_30;
   wire [3:0] stage3_31;
   wire [3:0] stage3_32;
   wire [3:0] stage3_33;
   wire [3:0] stage3_34;
   wire [3:0] stage3_35;
   wire [3:0] stage3_36;
   wire [3:0] stage3_37;
   wire [3:0] stage3_38;
   wire [3:0] stage3_39;
   wire [1:0] stage3_40;
   wire [2:0] stage3_41;
   wire [4:0] stage3_42;
   wire [3:0] stage3_43;
   wire [3:0] stage3_44;
   wire [3:0] stage3_45;
   wire [5:0] stage3_46;
   wire [4:0] stage3_47;
   wire [2:0] stage3_48;
   wire [2:0] stage3_49;
   wire [5:0] stage3_50;
   wire [3:0] stage3_51;
   wire [2:0] stage3_52;
   wire [2:0] stage3_53;
   wire [5:0] stage3_54;
   wire [2:0] stage3_55;
   wire [5:0] stage3_56;
   wire [2:0] stage3_57;
   wire [3:0] stage3_58;
   wire [5:0] stage3_59;
   wire [3:0] stage3_60;
   wire [2:0] stage3_61;
   wire [5:0] stage3_62;
   wire [2:0] stage3_63;
   wire [5:0] stage3_64;
   wire [3:0] stage3_65;
   wire [1:0] stage3_66;
   wire [0:0] stage3_67;
   wire [1:0] stage4_0;
   wire [1:0] stage4_1;
   wire [1:0] stage4_2;
   wire [1:0] stage4_3;
   wire [1:0] stage4_4;
   wire [1:0] stage4_5;
   wire [1:0] stage4_6;
   wire [1:0] stage4_7;
   wire [1:0] stage4_8;
   wire [1:0] stage4_9;
   wire [1:0] stage4_10;
   wire [1:0] stage4_11;
   wire [1:0] stage4_12;
   wire [1:0] stage4_13;
   wire [1:0] stage4_14;
   wire [1:0] stage4_15;
   wire [1:0] stage4_16;
   wire [1:0] stage4_17;
   wire [1:0] stage4_18;
   wire [1:0] stage4_19;
   wire [1:0] stage4_20;
   wire [1:0] stage4_21;
   wire [1:0] stage4_22;
   wire [1:0] stage4_23;
   wire [1:0] stage4_24;
   wire [1:0] stage4_25;
   wire [1:0] stage4_26;
   wire [1:0] stage4_27;
   wire [1:0] stage4_28;
   wire [1:0] stage4_29;
   wire [1:0] stage4_30;
   wire [1:0] stage4_31;
   wire [1:0] stage4_32;
   wire [1:0] stage4_33;
   wire [1:0] stage4_34;
   wire [1:0] stage4_35;
   wire [1:0] stage4_36;
   wire [1:0] stage4_37;
   wire [1:0] stage4_38;
   wire [1:0] stage4_39;
   wire [1:0] stage4_40;
   wire [1:0] stage4_41;
   wire [1:0] stage4_42;
   wire [1:0] stage4_43;
   wire [1:0] stage4_44;
   wire [1:0] stage4_45;
   wire [1:0] stage4_46;
   wire [1:0] stage4_47;
   wire [1:0] stage4_48;
   wire [1:0] stage4_49;
   wire [1:0] stage4_50;
   wire [1:0] stage4_51;
   wire [1:0] stage4_52;
   wire [1:0] stage4_53;
   wire [1:0] stage4_54;
   wire [1:0] stage4_55;
   wire [1:0] stage4_56;
   wire [1:0] stage4_57;
   wire [1:0] stage4_58;
   wire [1:0] stage4_59;
   wire [1:0] stage4_60;
   wire [1:0] stage4_61;
   wire [1:0] stage4_62;
   wire [1:0] stage4_63;
   wire [1:0] stage4_64;
   wire [1:0] stage4_65;
   wire [1:0] stage4_66;
   wire [1:0] stage4_67;
   wire [0:0] stage4_68;

   assign stage0_0 = src0;
   assign stage0_1 = src1;
   assign stage0_2 = src2;
   assign stage0_3 = src3;
   assign stage0_4 = src4;
   assign stage0_5 = src5;
   assign stage0_6 = src6;
   assign stage0_7 = src7;
   assign stage0_8 = src8;
   assign stage0_9 = src9;
   assign stage0_10 = src10;
   assign stage0_11 = src11;
   assign stage0_12 = src12;
   assign stage0_13 = src13;
   assign stage0_14 = src14;
   assign stage0_15 = src15;
   assign stage0_16 = src16;
   assign stage0_17 = src17;
   assign stage0_18 = src18;
   assign stage0_19 = src19;
   assign stage0_20 = src20;
   assign stage0_21 = src21;
   assign stage0_22 = src22;
   assign stage0_23 = src23;
   assign stage0_24 = src24;
   assign stage0_25 = src25;
   assign stage0_26 = src26;
   assign stage0_27 = src27;
   assign stage0_28 = src28;
   assign stage0_29 = src29;
   assign stage0_30 = src30;
   assign stage0_31 = src31;
   assign stage0_32 = src32;
   assign stage0_33 = src33;
   assign stage0_34 = src34;
   assign stage0_35 = src35;
   assign stage0_36 = src36;
   assign stage0_37 = src37;
   assign stage0_38 = src38;
   assign stage0_39 = src39;
   assign stage0_40 = src40;
   assign stage0_41 = src41;
   assign stage0_42 = src42;
   assign stage0_43 = src43;
   assign stage0_44 = src44;
   assign stage0_45 = src45;
   assign stage0_46 = src46;
   assign stage0_47 = src47;
   assign stage0_48 = src48;
   assign stage0_49 = src49;
   assign stage0_50 = src50;
   assign stage0_51 = src51;
   assign stage0_52 = src52;
   assign stage0_53 = src53;
   assign stage0_54 = src54;
   assign stage0_55 = src55;
   assign stage0_56 = src56;
   assign stage0_57 = src57;
   assign stage0_58 = src58;
   assign stage0_59 = src59;
   assign stage0_60 = src60;
   assign stage0_61 = src61;
   assign stage0_62 = src62;
   assign stage0_63 = src63;
   assign dst0 = stage4_0;
   assign dst1 = stage4_1;
   assign dst2 = stage4_2;
   assign dst3 = stage4_3;
   assign dst4 = stage4_4;
   assign dst5 = stage4_5;
   assign dst6 = stage4_6;
   assign dst7 = stage4_7;
   assign dst8 = stage4_8;
   assign dst9 = stage4_9;
   assign dst10 = stage4_10;
   assign dst11 = stage4_11;
   assign dst12 = stage4_12;
   assign dst13 = stage4_13;
   assign dst14 = stage4_14;
   assign dst15 = stage4_15;
   assign dst16 = stage4_16;
   assign dst17 = stage4_17;
   assign dst18 = stage4_18;
   assign dst19 = stage4_19;
   assign dst20 = stage4_20;
   assign dst21 = stage4_21;
   assign dst22 = stage4_22;
   assign dst23 = stage4_23;
   assign dst24 = stage4_24;
   assign dst25 = stage4_25;
   assign dst26 = stage4_26;
   assign dst27 = stage4_27;
   assign dst28 = stage4_28;
   assign dst29 = stage4_29;
   assign dst30 = stage4_30;
   assign dst31 = stage4_31;
   assign dst32 = stage4_32;
   assign dst33 = stage4_33;
   assign dst34 = stage4_34;
   assign dst35 = stage4_35;
   assign dst36 = stage4_36;
   assign dst37 = stage4_37;
   assign dst38 = stage4_38;
   assign dst39 = stage4_39;
   assign dst40 = stage4_40;
   assign dst41 = stage4_41;
   assign dst42 = stage4_42;
   assign dst43 = stage4_43;
   assign dst44 = stage4_44;
   assign dst45 = stage4_45;
   assign dst46 = stage4_46;
   assign dst47 = stage4_47;
   assign dst48 = stage4_48;
   assign dst49 = stage4_49;
   assign dst50 = stage4_50;
   assign dst51 = stage4_51;
   assign dst52 = stage4_52;
   assign dst53 = stage4_53;
   assign dst54 = stage4_54;
   assign dst55 = stage4_55;
   assign dst56 = stage4_56;
   assign dst57 = stage4_57;
   assign dst58 = stage4_58;
   assign dst59 = stage4_59;
   assign dst60 = stage4_60;
   assign dst61 = stage4_61;
   assign dst62 = stage4_62;
   assign dst63 = stage4_63;
   assign dst64 = stage4_64;
   assign dst65 = stage4_65;
   assign dst66 = stage4_66;
   assign dst67 = stage4_67;
   assign dst68 = stage4_68;

   gpc2116_5 gpc0 (
      {stage0_0[0], stage0_0[1], stage0_0[2], stage0_0[3], stage0_0[4], stage0_0[5]},
      {stage0_1[0]},
      {stage0_2[0]},
      {stage0_3[0], stage0_3[1]},
      {stage1_4[0],stage1_3[0],stage1_2[0],stage1_1[0],stage1_0[0]}
   );
   gpc2116_5 gpc1 (
      {stage0_0[6], stage0_0[7], stage0_0[8], stage0_0[9], stage0_0[10], stage0_0[11]},
      {stage0_1[1]},
      {stage0_2[1]},
      {stage0_3[2], stage0_3[3]},
      {stage1_4[1],stage1_3[1],stage1_2[1],stage1_1[1],stage1_0[1]}
   );
   gpc1163_5 gpc2 (
      {stage0_0[12], stage0_0[13], stage0_0[14]},
      {stage0_1[2], stage0_1[3], stage0_1[4], stage0_1[5], stage0_1[6], stage0_1[7]},
      {stage0_2[2]},
      {stage0_3[4]},
      {stage1_4[2],stage1_3[2],stage1_2[2],stage1_1[2],stage1_0[2]}
   );
   gpc1163_5 gpc3 (
      {stage0_0[15], stage0_0[16], stage0_0[17]},
      {stage0_1[8], stage0_1[9], stage0_1[10], stage0_1[11], stage0_1[12], stage0_1[13]},
      {stage0_2[3]},
      {stage0_3[5]},
      {stage1_4[3],stage1_3[3],stage1_2[3],stage1_1[3],stage1_0[3]}
   );
   gpc1163_5 gpc4 (
      {stage0_0[18], stage0_0[19], stage0_0[20]},
      {stage0_1[14], stage0_1[15], stage0_1[16], stage0_1[17], stage0_1[18], stage0_1[19]},
      {stage0_2[4]},
      {stage0_3[6]},
      {stage1_4[4],stage1_3[4],stage1_2[4],stage1_1[4],stage1_0[4]}
   );
   gpc606_5 gpc5 (
      {stage0_0[21], stage0_0[22], stage0_0[23], stage0_0[24], stage0_0[25], stage0_0[26]},
      {stage0_2[5], stage0_2[6], stage0_2[7], stage0_2[8], stage0_2[9], stage0_2[10]},
      {stage1_4[5],stage1_3[5],stage1_2[5],stage1_1[5],stage1_0[5]}
   );
   gpc606_5 gpc6 (
      {stage0_1[20], stage0_1[21], stage0_1[22], stage0_1[23], stage0_1[24], stage0_1[25]},
      {stage0_3[7], stage0_3[8], stage0_3[9], stage0_3[10], stage0_3[11], stage0_3[12]},
      {stage1_5[0],stage1_4[6],stage1_3[6],stage1_2[6],stage1_1[6]}
   );
   gpc606_5 gpc7 (
      {stage0_1[26], stage0_1[27], stage0_1[28], stage0_1[29], stage0_1[30], stage0_1[31]},
      {stage0_3[13], stage0_3[14], stage0_3[15], stage0_3[16], stage0_3[17], stage0_3[18]},
      {stage1_5[1],stage1_4[7],stage1_3[7],stage1_2[7],stage1_1[7]}
   );
   gpc615_5 gpc8 (
      {stage0_2[11], stage0_2[12], stage0_2[13], stage0_2[14], stage0_2[15]},
      {stage0_3[19]},
      {stage0_4[0], stage0_4[1], stage0_4[2], stage0_4[3], stage0_4[4], stage0_4[5]},
      {stage1_6[0],stage1_5[2],stage1_4[8],stage1_3[8],stage1_2[8]}
   );
   gpc615_5 gpc9 (
      {stage0_3[20], stage0_3[21], stage0_3[22], stage0_3[23], stage0_3[24]},
      {stage0_4[6]},
      {stage0_5[0], stage0_5[1], stage0_5[2], stage0_5[3], stage0_5[4], stage0_5[5]},
      {stage1_7[0],stage1_6[1],stage1_5[3],stage1_4[9],stage1_3[9]}
   );
   gpc606_5 gpc10 (
      {stage0_4[7], stage0_4[8], stage0_4[9], stage0_4[10], stage0_4[11], stage0_4[12]},
      {stage0_6[0], stage0_6[1], stage0_6[2], stage0_6[3], stage0_6[4], stage0_6[5]},
      {stage1_8[0],stage1_7[1],stage1_6[2],stage1_5[4],stage1_4[10]}
   );
   gpc1343_5 gpc11 (
      {stage0_5[6], stage0_5[7], stage0_5[8]},
      {stage0_6[6], stage0_6[7], stage0_6[8], stage0_6[9]},
      {stage0_7[0], stage0_7[1], stage0_7[2]},
      {stage0_8[0]},
      {stage1_9[0],stage1_8[1],stage1_7[2],stage1_6[3],stage1_5[5]}
   );
   gpc606_5 gpc12 (
      {stage0_5[9], stage0_5[10], stage0_5[11], stage0_5[12], stage0_5[13], stage0_5[14]},
      {stage0_7[3], stage0_7[4], stage0_7[5], stage0_7[6], stage0_7[7], stage0_7[8]},
      {stage1_9[1],stage1_8[2],stage1_7[3],stage1_6[4],stage1_5[6]}
   );
   gpc606_5 gpc13 (
      {stage0_5[15], stage0_5[16], stage0_5[17], stage0_5[18], stage0_5[19], stage0_5[20]},
      {stage0_7[9], stage0_7[10], stage0_7[11], stage0_7[12], stage0_7[13], stage0_7[14]},
      {stage1_9[2],stage1_8[3],stage1_7[4],stage1_6[5],stage1_5[7]}
   );
   gpc606_5 gpc14 (
      {stage0_5[21], stage0_5[22], stage0_5[23], stage0_5[24], stage0_5[25], stage0_5[26]},
      {stage0_7[15], stage0_7[16], stage0_7[17], stage0_7[18], stage0_7[19], stage0_7[20]},
      {stage1_9[3],stage1_8[4],stage1_7[5],stage1_6[6],stage1_5[8]}
   );
   gpc615_5 gpc15 (
      {stage0_7[21], stage0_7[22], stage0_7[23], stage0_7[24], stage0_7[25]},
      {stage0_8[1]},
      {stage0_9[0], stage0_9[1], stage0_9[2], stage0_9[3], stage0_9[4], stage0_9[5]},
      {stage1_11[0],stage1_10[0],stage1_9[4],stage1_8[5],stage1_7[6]}
   );
   gpc615_5 gpc16 (
      {stage0_7[26], stage0_7[27], stage0_7[28], stage0_7[29], stage0_7[30]},
      {stage0_8[2]},
      {stage0_9[6], stage0_9[7], stage0_9[8], stage0_9[9], stage0_9[10], stage0_9[11]},
      {stage1_11[1],stage1_10[1],stage1_9[5],stage1_8[6],stage1_7[7]}
   );
   gpc2135_5 gpc17 (
      {stage0_8[3], stage0_8[4], stage0_8[5], stage0_8[6], stage0_8[7]},
      {stage0_9[12], stage0_9[13], stage0_9[14]},
      {stage0_10[0]},
      {stage0_11[0], stage0_11[1]},
      {stage1_12[0],stage1_11[2],stage1_10[2],stage1_9[6],stage1_8[7]}
   );
   gpc606_5 gpc18 (
      {stage0_8[8], stage0_8[9], stage0_8[10], stage0_8[11], stage0_8[12], stage0_8[13]},
      {stage0_10[1], stage0_10[2], stage0_10[3], stage0_10[4], stage0_10[5], stage0_10[6]},
      {stage1_12[1],stage1_11[3],stage1_10[3],stage1_9[7],stage1_8[8]}
   );
   gpc615_5 gpc19 (
      {stage0_8[14], stage0_8[15], stage0_8[16], stage0_8[17], stage0_8[18]},
      {stage0_9[15]},
      {stage0_10[7], stage0_10[8], stage0_10[9], stage0_10[10], stage0_10[11], stage0_10[12]},
      {stage1_12[2],stage1_11[4],stage1_10[4],stage1_9[8],stage1_8[9]}
   );
   gpc615_5 gpc20 (
      {stage0_8[19], stage0_8[20], stage0_8[21], stage0_8[22], stage0_8[23]},
      {stage0_9[16]},
      {stage0_10[13], stage0_10[14], stage0_10[15], stage0_10[16], stage0_10[17], stage0_10[18]},
      {stage1_12[3],stage1_11[5],stage1_10[5],stage1_9[9],stage1_8[10]}
   );
   gpc606_5 gpc21 (
      {stage0_9[17], stage0_9[18], stage0_9[19], stage0_9[20], stage0_9[21], stage0_9[22]},
      {stage0_11[2], stage0_11[3], stage0_11[4], stage0_11[5], stage0_11[6], stage0_11[7]},
      {stage1_13[0],stage1_12[4],stage1_11[6],stage1_10[6],stage1_9[10]}
   );
   gpc623_5 gpc22 (
      {stage0_9[23], stage0_9[24], stage0_9[25]},
      {stage0_10[19], stage0_10[20]},
      {stage0_11[8], stage0_11[9], stage0_11[10], stage0_11[11], stage0_11[12], stage0_11[13]},
      {stage1_13[1],stage1_12[5],stage1_11[7],stage1_10[7],stage1_9[11]}
   );
   gpc623_5 gpc23 (
      {stage0_9[26], stage0_9[27], stage0_9[28]},
      {stage0_10[21], stage0_10[22]},
      {stage0_11[14], stage0_11[15], stage0_11[16], stage0_11[17], stage0_11[18], stage0_11[19]},
      {stage1_13[2],stage1_12[6],stage1_11[8],stage1_10[8],stage1_9[12]}
   );
   gpc615_5 gpc24 (
      {stage0_11[20], stage0_11[21], stage0_11[22], stage0_11[23], stage0_11[24]},
      {stage0_12[0]},
      {stage0_13[0], stage0_13[1], stage0_13[2], stage0_13[3], stage0_13[4], stage0_13[5]},
      {stage1_15[0],stage1_14[0],stage1_13[3],stage1_12[7],stage1_11[9]}
   );
   gpc606_5 gpc25 (
      {stage0_12[1], stage0_12[2], stage0_12[3], stage0_12[4], stage0_12[5], stage0_12[6]},
      {stage0_14[0], stage0_14[1], stage0_14[2], stage0_14[3], stage0_14[4], stage0_14[5]},
      {stage1_16[0],stage1_15[1],stage1_14[1],stage1_13[4],stage1_12[8]}
   );
   gpc606_5 gpc26 (
      {stage0_12[7], stage0_12[8], stage0_12[9], stage0_12[10], stage0_12[11], stage0_12[12]},
      {stage0_14[6], stage0_14[7], stage0_14[8], stage0_14[9], stage0_14[10], stage0_14[11]},
      {stage1_16[1],stage1_15[2],stage1_14[2],stage1_13[5],stage1_12[9]}
   );
   gpc606_5 gpc27 (
      {stage0_12[13], stage0_12[14], stage0_12[15], stage0_12[16], stage0_12[17], stage0_12[18]},
      {stage0_14[12], stage0_14[13], stage0_14[14], stage0_14[15], stage0_14[16], stage0_14[17]},
      {stage1_16[2],stage1_15[3],stage1_14[3],stage1_13[6],stage1_12[10]}
   );
   gpc606_5 gpc28 (
      {stage0_12[19], stage0_12[20], stage0_12[21], stage0_12[22], stage0_12[23], stage0_12[24]},
      {stage0_14[18], stage0_14[19], stage0_14[20], stage0_14[21], stage0_14[22], stage0_14[23]},
      {stage1_16[3],stage1_15[4],stage1_14[4],stage1_13[7],stage1_12[11]}
   );
   gpc606_5 gpc29 (
      {stage0_13[6], stage0_13[7], stage0_13[8], stage0_13[9], stage0_13[10], stage0_13[11]},
      {stage0_15[0], stage0_15[1], stage0_15[2], stage0_15[3], stage0_15[4], stage0_15[5]},
      {stage1_17[0],stage1_16[4],stage1_15[5],stage1_14[5],stage1_13[8]}
   );
   gpc606_5 gpc30 (
      {stage0_13[12], stage0_13[13], stage0_13[14], stage0_13[15], stage0_13[16], stage0_13[17]},
      {stage0_15[6], stage0_15[7], stage0_15[8], stage0_15[9], stage0_15[10], stage0_15[11]},
      {stage1_17[1],stage1_16[5],stage1_15[6],stage1_14[6],stage1_13[9]}
   );
   gpc606_5 gpc31 (
      {stage0_13[18], stage0_13[19], stage0_13[20], stage0_13[21], stage0_13[22], stage0_13[23]},
      {stage0_15[12], stage0_15[13], stage0_15[14], stage0_15[15], stage0_15[16], stage0_15[17]},
      {stage1_17[2],stage1_16[6],stage1_15[7],stage1_14[7],stage1_13[10]}
   );
   gpc606_5 gpc32 (
      {stage0_13[24], stage0_13[25], stage0_13[26], stage0_13[27], stage0_13[28], stage0_13[29]},
      {stage0_15[18], stage0_15[19], stage0_15[20], stage0_15[21], stage0_15[22], stage0_15[23]},
      {stage1_17[3],stage1_16[7],stage1_15[8],stage1_14[8],stage1_13[11]}
   );
   gpc615_5 gpc33 (
      {stage0_15[24], stage0_15[25], stage0_15[26], stage0_15[27], stage0_15[28]},
      {stage0_16[0]},
      {stage0_17[0], stage0_17[1], stage0_17[2], stage0_17[3], stage0_17[4], stage0_17[5]},
      {stage1_19[0],stage1_18[0],stage1_17[4],stage1_16[8],stage1_15[9]}
   );
   gpc606_5 gpc34 (
      {stage0_16[1], stage0_16[2], stage0_16[3], stage0_16[4], stage0_16[5], stage0_16[6]},
      {stage0_18[0], stage0_18[1], stage0_18[2], stage0_18[3], stage0_18[4], stage0_18[5]},
      {stage1_20[0],stage1_19[1],stage1_18[1],stage1_17[5],stage1_16[9]}
   );
   gpc615_5 gpc35 (
      {stage0_16[7], stage0_16[8], stage0_16[9], stage0_16[10], stage0_16[11]},
      {stage0_17[6]},
      {stage0_18[6], stage0_18[7], stage0_18[8], stage0_18[9], stage0_18[10], stage0_18[11]},
      {stage1_20[1],stage1_19[2],stage1_18[2],stage1_17[6],stage1_16[10]}
   );
   gpc606_5 gpc36 (
      {stage0_17[7], stage0_17[8], stage0_17[9], stage0_17[10], stage0_17[11], stage0_17[12]},
      {stage0_19[0], stage0_19[1], stage0_19[2], stage0_19[3], stage0_19[4], stage0_19[5]},
      {stage1_21[0],stage1_20[2],stage1_19[3],stage1_18[3],stage1_17[7]}
   );
   gpc606_5 gpc37 (
      {stage0_17[13], stage0_17[14], stage0_17[15], stage0_17[16], stage0_17[17], stage0_17[18]},
      {stage0_19[6], stage0_19[7], stage0_19[8], stage0_19[9], stage0_19[10], stage0_19[11]},
      {stage1_21[1],stage1_20[3],stage1_19[4],stage1_18[4],stage1_17[8]}
   );
   gpc1406_5 gpc38 (
      {stage0_18[12], stage0_18[13], stage0_18[14], stage0_18[15], stage0_18[16], stage0_18[17]},
      {stage0_20[0], stage0_20[1], stage0_20[2], stage0_20[3]},
      {stage0_21[0]},
      {stage1_22[0],stage1_21[2],stage1_20[4],stage1_19[5],stage1_18[5]}
   );
   gpc1406_5 gpc39 (
      {stage0_18[18], stage0_18[19], stage0_18[20], stage0_18[21], stage0_18[22], stage0_18[23]},
      {stage0_20[4], stage0_20[5], stage0_20[6], stage0_20[7]},
      {stage0_21[1]},
      {stage1_22[1],stage1_21[3],stage1_20[5],stage1_19[6],stage1_18[6]}
   );
   gpc615_5 gpc40 (
      {stage0_18[24], stage0_18[25], stage0_18[26], stage0_18[27], stage0_18[28]},
      {stage0_19[12]},
      {stage0_20[8], stage0_20[9], stage0_20[10], stage0_20[11], stage0_20[12], stage0_20[13]},
      {stage1_22[2],stage1_21[4],stage1_20[6],stage1_19[7],stage1_18[7]}
   );
   gpc615_5 gpc41 (
      {stage0_19[13], stage0_19[14], stage0_19[15], stage0_19[16], stage0_19[17]},
      {stage0_20[14]},
      {stage0_21[2], stage0_21[3], stage0_21[4], stage0_21[5], stage0_21[6], stage0_21[7]},
      {stage1_23[0],stage1_22[3],stage1_21[5],stage1_20[7],stage1_19[8]}
   );
   gpc615_5 gpc42 (
      {stage0_19[18], stage0_19[19], stage0_19[20], stage0_19[21], stage0_19[22]},
      {stage0_20[15]},
      {stage0_21[8], stage0_21[9], stage0_21[10], stage0_21[11], stage0_21[12], stage0_21[13]},
      {stage1_23[1],stage1_22[4],stage1_21[6],stage1_20[8],stage1_19[9]}
   );
   gpc606_5 gpc43 (
      {stage0_20[16], stage0_20[17], stage0_20[18], stage0_20[19], stage0_20[20], stage0_20[21]},
      {stage0_22[0], stage0_22[1], stage0_22[2], stage0_22[3], stage0_22[4], stage0_22[5]},
      {stage1_24[0],stage1_23[2],stage1_22[5],stage1_21[7],stage1_20[9]}
   );
   gpc606_5 gpc44 (
      {stage0_20[22], stage0_20[23], stage0_20[24], stage0_20[25], stage0_20[26], stage0_20[27]},
      {stage0_22[6], stage0_22[7], stage0_22[8], stage0_22[9], stage0_22[10], stage0_22[11]},
      {stage1_24[1],stage1_23[3],stage1_22[6],stage1_21[8],stage1_20[10]}
   );
   gpc606_5 gpc45 (
      {stage0_20[28], stage0_20[29], stage0_20[30], stage0_20[31], 1'b0, 1'b0},
      {stage0_22[12], stage0_22[13], stage0_22[14], stage0_22[15], stage0_22[16], stage0_22[17]},
      {stage1_24[2],stage1_23[4],stage1_22[7],stage1_21[9],stage1_20[11]}
   );
   gpc606_5 gpc46 (
      {stage0_21[14], stage0_21[15], stage0_21[16], stage0_21[17], stage0_21[18], stage0_21[19]},
      {stage0_23[0], stage0_23[1], stage0_23[2], stage0_23[3], stage0_23[4], stage0_23[5]},
      {stage1_25[0],stage1_24[3],stage1_23[5],stage1_22[8],stage1_21[10]}
   );
   gpc606_5 gpc47 (
      {stage0_21[20], stage0_21[21], stage0_21[22], stage0_21[23], stage0_21[24], stage0_21[25]},
      {stage0_23[6], stage0_23[7], stage0_23[8], stage0_23[9], stage0_23[10], stage0_23[11]},
      {stage1_25[1],stage1_24[4],stage1_23[6],stage1_22[9],stage1_21[11]}
   );
   gpc1163_5 gpc48 (
      {stage0_22[18], stage0_22[19], stage0_22[20]},
      {stage0_23[12], stage0_23[13], stage0_23[14], stage0_23[15], stage0_23[16], stage0_23[17]},
      {stage0_24[0]},
      {stage0_25[0]},
      {stage1_26[0],stage1_25[2],stage1_24[5],stage1_23[7],stage1_22[10]}
   );
   gpc615_5 gpc49 (
      {stage0_22[21], stage0_22[22], stage0_22[23], stage0_22[24], stage0_22[25]},
      {stage0_23[18]},
      {stage0_24[1], stage0_24[2], stage0_24[3], stage0_24[4], stage0_24[5], stage0_24[6]},
      {stage1_26[1],stage1_25[3],stage1_24[6],stage1_23[8],stage1_22[11]}
   );
   gpc615_5 gpc50 (
      {stage0_22[26], stage0_22[27], stage0_22[28], stage0_22[29], stage0_22[30]},
      {stage0_23[19]},
      {stage0_24[7], stage0_24[8], stage0_24[9], stage0_24[10], stage0_24[11], stage0_24[12]},
      {stage1_26[2],stage1_25[4],stage1_24[7],stage1_23[9],stage1_22[12]}
   );
   gpc615_5 gpc51 (
      {stage0_23[20], stage0_23[21], stage0_23[22], stage0_23[23], stage0_23[24]},
      {stage0_24[13]},
      {stage0_25[1], stage0_25[2], stage0_25[3], stage0_25[4], stage0_25[5], stage0_25[6]},
      {stage1_27[0],stage1_26[3],stage1_25[5],stage1_24[8],stage1_23[10]}
   );
   gpc606_5 gpc52 (
      {stage0_24[14], stage0_24[15], stage0_24[16], stage0_24[17], stage0_24[18], stage0_24[19]},
      {stage0_26[0], stage0_26[1], stage0_26[2], stage0_26[3], stage0_26[4], stage0_26[5]},
      {stage1_28[0],stage1_27[1],stage1_26[4],stage1_25[6],stage1_24[9]}
   );
   gpc606_5 gpc53 (
      {stage0_24[20], stage0_24[21], stage0_24[22], stage0_24[23], stage0_24[24], stage0_24[25]},
      {stage0_26[6], stage0_26[7], stage0_26[8], stage0_26[9], stage0_26[10], stage0_26[11]},
      {stage1_28[1],stage1_27[2],stage1_26[5],stage1_25[7],stage1_24[10]}
   );
   gpc606_5 gpc54 (
      {stage0_24[26], stage0_24[27], stage0_24[28], stage0_24[29], stage0_24[30], stage0_24[31]},
      {stage0_26[12], stage0_26[13], stage0_26[14], stage0_26[15], stage0_26[16], stage0_26[17]},
      {stage1_28[2],stage1_27[3],stage1_26[6],stage1_25[8],stage1_24[11]}
   );
   gpc615_5 gpc55 (
      {stage0_25[7], stage0_25[8], stage0_25[9], stage0_25[10], stage0_25[11]},
      {stage0_26[18]},
      {stage0_27[0], stage0_27[1], stage0_27[2], stage0_27[3], stage0_27[4], stage0_27[5]},
      {stage1_29[0],stage1_28[3],stage1_27[4],stage1_26[7],stage1_25[9]}
   );
   gpc615_5 gpc56 (
      {stage0_25[12], stage0_25[13], stage0_25[14], stage0_25[15], stage0_25[16]},
      {stage0_26[19]},
      {stage0_27[6], stage0_27[7], stage0_27[8], stage0_27[9], stage0_27[10], stage0_27[11]},
      {stage1_29[1],stage1_28[4],stage1_27[5],stage1_26[8],stage1_25[10]}
   );
   gpc615_5 gpc57 (
      {stage0_25[17], stage0_25[18], stage0_25[19], stage0_25[20], stage0_25[21]},
      {stage0_26[20]},
      {stage0_27[12], stage0_27[13], stage0_27[14], stage0_27[15], stage0_27[16], stage0_27[17]},
      {stage1_29[2],stage1_28[5],stage1_27[6],stage1_26[9],stage1_25[11]}
   );
   gpc615_5 gpc58 (
      {stage0_25[22], stage0_25[23], stage0_25[24], stage0_25[25], stage0_25[26]},
      {stage0_26[21]},
      {stage0_27[18], stage0_27[19], stage0_27[20], stage0_27[21], stage0_27[22], stage0_27[23]},
      {stage1_29[3],stage1_28[6],stage1_27[7],stage1_26[10],stage1_25[12]}
   );
   gpc615_5 gpc59 (
      {stage0_26[22], stage0_26[23], stage0_26[24], stage0_26[25], stage0_26[26]},
      {stage0_27[24]},
      {stage0_28[0], stage0_28[1], stage0_28[2], stage0_28[3], stage0_28[4], stage0_28[5]},
      {stage1_30[0],stage1_29[4],stage1_28[7],stage1_27[8],stage1_26[11]}
   );
   gpc606_5 gpc60 (
      {stage0_27[25], stage0_27[26], stage0_27[27], stage0_27[28], stage0_27[29], stage0_27[30]},
      {stage0_29[0], stage0_29[1], stage0_29[2], stage0_29[3], stage0_29[4], stage0_29[5]},
      {stage1_31[0],stage1_30[1],stage1_29[5],stage1_28[8],stage1_27[9]}
   );
   gpc606_5 gpc61 (
      {stage0_28[6], stage0_28[7], stage0_28[8], stage0_28[9], stage0_28[10], stage0_28[11]},
      {stage0_30[0], stage0_30[1], stage0_30[2], stage0_30[3], stage0_30[4], stage0_30[5]},
      {stage1_32[0],stage1_31[1],stage1_30[2],stage1_29[6],stage1_28[9]}
   );
   gpc606_5 gpc62 (
      {stage0_28[12], stage0_28[13], stage0_28[14], stage0_28[15], stage0_28[16], stage0_28[17]},
      {stage0_30[6], stage0_30[7], stage0_30[8], stage0_30[9], stage0_30[10], stage0_30[11]},
      {stage1_32[1],stage1_31[2],stage1_30[3],stage1_29[7],stage1_28[10]}
   );
   gpc606_5 gpc63 (
      {stage0_28[18], stage0_28[19], stage0_28[20], stage0_28[21], stage0_28[22], stage0_28[23]},
      {stage0_30[12], stage0_30[13], stage0_30[14], stage0_30[15], stage0_30[16], stage0_30[17]},
      {stage1_32[2],stage1_31[3],stage1_30[4],stage1_29[8],stage1_28[11]}
   );
   gpc615_5 gpc64 (
      {stage0_28[24], stage0_28[25], stage0_28[26], stage0_28[27], stage0_28[28]},
      {stage0_29[6]},
      {stage0_30[18], stage0_30[19], stage0_30[20], stage0_30[21], stage0_30[22], stage0_30[23]},
      {stage1_32[3],stage1_31[4],stage1_30[5],stage1_29[9],stage1_28[12]}
   );
   gpc606_5 gpc65 (
      {stage0_29[7], stage0_29[8], stage0_29[9], stage0_29[10], stage0_29[11], stage0_29[12]},
      {stage0_31[0], stage0_31[1], stage0_31[2], stage0_31[3], stage0_31[4], stage0_31[5]},
      {stage1_33[0],stage1_32[4],stage1_31[5],stage1_30[6],stage1_29[10]}
   );
   gpc615_5 gpc66 (
      {stage0_29[13], stage0_29[14], stage0_29[15], stage0_29[16], stage0_29[17]},
      {stage0_30[24]},
      {stage0_31[6], stage0_31[7], stage0_31[8], stage0_31[9], stage0_31[10], stage0_31[11]},
      {stage1_33[1],stage1_32[5],stage1_31[6],stage1_30[7],stage1_29[11]}
   );
   gpc615_5 gpc67 (
      {stage0_29[18], stage0_29[19], stage0_29[20], stage0_29[21], stage0_29[22]},
      {stage0_30[25]},
      {stage0_31[12], stage0_31[13], stage0_31[14], stage0_31[15], stage0_31[16], stage0_31[17]},
      {stage1_33[2],stage1_32[6],stage1_31[7],stage1_30[8],stage1_29[12]}
   );
   gpc615_5 gpc68 (
      {stage0_29[23], stage0_29[24], stage0_29[25], stage0_29[26], stage0_29[27]},
      {stage0_30[26]},
      {stage0_31[18], stage0_31[19], stage0_31[20], stage0_31[21], stage0_31[22], stage0_31[23]},
      {stage1_33[3],stage1_32[7],stage1_31[8],stage1_30[9],stage1_29[13]}
   );
   gpc615_5 gpc69 (
      {stage0_30[27], stage0_30[28], stage0_30[29], stage0_30[30], stage0_30[31]},
      {stage0_31[24]},
      {stage0_32[0], stage0_32[1], stage0_32[2], stage0_32[3], stage0_32[4], stage0_32[5]},
      {stage1_34[0],stage1_33[4],stage1_32[8],stage1_31[9],stage1_30[10]}
   );
   gpc606_5 gpc70 (
      {stage0_32[6], stage0_32[7], stage0_32[8], stage0_32[9], stage0_32[10], stage0_32[11]},
      {stage0_34[0], stage0_34[1], stage0_34[2], stage0_34[3], stage0_34[4], stage0_34[5]},
      {stage1_36[0],stage1_35[0],stage1_34[1],stage1_33[5],stage1_32[9]}
   );
   gpc606_5 gpc71 (
      {stage0_32[12], stage0_32[13], stage0_32[14], stage0_32[15], stage0_32[16], stage0_32[17]},
      {stage0_34[6], stage0_34[7], stage0_34[8], stage0_34[9], stage0_34[10], stage0_34[11]},
      {stage1_36[1],stage1_35[1],stage1_34[2],stage1_33[6],stage1_32[10]}
   );
   gpc606_5 gpc72 (
      {stage0_33[0], stage0_33[1], stage0_33[2], stage0_33[3], stage0_33[4], stage0_33[5]},
      {stage0_35[0], stage0_35[1], stage0_35[2], stage0_35[3], stage0_35[4], stage0_35[5]},
      {stage1_37[0],stage1_36[2],stage1_35[2],stage1_34[3],stage1_33[7]}
   );
   gpc606_5 gpc73 (
      {stage0_33[6], stage0_33[7], stage0_33[8], stage0_33[9], stage0_33[10], stage0_33[11]},
      {stage0_35[6], stage0_35[7], stage0_35[8], stage0_35[9], stage0_35[10], stage0_35[11]},
      {stage1_37[1],stage1_36[3],stage1_35[3],stage1_34[4],stage1_33[8]}
   );
   gpc606_5 gpc74 (
      {stage0_33[12], stage0_33[13], stage0_33[14], stage0_33[15], stage0_33[16], stage0_33[17]},
      {stage0_35[12], stage0_35[13], stage0_35[14], stage0_35[15], stage0_35[16], stage0_35[17]},
      {stage1_37[2],stage1_36[4],stage1_35[4],stage1_34[5],stage1_33[9]}
   );
   gpc606_5 gpc75 (
      {stage0_33[18], stage0_33[19], stage0_33[20], stage0_33[21], stage0_33[22], stage0_33[23]},
      {stage0_35[18], stage0_35[19], stage0_35[20], stage0_35[21], stage0_35[22], stage0_35[23]},
      {stage1_37[3],stage1_36[5],stage1_35[5],stage1_34[6],stage1_33[10]}
   );
   gpc615_5 gpc76 (
      {stage0_34[12], stage0_34[13], stage0_34[14], stage0_34[15], stage0_34[16]},
      {stage0_35[24]},
      {stage0_36[0], stage0_36[1], stage0_36[2], stage0_36[3], stage0_36[4], stage0_36[5]},
      {stage1_38[0],stage1_37[4],stage1_36[6],stage1_35[6],stage1_34[7]}
   );
   gpc623_5 gpc77 (
      {stage0_34[17], stage0_34[18], stage0_34[19]},
      {stage0_35[25], stage0_35[26]},
      {stage0_36[6], stage0_36[7], stage0_36[8], stage0_36[9], stage0_36[10], stage0_36[11]},
      {stage1_38[1],stage1_37[5],stage1_36[7],stage1_35[7],stage1_34[8]}
   );
   gpc606_5 gpc78 (
      {stage0_36[12], stage0_36[13], stage0_36[14], stage0_36[15], stage0_36[16], stage0_36[17]},
      {stage0_38[0], stage0_38[1], stage0_38[2], stage0_38[3], stage0_38[4], stage0_38[5]},
      {stage1_40[0],stage1_39[0],stage1_38[2],stage1_37[6],stage1_36[8]}
   );
   gpc606_5 gpc79 (
      {stage0_36[18], stage0_36[19], stage0_36[20], stage0_36[21], stage0_36[22], stage0_36[23]},
      {stage0_38[6], stage0_38[7], stage0_38[8], stage0_38[9], stage0_38[10], stage0_38[11]},
      {stage1_40[1],stage1_39[1],stage1_38[3],stage1_37[7],stage1_36[9]}
   );
   gpc606_5 gpc80 (
      {stage0_36[24], stage0_36[25], stage0_36[26], stage0_36[27], stage0_36[28], stage0_36[29]},
      {stage0_38[12], stage0_38[13], stage0_38[14], stage0_38[15], stage0_38[16], stage0_38[17]},
      {stage1_40[2],stage1_39[2],stage1_38[4],stage1_37[8],stage1_36[10]}
   );
   gpc117_4 gpc81 (
      {stage0_37[0], stage0_37[1], stage0_37[2], stage0_37[3], stage0_37[4], stage0_37[5], stage0_37[6]},
      {stage0_38[18]},
      {stage0_39[0]},
      {stage1_40[3],stage1_39[3],stage1_38[5],stage1_37[9]}
   );
   gpc117_4 gpc82 (
      {stage0_37[7], stage0_37[8], stage0_37[9], stage0_37[10], stage0_37[11], stage0_37[12], stage0_37[13]},
      {stage0_38[19]},
      {stage0_39[1]},
      {stage1_40[4],stage1_39[4],stage1_38[6],stage1_37[10]}
   );
   gpc606_5 gpc83 (
      {stage0_37[14], stage0_37[15], stage0_37[16], stage0_37[17], stage0_37[18], stage0_37[19]},
      {stage0_39[2], stage0_39[3], stage0_39[4], stage0_39[5], stage0_39[6], stage0_39[7]},
      {stage1_41[0],stage1_40[5],stage1_39[5],stage1_38[7],stage1_37[11]}
   );
   gpc606_5 gpc84 (
      {stage0_37[20], stage0_37[21], stage0_37[22], stage0_37[23], stage0_37[24], stage0_37[25]},
      {stage0_39[8], stage0_39[9], stage0_39[10], stage0_39[11], stage0_39[12], stage0_39[13]},
      {stage1_41[1],stage1_40[6],stage1_39[6],stage1_38[8],stage1_37[12]}
   );
   gpc606_5 gpc85 (
      {stage0_37[26], stage0_37[27], stage0_37[28], stage0_37[29], stage0_37[30], stage0_37[31]},
      {stage0_39[14], stage0_39[15], stage0_39[16], stage0_39[17], stage0_39[18], stage0_39[19]},
      {stage1_41[2],stage1_40[7],stage1_39[7],stage1_38[9],stage1_37[13]}
   );
   gpc615_5 gpc86 (
      {stage0_38[20], stage0_38[21], stage0_38[22], stage0_38[23], stage0_38[24]},
      {stage0_39[20]},
      {stage0_40[0], stage0_40[1], stage0_40[2], stage0_40[3], stage0_40[4], stage0_40[5]},
      {stage1_42[0],stage1_41[3],stage1_40[8],stage1_39[8],stage1_38[10]}
   );
   gpc606_5 gpc87 (
      {stage0_39[21], stage0_39[22], stage0_39[23], stage0_39[24], stage0_39[25], stage0_39[26]},
      {stage0_41[0], stage0_41[1], stage0_41[2], stage0_41[3], stage0_41[4], stage0_41[5]},
      {stage1_43[0],stage1_42[1],stage1_41[4],stage1_40[9],stage1_39[9]}
   );
   gpc606_5 gpc88 (
      {stage0_40[6], stage0_40[7], stage0_40[8], stage0_40[9], stage0_40[10], stage0_40[11]},
      {stage0_42[0], stage0_42[1], stage0_42[2], stage0_42[3], stage0_42[4], stage0_42[5]},
      {stage1_44[0],stage1_43[1],stage1_42[2],stage1_41[5],stage1_40[10]}
   );
   gpc606_5 gpc89 (
      {stage0_40[12], stage0_40[13], stage0_40[14], stage0_40[15], stage0_40[16], stage0_40[17]},
      {stage0_42[6], stage0_42[7], stage0_42[8], stage0_42[9], stage0_42[10], stage0_42[11]},
      {stage1_44[1],stage1_43[2],stage1_42[3],stage1_41[6],stage1_40[11]}
   );
   gpc606_5 gpc90 (
      {stage0_40[18], stage0_40[19], stage0_40[20], stage0_40[21], stage0_40[22], stage0_40[23]},
      {stage0_42[12], stage0_42[13], stage0_42[14], stage0_42[15], stage0_42[16], stage0_42[17]},
      {stage1_44[2],stage1_43[3],stage1_42[4],stage1_41[7],stage1_40[12]}
   );
   gpc606_5 gpc91 (
      {stage0_40[24], stage0_40[25], stage0_40[26], stage0_40[27], stage0_40[28], stage0_40[29]},
      {stage0_42[18], stage0_42[19], stage0_42[20], stage0_42[21], stage0_42[22], stage0_42[23]},
      {stage1_44[3],stage1_43[4],stage1_42[5],stage1_41[8],stage1_40[13]}
   );
   gpc606_5 gpc92 (
      {stage0_41[6], stage0_41[7], stage0_41[8], stage0_41[9], stage0_41[10], stage0_41[11]},
      {stage0_43[0], stage0_43[1], stage0_43[2], stage0_43[3], stage0_43[4], stage0_43[5]},
      {stage1_45[0],stage1_44[4],stage1_43[5],stage1_42[6],stage1_41[9]}
   );
   gpc606_5 gpc93 (
      {stage0_41[12], stage0_41[13], stage0_41[14], stage0_41[15], stage0_41[16], stage0_41[17]},
      {stage0_43[6], stage0_43[7], stage0_43[8], stage0_43[9], stage0_43[10], stage0_43[11]},
      {stage1_45[1],stage1_44[5],stage1_43[6],stage1_42[7],stage1_41[10]}
   );
   gpc606_5 gpc94 (
      {stage0_41[18], stage0_41[19], stage0_41[20], stage0_41[21], stage0_41[22], stage0_41[23]},
      {stage0_43[12], stage0_43[13], stage0_43[14], stage0_43[15], stage0_43[16], stage0_43[17]},
      {stage1_45[2],stage1_44[6],stage1_43[7],stage1_42[8],stage1_41[11]}
   );
   gpc615_5 gpc95 (
      {stage0_42[24], stage0_42[25], stage0_42[26], stage0_42[27], stage0_42[28]},
      {stage0_43[18]},
      {stage0_44[0], stage0_44[1], stage0_44[2], stage0_44[3], stage0_44[4], stage0_44[5]},
      {stage1_46[0],stage1_45[3],stage1_44[7],stage1_43[8],stage1_42[9]}
   );
   gpc615_5 gpc96 (
      {stage0_43[19], stage0_43[20], stage0_43[21], stage0_43[22], stage0_43[23]},
      {stage0_44[6]},
      {stage0_45[0], stage0_45[1], stage0_45[2], stage0_45[3], stage0_45[4], stage0_45[5]},
      {stage1_47[0],stage1_46[1],stage1_45[4],stage1_44[8],stage1_43[9]}
   );
   gpc615_5 gpc97 (
      {stage0_43[24], stage0_43[25], stage0_43[26], stage0_43[27], stage0_43[28]},
      {stage0_44[7]},
      {stage0_45[6], stage0_45[7], stage0_45[8], stage0_45[9], stage0_45[10], stage0_45[11]},
      {stage1_47[1],stage1_46[2],stage1_45[5],stage1_44[9],stage1_43[10]}
   );
   gpc606_5 gpc98 (
      {stage0_44[8], stage0_44[9], stage0_44[10], stage0_44[11], stage0_44[12], stage0_44[13]},
      {stage0_46[0], stage0_46[1], stage0_46[2], stage0_46[3], stage0_46[4], stage0_46[5]},
      {stage1_48[0],stage1_47[2],stage1_46[3],stage1_45[6],stage1_44[10]}
   );
   gpc606_5 gpc99 (
      {stage0_44[14], stage0_44[15], stage0_44[16], stage0_44[17], stage0_44[18], stage0_44[19]},
      {stage0_46[6], stage0_46[7], stage0_46[8], stage0_46[9], stage0_46[10], stage0_46[11]},
      {stage1_48[1],stage1_47[3],stage1_46[4],stage1_45[7],stage1_44[11]}
   );
   gpc606_5 gpc100 (
      {stage0_44[20], stage0_44[21], stage0_44[22], stage0_44[23], stage0_44[24], stage0_44[25]},
      {stage0_46[12], stage0_46[13], stage0_46[14], stage0_46[15], stage0_46[16], stage0_46[17]},
      {stage1_48[2],stage1_47[4],stage1_46[5],stage1_45[8],stage1_44[12]}
   );
   gpc606_5 gpc101 (
      {stage0_44[26], stage0_44[27], stage0_44[28], stage0_44[29], stage0_44[30], stage0_44[31]},
      {stage0_46[18], stage0_46[19], stage0_46[20], stage0_46[21], stage0_46[22], stage0_46[23]},
      {stage1_48[3],stage1_47[5],stage1_46[6],stage1_45[9],stage1_44[13]}
   );
   gpc606_5 gpc102 (
      {stage0_45[12], stage0_45[13], stage0_45[14], stage0_45[15], stage0_45[16], stage0_45[17]},
      {stage0_47[0], stage0_47[1], stage0_47[2], stage0_47[3], stage0_47[4], stage0_47[5]},
      {stage1_49[0],stage1_48[4],stage1_47[6],stage1_46[7],stage1_45[10]}
   );
   gpc615_5 gpc103 (
      {stage0_46[24], stage0_46[25], stage0_46[26], stage0_46[27], stage0_46[28]},
      {stage0_47[6]},
      {stage0_48[0], stage0_48[1], stage0_48[2], stage0_48[3], stage0_48[4], stage0_48[5]},
      {stage1_50[0],stage1_49[1],stage1_48[5],stage1_47[7],stage1_46[8]}
   );
   gpc606_5 gpc104 (
      {stage0_47[7], stage0_47[8], stage0_47[9], stage0_47[10], stage0_47[11], stage0_47[12]},
      {stage0_49[0], stage0_49[1], stage0_49[2], stage0_49[3], stage0_49[4], stage0_49[5]},
      {stage1_51[0],stage1_50[1],stage1_49[2],stage1_48[6],stage1_47[8]}
   );
   gpc606_5 gpc105 (
      {stage0_47[13], stage0_47[14], stage0_47[15], stage0_47[16], stage0_47[17], stage0_47[18]},
      {stage0_49[6], stage0_49[7], stage0_49[8], stage0_49[9], stage0_49[10], stage0_49[11]},
      {stage1_51[1],stage1_50[2],stage1_49[3],stage1_48[7],stage1_47[9]}
   );
   gpc606_5 gpc106 (
      {stage0_47[19], stage0_47[20], stage0_47[21], stage0_47[22], stage0_47[23], stage0_47[24]},
      {stage0_49[12], stage0_49[13], stage0_49[14], stage0_49[15], stage0_49[16], stage0_49[17]},
      {stage1_51[2],stage1_50[3],stage1_49[4],stage1_48[8],stage1_47[10]}
   );
   gpc606_5 gpc107 (
      {stage0_48[6], stage0_48[7], stage0_48[8], stage0_48[9], stage0_48[10], stage0_48[11]},
      {stage0_50[0], stage0_50[1], stage0_50[2], stage0_50[3], stage0_50[4], stage0_50[5]},
      {stage1_52[0],stage1_51[3],stage1_50[4],stage1_49[5],stage1_48[9]}
   );
   gpc606_5 gpc108 (
      {stage0_48[12], stage0_48[13], stage0_48[14], stage0_48[15], stage0_48[16], stage0_48[17]},
      {stage0_50[6], stage0_50[7], stage0_50[8], stage0_50[9], stage0_50[10], stage0_50[11]},
      {stage1_52[1],stage1_51[4],stage1_50[5],stage1_49[6],stage1_48[10]}
   );
   gpc606_5 gpc109 (
      {stage0_48[18], stage0_48[19], stage0_48[20], stage0_48[21], stage0_48[22], stage0_48[23]},
      {stage0_50[12], stage0_50[13], stage0_50[14], stage0_50[15], stage0_50[16], stage0_50[17]},
      {stage1_52[2],stage1_51[5],stage1_50[6],stage1_49[7],stage1_48[11]}
   );
   gpc623_5 gpc110 (
      {stage0_49[18], stage0_49[19], stage0_49[20]},
      {stage0_50[18], stage0_50[19]},
      {stage0_51[0], stage0_51[1], stage0_51[2], stage0_51[3], stage0_51[4], stage0_51[5]},
      {stage1_53[0],stage1_52[3],stage1_51[6],stage1_50[7],stage1_49[8]}
   );
   gpc615_5 gpc111 (
      {stage0_50[20], stage0_50[21], stage0_50[22], stage0_50[23], stage0_50[24]},
      {stage0_51[6]},
      {stage0_52[0], stage0_52[1], stage0_52[2], stage0_52[3], stage0_52[4], stage0_52[5]},
      {stage1_54[0],stage1_53[1],stage1_52[4],stage1_51[7],stage1_50[8]}
   );
   gpc615_5 gpc112 (
      {stage0_50[25], stage0_50[26], stage0_50[27], stage0_50[28], stage0_50[29]},
      {stage0_51[7]},
      {stage0_52[6], stage0_52[7], stage0_52[8], stage0_52[9], stage0_52[10], stage0_52[11]},
      {stage1_54[1],stage1_53[2],stage1_52[5],stage1_51[8],stage1_50[9]}
   );
   gpc615_5 gpc113 (
      {stage0_51[8], stage0_51[9], stage0_51[10], stage0_51[11], stage0_51[12]},
      {stage0_52[12]},
      {stage0_53[0], stage0_53[1], stage0_53[2], stage0_53[3], stage0_53[4], stage0_53[5]},
      {stage1_55[0],stage1_54[2],stage1_53[3],stage1_52[6],stage1_51[9]}
   );
   gpc615_5 gpc114 (
      {stage0_51[13], stage0_51[14], stage0_51[15], stage0_51[16], stage0_51[17]},
      {stage0_52[13]},
      {stage0_53[6], stage0_53[7], stage0_53[8], stage0_53[9], stage0_53[10], stage0_53[11]},
      {stage1_55[1],stage1_54[3],stage1_53[4],stage1_52[7],stage1_51[10]}
   );
   gpc615_5 gpc115 (
      {stage0_51[18], stage0_51[19], stage0_51[20], stage0_51[21], stage0_51[22]},
      {stage0_52[14]},
      {stage0_53[12], stage0_53[13], stage0_53[14], stage0_53[15], stage0_53[16], stage0_53[17]},
      {stage1_55[2],stage1_54[4],stage1_53[5],stage1_52[8],stage1_51[11]}
   );
   gpc606_5 gpc116 (
      {stage0_52[15], stage0_52[16], stage0_52[17], stage0_52[18], stage0_52[19], stage0_52[20]},
      {stage0_54[0], stage0_54[1], stage0_54[2], stage0_54[3], stage0_54[4], stage0_54[5]},
      {stage1_56[0],stage1_55[3],stage1_54[5],stage1_53[6],stage1_52[9]}
   );
   gpc606_5 gpc117 (
      {stage0_52[21], stage0_52[22], stage0_52[23], stage0_52[24], stage0_52[25], stage0_52[26]},
      {stage0_54[6], stage0_54[7], stage0_54[8], stage0_54[9], stage0_54[10], stage0_54[11]},
      {stage1_56[1],stage1_55[4],stage1_54[6],stage1_53[7],stage1_52[10]}
   );
   gpc606_5 gpc118 (
      {stage0_52[27], stage0_52[28], stage0_52[29], stage0_52[30], stage0_52[31], 1'b0},
      {stage0_54[12], stage0_54[13], stage0_54[14], stage0_54[15], stage0_54[16], stage0_54[17]},
      {stage1_56[2],stage1_55[5],stage1_54[7],stage1_53[8],stage1_52[11]}
   );
   gpc207_4 gpc119 (
      {stage0_54[18], stage0_54[19], stage0_54[20], stage0_54[21], stage0_54[22], stage0_54[23], stage0_54[24]},
      {stage0_56[0], stage0_56[1]},
      {stage1_57[0],stage1_56[3],stage1_55[6],stage1_54[8]}
   );
   gpc207_4 gpc120 (
      {stage0_54[25], stage0_54[26], stage0_54[27], stage0_54[28], stage0_54[29], stage0_54[30], stage0_54[31]},
      {stage0_56[2], stage0_56[3]},
      {stage1_57[1],stage1_56[4],stage1_55[7],stage1_54[9]}
   );
   gpc1163_5 gpc121 (
      {stage0_55[0], stage0_55[1], stage0_55[2]},
      {stage0_56[4], stage0_56[5], stage0_56[6], stage0_56[7], stage0_56[8], stage0_56[9]},
      {stage0_57[0]},
      {stage0_58[0]},
      {stage1_59[0],stage1_58[0],stage1_57[2],stage1_56[5],stage1_55[8]}
   );
   gpc615_5 gpc122 (
      {stage0_55[3], stage0_55[4], stage0_55[5], stage0_55[6], stage0_55[7]},
      {stage0_56[10]},
      {stage0_57[1], stage0_57[2], stage0_57[3], stage0_57[4], stage0_57[5], stage0_57[6]},
      {stage1_59[1],stage1_58[1],stage1_57[3],stage1_56[6],stage1_55[9]}
   );
   gpc615_5 gpc123 (
      {stage0_55[8], stage0_55[9], stage0_55[10], stage0_55[11], stage0_55[12]},
      {stage0_56[11]},
      {stage0_57[7], stage0_57[8], stage0_57[9], stage0_57[10], stage0_57[11], stage0_57[12]},
      {stage1_59[2],stage1_58[2],stage1_57[4],stage1_56[7],stage1_55[10]}
   );
   gpc606_5 gpc124 (
      {stage0_56[12], stage0_56[13], stage0_56[14], stage0_56[15], stage0_56[16], stage0_56[17]},
      {stage0_58[1], stage0_58[2], stage0_58[3], stage0_58[4], stage0_58[5], stage0_58[6]},
      {stage1_60[0],stage1_59[3],stage1_58[3],stage1_57[5],stage1_56[8]}
   );
   gpc615_5 gpc125 (
      {stage0_56[18], stage0_56[19], stage0_56[20], stage0_56[21], stage0_56[22]},
      {stage0_57[13]},
      {stage0_58[7], stage0_58[8], stage0_58[9], stage0_58[10], stage0_58[11], stage0_58[12]},
      {stage1_60[1],stage1_59[4],stage1_58[4],stage1_57[6],stage1_56[9]}
   );
   gpc615_5 gpc126 (
      {stage0_56[23], stage0_56[24], stage0_56[25], stage0_56[26], stage0_56[27]},
      {stage0_57[14]},
      {stage0_58[13], stage0_58[14], stage0_58[15], stage0_58[16], stage0_58[17], stage0_58[18]},
      {stage1_60[2],stage1_59[5],stage1_58[5],stage1_57[7],stage1_56[10]}
   );
   gpc615_5 gpc127 (
      {stage0_57[15], stage0_57[16], stage0_57[17], stage0_57[18], stage0_57[19]},
      {stage0_58[19]},
      {stage0_59[0], stage0_59[1], stage0_59[2], stage0_59[3], stage0_59[4], stage0_59[5]},
      {stage1_61[0],stage1_60[3],stage1_59[6],stage1_58[6],stage1_57[8]}
   );
   gpc615_5 gpc128 (
      {stage0_57[20], stage0_57[21], stage0_57[22], stage0_57[23], stage0_57[24]},
      {stage0_58[20]},
      {stage0_59[6], stage0_59[7], stage0_59[8], stage0_59[9], stage0_59[10], stage0_59[11]},
      {stage1_61[1],stage1_60[4],stage1_59[7],stage1_58[7],stage1_57[9]}
   );
   gpc606_5 gpc129 (
      {stage0_58[21], stage0_58[22], stage0_58[23], stage0_58[24], stage0_58[25], stage0_58[26]},
      {stage0_60[0], stage0_60[1], stage0_60[2], stage0_60[3], stage0_60[4], stage0_60[5]},
      {stage1_62[0],stage1_61[2],stage1_60[5],stage1_59[8],stage1_58[8]}
   );
   gpc606_5 gpc130 (
      {stage0_59[12], stage0_59[13], stage0_59[14], stage0_59[15], stage0_59[16], stage0_59[17]},
      {stage0_61[0], stage0_61[1], stage0_61[2], stage0_61[3], stage0_61[4], stage0_61[5]},
      {stage1_63[0],stage1_62[1],stage1_61[3],stage1_60[6],stage1_59[9]}
   );
   gpc1406_5 gpc131 (
      {stage0_60[6], stage0_60[7], stage0_60[8], stage0_60[9], stage0_60[10], stage0_60[11]},
      {stage0_62[0], stage0_62[1], stage0_62[2], stage0_62[3]},
      {stage0_63[0]},
      {stage1_64[0],stage1_63[1],stage1_62[2],stage1_61[4],stage1_60[7]}
   );
   gpc606_5 gpc132 (
      {stage0_60[12], stage0_60[13], stage0_60[14], stage0_60[15], stage0_60[16], stage0_60[17]},
      {stage0_62[4], stage0_62[5], stage0_62[6], stage0_62[7], stage0_62[8], stage0_62[9]},
      {stage1_64[1],stage1_63[2],stage1_62[3],stage1_61[5],stage1_60[8]}
   );
   gpc606_5 gpc133 (
      {stage0_60[18], stage0_60[19], stage0_60[20], stage0_60[21], stage0_60[22], stage0_60[23]},
      {stage0_62[10], stage0_62[11], stage0_62[12], stage0_62[13], stage0_62[14], stage0_62[15]},
      {stage1_64[2],stage1_63[3],stage1_62[4],stage1_61[6],stage1_60[9]}
   );
   gpc606_5 gpc134 (
      {stage0_60[24], stage0_60[25], stage0_60[26], stage0_60[27], stage0_60[28], stage0_60[29]},
      {stage0_62[16], stage0_62[17], stage0_62[18], stage0_62[19], stage0_62[20], stage0_62[21]},
      {stage1_64[3],stage1_63[4],stage1_62[5],stage1_61[7],stage1_60[10]}
   );
   gpc606_5 gpc135 (
      {stage0_61[6], stage0_61[7], stage0_61[8], stage0_61[9], stage0_61[10], stage0_61[11]},
      {stage0_63[1], stage0_63[2], stage0_63[3], stage0_63[4], stage0_63[5], stage0_63[6]},
      {stage1_65[0],stage1_64[4],stage1_63[5],stage1_62[6],stage1_61[8]}
   );
   gpc615_5 gpc136 (
      {stage0_61[12], stage0_61[13], stage0_61[14], stage0_61[15], stage0_61[16]},
      {stage0_62[22]},
      {stage0_63[7], stage0_63[8], stage0_63[9], stage0_63[10], stage0_63[11], stage0_63[12]},
      {stage1_65[1],stage1_64[5],stage1_63[6],stage1_62[7],stage1_61[9]}
   );
   gpc615_5 gpc137 (
      {stage0_61[17], stage0_61[18], stage0_61[19], stage0_61[20], stage0_61[21]},
      {stage0_62[23]},
      {stage0_63[13], stage0_63[14], stage0_63[15], stage0_63[16], stage0_63[17], stage0_63[18]},
      {stage1_65[2],stage1_64[6],stage1_63[7],stage1_62[8],stage1_61[10]}
   );
   gpc615_5 gpc138 (
      {stage0_61[22], stage0_61[23], stage0_61[24], stage0_61[25], stage0_61[26]},
      {stage0_62[24]},
      {stage0_63[19], stage0_63[20], stage0_63[21], stage0_63[22], stage0_63[23], stage0_63[24]},
      {stage1_65[3],stage1_64[7],stage1_63[8],stage1_62[9],stage1_61[11]}
   );
   gpc615_5 gpc139 (
      {stage0_61[27], stage0_61[28], stage0_61[29], stage0_61[30], stage0_61[31]},
      {stage0_62[25]},
      {stage0_63[25], stage0_63[26], stage0_63[27], stage0_63[28], stage0_63[29], stage0_63[30]},
      {stage1_65[4],stage1_64[8],stage1_63[9],stage1_62[10],stage1_61[12]}
   );
   gpc1_1 gpc140 (
      {stage0_0[27]},
      {stage1_0[6]}
   );
   gpc1_1 gpc141 (
      {stage0_0[28]},
      {stage1_0[7]}
   );
   gpc1_1 gpc142 (
      {stage0_0[29]},
      {stage1_0[8]}
   );
   gpc1_1 gpc143 (
      {stage0_0[30]},
      {stage1_0[9]}
   );
   gpc1_1 gpc144 (
      {stage0_0[31]},
      {stage1_0[10]}
   );
   gpc1_1 gpc145 (
      {stage0_2[16]},
      {stage1_2[9]}
   );
   gpc1_1 gpc146 (
      {stage0_2[17]},
      {stage1_2[10]}
   );
   gpc1_1 gpc147 (
      {stage0_2[18]},
      {stage1_2[11]}
   );
   gpc1_1 gpc148 (
      {stage0_2[19]},
      {stage1_2[12]}
   );
   gpc1_1 gpc149 (
      {stage0_2[20]},
      {stage1_2[13]}
   );
   gpc1_1 gpc150 (
      {stage0_2[21]},
      {stage1_2[14]}
   );
   gpc1_1 gpc151 (
      {stage0_2[22]},
      {stage1_2[15]}
   );
   gpc1_1 gpc152 (
      {stage0_2[23]},
      {stage1_2[16]}
   );
   gpc1_1 gpc153 (
      {stage0_2[24]},
      {stage1_2[17]}
   );
   gpc1_1 gpc154 (
      {stage0_2[25]},
      {stage1_2[18]}
   );
   gpc1_1 gpc155 (
      {stage0_2[26]},
      {stage1_2[19]}
   );
   gpc1_1 gpc156 (
      {stage0_2[27]},
      {stage1_2[20]}
   );
   gpc1_1 gpc157 (
      {stage0_2[28]},
      {stage1_2[21]}
   );
   gpc1_1 gpc158 (
      {stage0_2[29]},
      {stage1_2[22]}
   );
   gpc1_1 gpc159 (
      {stage0_2[30]},
      {stage1_2[23]}
   );
   gpc1_1 gpc160 (
      {stage0_2[31]},
      {stage1_2[24]}
   );
   gpc1_1 gpc161 (
      {stage0_3[25]},
      {stage1_3[10]}
   );
   gpc1_1 gpc162 (
      {stage0_3[26]},
      {stage1_3[11]}
   );
   gpc1_1 gpc163 (
      {stage0_3[27]},
      {stage1_3[12]}
   );
   gpc1_1 gpc164 (
      {stage0_3[28]},
      {stage1_3[13]}
   );
   gpc1_1 gpc165 (
      {stage0_3[29]},
      {stage1_3[14]}
   );
   gpc1_1 gpc166 (
      {stage0_3[30]},
      {stage1_3[15]}
   );
   gpc1_1 gpc167 (
      {stage0_3[31]},
      {stage1_3[16]}
   );
   gpc1_1 gpc168 (
      {stage0_4[13]},
      {stage1_4[11]}
   );
   gpc1_1 gpc169 (
      {stage0_4[14]},
      {stage1_4[12]}
   );
   gpc1_1 gpc170 (
      {stage0_4[15]},
      {stage1_4[13]}
   );
   gpc1_1 gpc171 (
      {stage0_4[16]},
      {stage1_4[14]}
   );
   gpc1_1 gpc172 (
      {stage0_4[17]},
      {stage1_4[15]}
   );
   gpc1_1 gpc173 (
      {stage0_4[18]},
      {stage1_4[16]}
   );
   gpc1_1 gpc174 (
      {stage0_4[19]},
      {stage1_4[17]}
   );
   gpc1_1 gpc175 (
      {stage0_4[20]},
      {stage1_4[18]}
   );
   gpc1_1 gpc176 (
      {stage0_4[21]},
      {stage1_4[19]}
   );
   gpc1_1 gpc177 (
      {stage0_4[22]},
      {stage1_4[20]}
   );
   gpc1_1 gpc178 (
      {stage0_4[23]},
      {stage1_4[21]}
   );
   gpc1_1 gpc179 (
      {stage0_4[24]},
      {stage1_4[22]}
   );
   gpc1_1 gpc180 (
      {stage0_4[25]},
      {stage1_4[23]}
   );
   gpc1_1 gpc181 (
      {stage0_4[26]},
      {stage1_4[24]}
   );
   gpc1_1 gpc182 (
      {stage0_4[27]},
      {stage1_4[25]}
   );
   gpc1_1 gpc183 (
      {stage0_4[28]},
      {stage1_4[26]}
   );
   gpc1_1 gpc184 (
      {stage0_4[29]},
      {stage1_4[27]}
   );
   gpc1_1 gpc185 (
      {stage0_4[30]},
      {stage1_4[28]}
   );
   gpc1_1 gpc186 (
      {stage0_4[31]},
      {stage1_4[29]}
   );
   gpc1_1 gpc187 (
      {stage0_5[27]},
      {stage1_5[9]}
   );
   gpc1_1 gpc188 (
      {stage0_5[28]},
      {stage1_5[10]}
   );
   gpc1_1 gpc189 (
      {stage0_5[29]},
      {stage1_5[11]}
   );
   gpc1_1 gpc190 (
      {stage0_5[30]},
      {stage1_5[12]}
   );
   gpc1_1 gpc191 (
      {stage0_5[31]},
      {stage1_5[13]}
   );
   gpc1_1 gpc192 (
      {stage0_6[10]},
      {stage1_6[7]}
   );
   gpc1_1 gpc193 (
      {stage0_6[11]},
      {stage1_6[8]}
   );
   gpc1_1 gpc194 (
      {stage0_6[12]},
      {stage1_6[9]}
   );
   gpc1_1 gpc195 (
      {stage0_6[13]},
      {stage1_6[10]}
   );
   gpc1_1 gpc196 (
      {stage0_6[14]},
      {stage1_6[11]}
   );
   gpc1_1 gpc197 (
      {stage0_6[15]},
      {stage1_6[12]}
   );
   gpc1_1 gpc198 (
      {stage0_6[16]},
      {stage1_6[13]}
   );
   gpc1_1 gpc199 (
      {stage0_6[17]},
      {stage1_6[14]}
   );
   gpc1_1 gpc200 (
      {stage0_6[18]},
      {stage1_6[15]}
   );
   gpc1_1 gpc201 (
      {stage0_6[19]},
      {stage1_6[16]}
   );
   gpc1_1 gpc202 (
      {stage0_6[20]},
      {stage1_6[17]}
   );
   gpc1_1 gpc203 (
      {stage0_6[21]},
      {stage1_6[18]}
   );
   gpc1_1 gpc204 (
      {stage0_6[22]},
      {stage1_6[19]}
   );
   gpc1_1 gpc205 (
      {stage0_6[23]},
      {stage1_6[20]}
   );
   gpc1_1 gpc206 (
      {stage0_6[24]},
      {stage1_6[21]}
   );
   gpc1_1 gpc207 (
      {stage0_6[25]},
      {stage1_6[22]}
   );
   gpc1_1 gpc208 (
      {stage0_6[26]},
      {stage1_6[23]}
   );
   gpc1_1 gpc209 (
      {stage0_6[27]},
      {stage1_6[24]}
   );
   gpc1_1 gpc210 (
      {stage0_6[28]},
      {stage1_6[25]}
   );
   gpc1_1 gpc211 (
      {stage0_6[29]},
      {stage1_6[26]}
   );
   gpc1_1 gpc212 (
      {stage0_6[30]},
      {stage1_6[27]}
   );
   gpc1_1 gpc213 (
      {stage0_6[31]},
      {stage1_6[28]}
   );
   gpc1_1 gpc214 (
      {stage0_7[31]},
      {stage1_7[8]}
   );
   gpc1_1 gpc215 (
      {stage0_8[24]},
      {stage1_8[11]}
   );
   gpc1_1 gpc216 (
      {stage0_8[25]},
      {stage1_8[12]}
   );
   gpc1_1 gpc217 (
      {stage0_8[26]},
      {stage1_8[13]}
   );
   gpc1_1 gpc218 (
      {stage0_8[27]},
      {stage1_8[14]}
   );
   gpc1_1 gpc219 (
      {stage0_8[28]},
      {stage1_8[15]}
   );
   gpc1_1 gpc220 (
      {stage0_8[29]},
      {stage1_8[16]}
   );
   gpc1_1 gpc221 (
      {stage0_8[30]},
      {stage1_8[17]}
   );
   gpc1_1 gpc222 (
      {stage0_8[31]},
      {stage1_8[18]}
   );
   gpc1_1 gpc223 (
      {stage0_9[29]},
      {stage1_9[13]}
   );
   gpc1_1 gpc224 (
      {stage0_9[30]},
      {stage1_9[14]}
   );
   gpc1_1 gpc225 (
      {stage0_9[31]},
      {stage1_9[15]}
   );
   gpc1_1 gpc226 (
      {stage0_10[23]},
      {stage1_10[9]}
   );
   gpc1_1 gpc227 (
      {stage0_10[24]},
      {stage1_10[10]}
   );
   gpc1_1 gpc228 (
      {stage0_10[25]},
      {stage1_10[11]}
   );
   gpc1_1 gpc229 (
      {stage0_10[26]},
      {stage1_10[12]}
   );
   gpc1_1 gpc230 (
      {stage0_10[27]},
      {stage1_10[13]}
   );
   gpc1_1 gpc231 (
      {stage0_10[28]},
      {stage1_10[14]}
   );
   gpc1_1 gpc232 (
      {stage0_10[29]},
      {stage1_10[15]}
   );
   gpc1_1 gpc233 (
      {stage0_10[30]},
      {stage1_10[16]}
   );
   gpc1_1 gpc234 (
      {stage0_10[31]},
      {stage1_10[17]}
   );
   gpc1_1 gpc235 (
      {stage0_11[25]},
      {stage1_11[10]}
   );
   gpc1_1 gpc236 (
      {stage0_11[26]},
      {stage1_11[11]}
   );
   gpc1_1 gpc237 (
      {stage0_11[27]},
      {stage1_11[12]}
   );
   gpc1_1 gpc238 (
      {stage0_11[28]},
      {stage1_11[13]}
   );
   gpc1_1 gpc239 (
      {stage0_11[29]},
      {stage1_11[14]}
   );
   gpc1_1 gpc240 (
      {stage0_11[30]},
      {stage1_11[15]}
   );
   gpc1_1 gpc241 (
      {stage0_11[31]},
      {stage1_11[16]}
   );
   gpc1_1 gpc242 (
      {stage0_12[25]},
      {stage1_12[12]}
   );
   gpc1_1 gpc243 (
      {stage0_12[26]},
      {stage1_12[13]}
   );
   gpc1_1 gpc244 (
      {stage0_12[27]},
      {stage1_12[14]}
   );
   gpc1_1 gpc245 (
      {stage0_12[28]},
      {stage1_12[15]}
   );
   gpc1_1 gpc246 (
      {stage0_12[29]},
      {stage1_12[16]}
   );
   gpc1_1 gpc247 (
      {stage0_12[30]},
      {stage1_12[17]}
   );
   gpc1_1 gpc248 (
      {stage0_12[31]},
      {stage1_12[18]}
   );
   gpc1_1 gpc249 (
      {stage0_13[30]},
      {stage1_13[12]}
   );
   gpc1_1 gpc250 (
      {stage0_13[31]},
      {stage1_13[13]}
   );
   gpc1_1 gpc251 (
      {stage0_14[24]},
      {stage1_14[9]}
   );
   gpc1_1 gpc252 (
      {stage0_14[25]},
      {stage1_14[10]}
   );
   gpc1_1 gpc253 (
      {stage0_14[26]},
      {stage1_14[11]}
   );
   gpc1_1 gpc254 (
      {stage0_14[27]},
      {stage1_14[12]}
   );
   gpc1_1 gpc255 (
      {stage0_14[28]},
      {stage1_14[13]}
   );
   gpc1_1 gpc256 (
      {stage0_14[29]},
      {stage1_14[14]}
   );
   gpc1_1 gpc257 (
      {stage0_14[30]},
      {stage1_14[15]}
   );
   gpc1_1 gpc258 (
      {stage0_14[31]},
      {stage1_14[16]}
   );
   gpc1_1 gpc259 (
      {stage0_15[29]},
      {stage1_15[10]}
   );
   gpc1_1 gpc260 (
      {stage0_15[30]},
      {stage1_15[11]}
   );
   gpc1_1 gpc261 (
      {stage0_15[31]},
      {stage1_15[12]}
   );
   gpc1_1 gpc262 (
      {stage0_16[12]},
      {stage1_16[11]}
   );
   gpc1_1 gpc263 (
      {stage0_16[13]},
      {stage1_16[12]}
   );
   gpc1_1 gpc264 (
      {stage0_16[14]},
      {stage1_16[13]}
   );
   gpc1_1 gpc265 (
      {stage0_16[15]},
      {stage1_16[14]}
   );
   gpc1_1 gpc266 (
      {stage0_16[16]},
      {stage1_16[15]}
   );
   gpc1_1 gpc267 (
      {stage0_16[17]},
      {stage1_16[16]}
   );
   gpc1_1 gpc268 (
      {stage0_16[18]},
      {stage1_16[17]}
   );
   gpc1_1 gpc269 (
      {stage0_16[19]},
      {stage1_16[18]}
   );
   gpc1_1 gpc270 (
      {stage0_16[20]},
      {stage1_16[19]}
   );
   gpc1_1 gpc271 (
      {stage0_16[21]},
      {stage1_16[20]}
   );
   gpc1_1 gpc272 (
      {stage0_16[22]},
      {stage1_16[21]}
   );
   gpc1_1 gpc273 (
      {stage0_16[23]},
      {stage1_16[22]}
   );
   gpc1_1 gpc274 (
      {stage0_16[24]},
      {stage1_16[23]}
   );
   gpc1_1 gpc275 (
      {stage0_16[25]},
      {stage1_16[24]}
   );
   gpc1_1 gpc276 (
      {stage0_16[26]},
      {stage1_16[25]}
   );
   gpc1_1 gpc277 (
      {stage0_16[27]},
      {stage1_16[26]}
   );
   gpc1_1 gpc278 (
      {stage0_16[28]},
      {stage1_16[27]}
   );
   gpc1_1 gpc279 (
      {stage0_16[29]},
      {stage1_16[28]}
   );
   gpc1_1 gpc280 (
      {stage0_16[30]},
      {stage1_16[29]}
   );
   gpc1_1 gpc281 (
      {stage0_16[31]},
      {stage1_16[30]}
   );
   gpc1_1 gpc282 (
      {stage0_17[19]},
      {stage1_17[9]}
   );
   gpc1_1 gpc283 (
      {stage0_17[20]},
      {stage1_17[10]}
   );
   gpc1_1 gpc284 (
      {stage0_17[21]},
      {stage1_17[11]}
   );
   gpc1_1 gpc285 (
      {stage0_17[22]},
      {stage1_17[12]}
   );
   gpc1_1 gpc286 (
      {stage0_17[23]},
      {stage1_17[13]}
   );
   gpc1_1 gpc287 (
      {stage0_17[24]},
      {stage1_17[14]}
   );
   gpc1_1 gpc288 (
      {stage0_17[25]},
      {stage1_17[15]}
   );
   gpc1_1 gpc289 (
      {stage0_17[26]},
      {stage1_17[16]}
   );
   gpc1_1 gpc290 (
      {stage0_17[27]},
      {stage1_17[17]}
   );
   gpc1_1 gpc291 (
      {stage0_17[28]},
      {stage1_17[18]}
   );
   gpc1_1 gpc292 (
      {stage0_17[29]},
      {stage1_17[19]}
   );
   gpc1_1 gpc293 (
      {stage0_17[30]},
      {stage1_17[20]}
   );
   gpc1_1 gpc294 (
      {stage0_17[31]},
      {stage1_17[21]}
   );
   gpc1_1 gpc295 (
      {stage0_18[29]},
      {stage1_18[8]}
   );
   gpc1_1 gpc296 (
      {stage0_18[30]},
      {stage1_18[9]}
   );
   gpc1_1 gpc297 (
      {stage0_18[31]},
      {stage1_18[10]}
   );
   gpc1_1 gpc298 (
      {stage0_19[23]},
      {stage1_19[10]}
   );
   gpc1_1 gpc299 (
      {stage0_19[24]},
      {stage1_19[11]}
   );
   gpc1_1 gpc300 (
      {stage0_19[25]},
      {stage1_19[12]}
   );
   gpc1_1 gpc301 (
      {stage0_19[26]},
      {stage1_19[13]}
   );
   gpc1_1 gpc302 (
      {stage0_19[27]},
      {stage1_19[14]}
   );
   gpc1_1 gpc303 (
      {stage0_19[28]},
      {stage1_19[15]}
   );
   gpc1_1 gpc304 (
      {stage0_19[29]},
      {stage1_19[16]}
   );
   gpc1_1 gpc305 (
      {stage0_19[30]},
      {stage1_19[17]}
   );
   gpc1_1 gpc306 (
      {stage0_19[31]},
      {stage1_19[18]}
   );
   gpc1_1 gpc307 (
      {stage0_21[26]},
      {stage1_21[12]}
   );
   gpc1_1 gpc308 (
      {stage0_21[27]},
      {stage1_21[13]}
   );
   gpc1_1 gpc309 (
      {stage0_21[28]},
      {stage1_21[14]}
   );
   gpc1_1 gpc310 (
      {stage0_21[29]},
      {stage1_21[15]}
   );
   gpc1_1 gpc311 (
      {stage0_21[30]},
      {stage1_21[16]}
   );
   gpc1_1 gpc312 (
      {stage0_21[31]},
      {stage1_21[17]}
   );
   gpc1_1 gpc313 (
      {stage0_22[31]},
      {stage1_22[13]}
   );
   gpc1_1 gpc314 (
      {stage0_23[25]},
      {stage1_23[11]}
   );
   gpc1_1 gpc315 (
      {stage0_23[26]},
      {stage1_23[12]}
   );
   gpc1_1 gpc316 (
      {stage0_23[27]},
      {stage1_23[13]}
   );
   gpc1_1 gpc317 (
      {stage0_23[28]},
      {stage1_23[14]}
   );
   gpc1_1 gpc318 (
      {stage0_23[29]},
      {stage1_23[15]}
   );
   gpc1_1 gpc319 (
      {stage0_23[30]},
      {stage1_23[16]}
   );
   gpc1_1 gpc320 (
      {stage0_23[31]},
      {stage1_23[17]}
   );
   gpc1_1 gpc321 (
      {stage0_25[27]},
      {stage1_25[13]}
   );
   gpc1_1 gpc322 (
      {stage0_25[28]},
      {stage1_25[14]}
   );
   gpc1_1 gpc323 (
      {stage0_25[29]},
      {stage1_25[15]}
   );
   gpc1_1 gpc324 (
      {stage0_25[30]},
      {stage1_25[16]}
   );
   gpc1_1 gpc325 (
      {stage0_25[31]},
      {stage1_25[17]}
   );
   gpc1_1 gpc326 (
      {stage0_26[27]},
      {stage1_26[12]}
   );
   gpc1_1 gpc327 (
      {stage0_26[28]},
      {stage1_26[13]}
   );
   gpc1_1 gpc328 (
      {stage0_26[29]},
      {stage1_26[14]}
   );
   gpc1_1 gpc329 (
      {stage0_26[30]},
      {stage1_26[15]}
   );
   gpc1_1 gpc330 (
      {stage0_26[31]},
      {stage1_26[16]}
   );
   gpc1_1 gpc331 (
      {stage0_27[31]},
      {stage1_27[10]}
   );
   gpc1_1 gpc332 (
      {stage0_28[29]},
      {stage1_28[13]}
   );
   gpc1_1 gpc333 (
      {stage0_28[30]},
      {stage1_28[14]}
   );
   gpc1_1 gpc334 (
      {stage0_28[31]},
      {stage1_28[15]}
   );
   gpc1_1 gpc335 (
      {stage0_29[28]},
      {stage1_29[14]}
   );
   gpc1_1 gpc336 (
      {stage0_29[29]},
      {stage1_29[15]}
   );
   gpc1_1 gpc337 (
      {stage0_29[30]},
      {stage1_29[16]}
   );
   gpc1_1 gpc338 (
      {stage0_29[31]},
      {stage1_29[17]}
   );
   gpc1_1 gpc339 (
      {stage0_31[25]},
      {stage1_31[10]}
   );
   gpc1_1 gpc340 (
      {stage0_31[26]},
      {stage1_31[11]}
   );
   gpc1_1 gpc341 (
      {stage0_31[27]},
      {stage1_31[12]}
   );
   gpc1_1 gpc342 (
      {stage0_31[28]},
      {stage1_31[13]}
   );
   gpc1_1 gpc343 (
      {stage0_31[29]},
      {stage1_31[14]}
   );
   gpc1_1 gpc344 (
      {stage0_31[30]},
      {stage1_31[15]}
   );
   gpc1_1 gpc345 (
      {stage0_31[31]},
      {stage1_31[16]}
   );
   gpc1_1 gpc346 (
      {stage0_32[18]},
      {stage1_32[11]}
   );
   gpc1_1 gpc347 (
      {stage0_32[19]},
      {stage1_32[12]}
   );
   gpc1_1 gpc348 (
      {stage0_32[20]},
      {stage1_32[13]}
   );
   gpc1_1 gpc349 (
      {stage0_32[21]},
      {stage1_32[14]}
   );
   gpc1_1 gpc350 (
      {stage0_32[22]},
      {stage1_32[15]}
   );
   gpc1_1 gpc351 (
      {stage0_32[23]},
      {stage1_32[16]}
   );
   gpc1_1 gpc352 (
      {stage0_32[24]},
      {stage1_32[17]}
   );
   gpc1_1 gpc353 (
      {stage0_32[25]},
      {stage1_32[18]}
   );
   gpc1_1 gpc354 (
      {stage0_32[26]},
      {stage1_32[19]}
   );
   gpc1_1 gpc355 (
      {stage0_32[27]},
      {stage1_32[20]}
   );
   gpc1_1 gpc356 (
      {stage0_32[28]},
      {stage1_32[21]}
   );
   gpc1_1 gpc357 (
      {stage0_32[29]},
      {stage1_32[22]}
   );
   gpc1_1 gpc358 (
      {stage0_32[30]},
      {stage1_32[23]}
   );
   gpc1_1 gpc359 (
      {stage0_32[31]},
      {stage1_32[24]}
   );
   gpc1_1 gpc360 (
      {stage0_33[24]},
      {stage1_33[11]}
   );
   gpc1_1 gpc361 (
      {stage0_33[25]},
      {stage1_33[12]}
   );
   gpc1_1 gpc362 (
      {stage0_33[26]},
      {stage1_33[13]}
   );
   gpc1_1 gpc363 (
      {stage0_33[27]},
      {stage1_33[14]}
   );
   gpc1_1 gpc364 (
      {stage0_33[28]},
      {stage1_33[15]}
   );
   gpc1_1 gpc365 (
      {stage0_33[29]},
      {stage1_33[16]}
   );
   gpc1_1 gpc366 (
      {stage0_33[30]},
      {stage1_33[17]}
   );
   gpc1_1 gpc367 (
      {stage0_33[31]},
      {stage1_33[18]}
   );
   gpc1_1 gpc368 (
      {stage0_34[20]},
      {stage1_34[9]}
   );
   gpc1_1 gpc369 (
      {stage0_34[21]},
      {stage1_34[10]}
   );
   gpc1_1 gpc370 (
      {stage0_34[22]},
      {stage1_34[11]}
   );
   gpc1_1 gpc371 (
      {stage0_34[23]},
      {stage1_34[12]}
   );
   gpc1_1 gpc372 (
      {stage0_34[24]},
      {stage1_34[13]}
   );
   gpc1_1 gpc373 (
      {stage0_34[25]},
      {stage1_34[14]}
   );
   gpc1_1 gpc374 (
      {stage0_34[26]},
      {stage1_34[15]}
   );
   gpc1_1 gpc375 (
      {stage0_34[27]},
      {stage1_34[16]}
   );
   gpc1_1 gpc376 (
      {stage0_34[28]},
      {stage1_34[17]}
   );
   gpc1_1 gpc377 (
      {stage0_34[29]},
      {stage1_34[18]}
   );
   gpc1_1 gpc378 (
      {stage0_34[30]},
      {stage1_34[19]}
   );
   gpc1_1 gpc379 (
      {stage0_34[31]},
      {stage1_34[20]}
   );
   gpc1_1 gpc380 (
      {stage0_35[27]},
      {stage1_35[8]}
   );
   gpc1_1 gpc381 (
      {stage0_35[28]},
      {stage1_35[9]}
   );
   gpc1_1 gpc382 (
      {stage0_35[29]},
      {stage1_35[10]}
   );
   gpc1_1 gpc383 (
      {stage0_35[30]},
      {stage1_35[11]}
   );
   gpc1_1 gpc384 (
      {stage0_35[31]},
      {stage1_35[12]}
   );
   gpc1_1 gpc385 (
      {stage0_36[30]},
      {stage1_36[11]}
   );
   gpc1_1 gpc386 (
      {stage0_36[31]},
      {stage1_36[12]}
   );
   gpc1_1 gpc387 (
      {stage0_38[25]},
      {stage1_38[11]}
   );
   gpc1_1 gpc388 (
      {stage0_38[26]},
      {stage1_38[12]}
   );
   gpc1_1 gpc389 (
      {stage0_38[27]},
      {stage1_38[13]}
   );
   gpc1_1 gpc390 (
      {stage0_38[28]},
      {stage1_38[14]}
   );
   gpc1_1 gpc391 (
      {stage0_38[29]},
      {stage1_38[15]}
   );
   gpc1_1 gpc392 (
      {stage0_38[30]},
      {stage1_38[16]}
   );
   gpc1_1 gpc393 (
      {stage0_38[31]},
      {stage1_38[17]}
   );
   gpc1_1 gpc394 (
      {stage0_39[27]},
      {stage1_39[10]}
   );
   gpc1_1 gpc395 (
      {stage0_39[28]},
      {stage1_39[11]}
   );
   gpc1_1 gpc396 (
      {stage0_39[29]},
      {stage1_39[12]}
   );
   gpc1_1 gpc397 (
      {stage0_39[30]},
      {stage1_39[13]}
   );
   gpc1_1 gpc398 (
      {stage0_39[31]},
      {stage1_39[14]}
   );
   gpc1_1 gpc399 (
      {stage0_40[30]},
      {stage1_40[14]}
   );
   gpc1_1 gpc400 (
      {stage0_40[31]},
      {stage1_40[15]}
   );
   gpc1_1 gpc401 (
      {stage0_41[24]},
      {stage1_41[12]}
   );
   gpc1_1 gpc402 (
      {stage0_41[25]},
      {stage1_41[13]}
   );
   gpc1_1 gpc403 (
      {stage0_41[26]},
      {stage1_41[14]}
   );
   gpc1_1 gpc404 (
      {stage0_41[27]},
      {stage1_41[15]}
   );
   gpc1_1 gpc405 (
      {stage0_41[28]},
      {stage1_41[16]}
   );
   gpc1_1 gpc406 (
      {stage0_41[29]},
      {stage1_41[17]}
   );
   gpc1_1 gpc407 (
      {stage0_41[30]},
      {stage1_41[18]}
   );
   gpc1_1 gpc408 (
      {stage0_41[31]},
      {stage1_41[19]}
   );
   gpc1_1 gpc409 (
      {stage0_42[29]},
      {stage1_42[10]}
   );
   gpc1_1 gpc410 (
      {stage0_42[30]},
      {stage1_42[11]}
   );
   gpc1_1 gpc411 (
      {stage0_42[31]},
      {stage1_42[12]}
   );
   gpc1_1 gpc412 (
      {stage0_43[29]},
      {stage1_43[11]}
   );
   gpc1_1 gpc413 (
      {stage0_43[30]},
      {stage1_43[12]}
   );
   gpc1_1 gpc414 (
      {stage0_43[31]},
      {stage1_43[13]}
   );
   gpc1_1 gpc415 (
      {stage0_45[18]},
      {stage1_45[11]}
   );
   gpc1_1 gpc416 (
      {stage0_45[19]},
      {stage1_45[12]}
   );
   gpc1_1 gpc417 (
      {stage0_45[20]},
      {stage1_45[13]}
   );
   gpc1_1 gpc418 (
      {stage0_45[21]},
      {stage1_45[14]}
   );
   gpc1_1 gpc419 (
      {stage0_45[22]},
      {stage1_45[15]}
   );
   gpc1_1 gpc420 (
      {stage0_45[23]},
      {stage1_45[16]}
   );
   gpc1_1 gpc421 (
      {stage0_45[24]},
      {stage1_45[17]}
   );
   gpc1_1 gpc422 (
      {stage0_45[25]},
      {stage1_45[18]}
   );
   gpc1_1 gpc423 (
      {stage0_45[26]},
      {stage1_45[19]}
   );
   gpc1_1 gpc424 (
      {stage0_45[27]},
      {stage1_45[20]}
   );
   gpc1_1 gpc425 (
      {stage0_45[28]},
      {stage1_45[21]}
   );
   gpc1_1 gpc426 (
      {stage0_45[29]},
      {stage1_45[22]}
   );
   gpc1_1 gpc427 (
      {stage0_45[30]},
      {stage1_45[23]}
   );
   gpc1_1 gpc428 (
      {stage0_45[31]},
      {stage1_45[24]}
   );
   gpc1_1 gpc429 (
      {stage0_46[29]},
      {stage1_46[9]}
   );
   gpc1_1 gpc430 (
      {stage0_46[30]},
      {stage1_46[10]}
   );
   gpc1_1 gpc431 (
      {stage0_46[31]},
      {stage1_46[11]}
   );
   gpc1_1 gpc432 (
      {stage0_47[25]},
      {stage1_47[11]}
   );
   gpc1_1 gpc433 (
      {stage0_47[26]},
      {stage1_47[12]}
   );
   gpc1_1 gpc434 (
      {stage0_47[27]},
      {stage1_47[13]}
   );
   gpc1_1 gpc435 (
      {stage0_47[28]},
      {stage1_47[14]}
   );
   gpc1_1 gpc436 (
      {stage0_47[29]},
      {stage1_47[15]}
   );
   gpc1_1 gpc437 (
      {stage0_47[30]},
      {stage1_47[16]}
   );
   gpc1_1 gpc438 (
      {stage0_47[31]},
      {stage1_47[17]}
   );
   gpc1_1 gpc439 (
      {stage0_48[24]},
      {stage1_48[12]}
   );
   gpc1_1 gpc440 (
      {stage0_48[25]},
      {stage1_48[13]}
   );
   gpc1_1 gpc441 (
      {stage0_48[26]},
      {stage1_48[14]}
   );
   gpc1_1 gpc442 (
      {stage0_48[27]},
      {stage1_48[15]}
   );
   gpc1_1 gpc443 (
      {stage0_48[28]},
      {stage1_48[16]}
   );
   gpc1_1 gpc444 (
      {stage0_48[29]},
      {stage1_48[17]}
   );
   gpc1_1 gpc445 (
      {stage0_48[30]},
      {stage1_48[18]}
   );
   gpc1_1 gpc446 (
      {stage0_48[31]},
      {stage1_48[19]}
   );
   gpc1_1 gpc447 (
      {stage0_49[21]},
      {stage1_49[9]}
   );
   gpc1_1 gpc448 (
      {stage0_49[22]},
      {stage1_49[10]}
   );
   gpc1_1 gpc449 (
      {stage0_49[23]},
      {stage1_49[11]}
   );
   gpc1_1 gpc450 (
      {stage0_49[24]},
      {stage1_49[12]}
   );
   gpc1_1 gpc451 (
      {stage0_49[25]},
      {stage1_49[13]}
   );
   gpc1_1 gpc452 (
      {stage0_49[26]},
      {stage1_49[14]}
   );
   gpc1_1 gpc453 (
      {stage0_49[27]},
      {stage1_49[15]}
   );
   gpc1_1 gpc454 (
      {stage0_49[28]},
      {stage1_49[16]}
   );
   gpc1_1 gpc455 (
      {stage0_49[29]},
      {stage1_49[17]}
   );
   gpc1_1 gpc456 (
      {stage0_49[30]},
      {stage1_49[18]}
   );
   gpc1_1 gpc457 (
      {stage0_49[31]},
      {stage1_49[19]}
   );
   gpc1_1 gpc458 (
      {stage0_50[30]},
      {stage1_50[10]}
   );
   gpc1_1 gpc459 (
      {stage0_50[31]},
      {stage1_50[11]}
   );
   gpc1_1 gpc460 (
      {stage0_51[23]},
      {stage1_51[12]}
   );
   gpc1_1 gpc461 (
      {stage0_51[24]},
      {stage1_51[13]}
   );
   gpc1_1 gpc462 (
      {stage0_51[25]},
      {stage1_51[14]}
   );
   gpc1_1 gpc463 (
      {stage0_51[26]},
      {stage1_51[15]}
   );
   gpc1_1 gpc464 (
      {stage0_51[27]},
      {stage1_51[16]}
   );
   gpc1_1 gpc465 (
      {stage0_51[28]},
      {stage1_51[17]}
   );
   gpc1_1 gpc466 (
      {stage0_51[29]},
      {stage1_51[18]}
   );
   gpc1_1 gpc467 (
      {stage0_51[30]},
      {stage1_51[19]}
   );
   gpc1_1 gpc468 (
      {stage0_51[31]},
      {stage1_51[20]}
   );
   gpc1_1 gpc469 (
      {stage0_53[18]},
      {stage1_53[9]}
   );
   gpc1_1 gpc470 (
      {stage0_53[19]},
      {stage1_53[10]}
   );
   gpc1_1 gpc471 (
      {stage0_53[20]},
      {stage1_53[11]}
   );
   gpc1_1 gpc472 (
      {stage0_53[21]},
      {stage1_53[12]}
   );
   gpc1_1 gpc473 (
      {stage0_53[22]},
      {stage1_53[13]}
   );
   gpc1_1 gpc474 (
      {stage0_53[23]},
      {stage1_53[14]}
   );
   gpc1_1 gpc475 (
      {stage0_53[24]},
      {stage1_53[15]}
   );
   gpc1_1 gpc476 (
      {stage0_53[25]},
      {stage1_53[16]}
   );
   gpc1_1 gpc477 (
      {stage0_53[26]},
      {stage1_53[17]}
   );
   gpc1_1 gpc478 (
      {stage0_53[27]},
      {stage1_53[18]}
   );
   gpc1_1 gpc479 (
      {stage0_53[28]},
      {stage1_53[19]}
   );
   gpc1_1 gpc480 (
      {stage0_53[29]},
      {stage1_53[20]}
   );
   gpc1_1 gpc481 (
      {stage0_53[30]},
      {stage1_53[21]}
   );
   gpc1_1 gpc482 (
      {stage0_53[31]},
      {stage1_53[22]}
   );
   gpc1_1 gpc483 (
      {stage0_55[13]},
      {stage1_55[11]}
   );
   gpc1_1 gpc484 (
      {stage0_55[14]},
      {stage1_55[12]}
   );
   gpc1_1 gpc485 (
      {stage0_55[15]},
      {stage1_55[13]}
   );
   gpc1_1 gpc486 (
      {stage0_55[16]},
      {stage1_55[14]}
   );
   gpc1_1 gpc487 (
      {stage0_55[17]},
      {stage1_55[15]}
   );
   gpc1_1 gpc488 (
      {stage0_55[18]},
      {stage1_55[16]}
   );
   gpc1_1 gpc489 (
      {stage0_55[19]},
      {stage1_55[17]}
   );
   gpc1_1 gpc490 (
      {stage0_55[20]},
      {stage1_55[18]}
   );
   gpc1_1 gpc491 (
      {stage0_55[21]},
      {stage1_55[19]}
   );
   gpc1_1 gpc492 (
      {stage0_55[22]},
      {stage1_55[20]}
   );
   gpc1_1 gpc493 (
      {stage0_55[23]},
      {stage1_55[21]}
   );
   gpc1_1 gpc494 (
      {stage0_55[24]},
      {stage1_55[22]}
   );
   gpc1_1 gpc495 (
      {stage0_55[25]},
      {stage1_55[23]}
   );
   gpc1_1 gpc496 (
      {stage0_55[26]},
      {stage1_55[24]}
   );
   gpc1_1 gpc497 (
      {stage0_55[27]},
      {stage1_55[25]}
   );
   gpc1_1 gpc498 (
      {stage0_55[28]},
      {stage1_55[26]}
   );
   gpc1_1 gpc499 (
      {stage0_55[29]},
      {stage1_55[27]}
   );
   gpc1_1 gpc500 (
      {stage0_55[30]},
      {stage1_55[28]}
   );
   gpc1_1 gpc501 (
      {stage0_55[31]},
      {stage1_55[29]}
   );
   gpc1_1 gpc502 (
      {stage0_56[28]},
      {stage1_56[11]}
   );
   gpc1_1 gpc503 (
      {stage0_56[29]},
      {stage1_56[12]}
   );
   gpc1_1 gpc504 (
      {stage0_56[30]},
      {stage1_56[13]}
   );
   gpc1_1 gpc505 (
      {stage0_56[31]},
      {stage1_56[14]}
   );
   gpc1_1 gpc506 (
      {stage0_57[25]},
      {stage1_57[10]}
   );
   gpc1_1 gpc507 (
      {stage0_57[26]},
      {stage1_57[11]}
   );
   gpc1_1 gpc508 (
      {stage0_57[27]},
      {stage1_57[12]}
   );
   gpc1_1 gpc509 (
      {stage0_57[28]},
      {stage1_57[13]}
   );
   gpc1_1 gpc510 (
      {stage0_57[29]},
      {stage1_57[14]}
   );
   gpc1_1 gpc511 (
      {stage0_57[30]},
      {stage1_57[15]}
   );
   gpc1_1 gpc512 (
      {stage0_57[31]},
      {stage1_57[16]}
   );
   gpc1_1 gpc513 (
      {stage0_58[27]},
      {stage1_58[9]}
   );
   gpc1_1 gpc514 (
      {stage0_58[28]},
      {stage1_58[10]}
   );
   gpc1_1 gpc515 (
      {stage0_58[29]},
      {stage1_58[11]}
   );
   gpc1_1 gpc516 (
      {stage0_58[30]},
      {stage1_58[12]}
   );
   gpc1_1 gpc517 (
      {stage0_58[31]},
      {stage1_58[13]}
   );
   gpc1_1 gpc518 (
      {stage0_59[18]},
      {stage1_59[10]}
   );
   gpc1_1 gpc519 (
      {stage0_59[19]},
      {stage1_59[11]}
   );
   gpc1_1 gpc520 (
      {stage0_59[20]},
      {stage1_59[12]}
   );
   gpc1_1 gpc521 (
      {stage0_59[21]},
      {stage1_59[13]}
   );
   gpc1_1 gpc522 (
      {stage0_59[22]},
      {stage1_59[14]}
   );
   gpc1_1 gpc523 (
      {stage0_59[23]},
      {stage1_59[15]}
   );
   gpc1_1 gpc524 (
      {stage0_59[24]},
      {stage1_59[16]}
   );
   gpc1_1 gpc525 (
      {stage0_59[25]},
      {stage1_59[17]}
   );
   gpc1_1 gpc526 (
      {stage0_59[26]},
      {stage1_59[18]}
   );
   gpc1_1 gpc527 (
      {stage0_59[27]},
      {stage1_59[19]}
   );
   gpc1_1 gpc528 (
      {stage0_59[28]},
      {stage1_59[20]}
   );
   gpc1_1 gpc529 (
      {stage0_59[29]},
      {stage1_59[21]}
   );
   gpc1_1 gpc530 (
      {stage0_59[30]},
      {stage1_59[22]}
   );
   gpc1_1 gpc531 (
      {stage0_59[31]},
      {stage1_59[23]}
   );
   gpc1_1 gpc532 (
      {stage0_60[30]},
      {stage1_60[11]}
   );
   gpc1_1 gpc533 (
      {stage0_60[31]},
      {stage1_60[12]}
   );
   gpc1_1 gpc534 (
      {stage0_62[26]},
      {stage1_62[11]}
   );
   gpc1_1 gpc535 (
      {stage0_62[27]},
      {stage1_62[12]}
   );
   gpc1_1 gpc536 (
      {stage0_62[28]},
      {stage1_62[13]}
   );
   gpc1_1 gpc537 (
      {stage0_62[29]},
      {stage1_62[14]}
   );
   gpc1_1 gpc538 (
      {stage0_62[30]},
      {stage1_62[15]}
   );
   gpc1_1 gpc539 (
      {stage0_62[31]},
      {stage1_62[16]}
   );
   gpc1_1 gpc540 (
      {stage0_63[31]},
      {stage1_63[10]}
   );
   gpc606_5 gpc541 (
      {stage1_1[0], stage1_1[1], stage1_1[2], stage1_1[3], stage1_1[4], stage1_1[5]},
      {stage1_3[0], stage1_3[1], stage1_3[2], stage1_3[3], stage1_3[4], stage1_3[5]},
      {stage2_5[0],stage2_4[0],stage2_3[0],stage2_2[0],stage2_1[0]}
   );
   gpc606_5 gpc542 (
      {stage1_2[0], stage1_2[1], stage1_2[2], stage1_2[3], stage1_2[4], stage1_2[5]},
      {stage1_4[0], stage1_4[1], stage1_4[2], stage1_4[3], stage1_4[4], stage1_4[5]},
      {stage2_6[0],stage2_5[1],stage2_4[1],stage2_3[1],stage2_2[1]}
   );
   gpc615_5 gpc543 (
      {stage1_2[6], stage1_2[7], stage1_2[8], stage1_2[9], stage1_2[10]},
      {stage1_3[6]},
      {stage1_4[6], stage1_4[7], stage1_4[8], stage1_4[9], stage1_4[10], stage1_4[11]},
      {stage2_6[1],stage2_5[2],stage2_4[2],stage2_3[2],stage2_2[2]}
   );
   gpc615_5 gpc544 (
      {stage1_2[11], stage1_2[12], stage1_2[13], stage1_2[14], stage1_2[15]},
      {stage1_3[7]},
      {stage1_4[12], stage1_4[13], stage1_4[14], stage1_4[15], stage1_4[16], stage1_4[17]},
      {stage2_6[2],stage2_5[3],stage2_4[3],stage2_3[3],stage2_2[3]}
   );
   gpc615_5 gpc545 (
      {stage1_2[16], stage1_2[17], stage1_2[18], stage1_2[19], stage1_2[20]},
      {stage1_3[8]},
      {stage1_4[18], stage1_4[19], stage1_4[20], stage1_4[21], stage1_4[22], stage1_4[23]},
      {stage2_6[3],stage2_5[4],stage2_4[4],stage2_3[4],stage2_2[4]}
   );
   gpc615_5 gpc546 (
      {stage1_3[9], stage1_3[10], stage1_3[11], stage1_3[12], stage1_3[13]},
      {stage1_4[24]},
      {stage1_5[0], stage1_5[1], stage1_5[2], stage1_5[3], stage1_5[4], stage1_5[5]},
      {stage2_7[0],stage2_6[4],stage2_5[5],stage2_4[5],stage2_3[5]}
   );
   gpc606_5 gpc547 (
      {stage1_4[25], stage1_4[26], stage1_4[27], stage1_4[28], stage1_4[29], 1'b0},
      {stage1_6[0], stage1_6[1], stage1_6[2], stage1_6[3], stage1_6[4], stage1_6[5]},
      {stage2_8[0],stage2_7[1],stage2_6[5],stage2_5[6],stage2_4[6]}
   );
   gpc606_5 gpc548 (
      {stage1_5[6], stage1_5[7], stage1_5[8], stage1_5[9], stage1_5[10], stage1_5[11]},
      {stage1_7[0], stage1_7[1], stage1_7[2], stage1_7[3], stage1_7[4], stage1_7[5]},
      {stage2_9[0],stage2_8[1],stage2_7[2],stage2_6[6],stage2_5[7]}
   );
   gpc615_5 gpc549 (
      {stage1_6[6], stage1_6[7], stage1_6[8], stage1_6[9], stage1_6[10]},
      {stage1_7[6]},
      {stage1_8[0], stage1_8[1], stage1_8[2], stage1_8[3], stage1_8[4], stage1_8[5]},
      {stage2_10[0],stage2_9[1],stage2_8[2],stage2_7[3],stage2_6[7]}
   );
   gpc615_5 gpc550 (
      {stage1_6[11], stage1_6[12], stage1_6[13], stage1_6[14], stage1_6[15]},
      {stage1_7[7]},
      {stage1_8[6], stage1_8[7], stage1_8[8], stage1_8[9], stage1_8[10], stage1_8[11]},
      {stage2_10[1],stage2_9[2],stage2_8[3],stage2_7[4],stage2_6[8]}
   );
   gpc615_5 gpc551 (
      {stage1_6[16], stage1_6[17], stage1_6[18], stage1_6[19], stage1_6[20]},
      {stage1_7[8]},
      {stage1_8[12], stage1_8[13], stage1_8[14], stage1_8[15], stage1_8[16], stage1_8[17]},
      {stage2_10[2],stage2_9[3],stage2_8[4],stage2_7[5],stage2_6[9]}
   );
   gpc606_5 gpc552 (
      {stage1_9[0], stage1_9[1], stage1_9[2], stage1_9[3], stage1_9[4], stage1_9[5]},
      {stage1_11[0], stage1_11[1], stage1_11[2], stage1_11[3], stage1_11[4], stage1_11[5]},
      {stage2_13[0],stage2_12[0],stage2_11[0],stage2_10[3],stage2_9[4]}
   );
   gpc606_5 gpc553 (
      {stage1_9[6], stage1_9[7], stage1_9[8], stage1_9[9], stage1_9[10], stage1_9[11]},
      {stage1_11[6], stage1_11[7], stage1_11[8], stage1_11[9], stage1_11[10], stage1_11[11]},
      {stage2_13[1],stage2_12[1],stage2_11[1],stage2_10[4],stage2_9[5]}
   );
   gpc606_5 gpc554 (
      {stage1_10[0], stage1_10[1], stage1_10[2], stage1_10[3], stage1_10[4], stage1_10[5]},
      {stage1_12[0], stage1_12[1], stage1_12[2], stage1_12[3], stage1_12[4], stage1_12[5]},
      {stage2_14[0],stage2_13[2],stage2_12[2],stage2_11[2],stage2_10[5]}
   );
   gpc606_5 gpc555 (
      {stage1_10[6], stage1_10[7], stage1_10[8], stage1_10[9], stage1_10[10], stage1_10[11]},
      {stage1_12[6], stage1_12[7], stage1_12[8], stage1_12[9], stage1_12[10], stage1_12[11]},
      {stage2_14[1],stage2_13[3],stage2_12[3],stage2_11[3],stage2_10[6]}
   );
   gpc606_5 gpc556 (
      {stage1_10[12], stage1_10[13], stage1_10[14], stage1_10[15], stage1_10[16], stage1_10[17]},
      {stage1_12[12], stage1_12[13], stage1_12[14], stage1_12[15], stage1_12[16], stage1_12[17]},
      {stage2_14[2],stage2_13[4],stage2_12[4],stage2_11[4],stage2_10[7]}
   );
   gpc615_5 gpc557 (
      {stage1_11[12], stage1_11[13], stage1_11[14], stage1_11[15], stage1_11[16]},
      {stage1_12[18]},
      {stage1_13[0], stage1_13[1], stage1_13[2], stage1_13[3], stage1_13[4], stage1_13[5]},
      {stage2_15[0],stage2_14[3],stage2_13[5],stage2_12[5],stage2_11[5]}
   );
   gpc606_5 gpc558 (
      {stage1_13[6], stage1_13[7], stage1_13[8], stage1_13[9], stage1_13[10], stage1_13[11]},
      {stage1_15[0], stage1_15[1], stage1_15[2], stage1_15[3], stage1_15[4], stage1_15[5]},
      {stage2_17[0],stage2_16[0],stage2_15[1],stage2_14[4],stage2_13[6]}
   );
   gpc1163_5 gpc559 (
      {stage1_14[0], stage1_14[1], stage1_14[2]},
      {stage1_15[6], stage1_15[7], stage1_15[8], stage1_15[9], stage1_15[10], stage1_15[11]},
      {stage1_16[0]},
      {stage1_17[0]},
      {stage2_18[0],stage2_17[1],stage2_16[1],stage2_15[2],stage2_14[5]}
   );
   gpc615_5 gpc560 (
      {stage1_14[3], stage1_14[4], stage1_14[5], stage1_14[6], stage1_14[7]},
      {stage1_15[12]},
      {stage1_16[1], stage1_16[2], stage1_16[3], stage1_16[4], stage1_16[5], stage1_16[6]},
      {stage2_18[1],stage2_17[2],stage2_16[2],stage2_15[3],stage2_14[6]}
   );
   gpc615_5 gpc561 (
      {stage1_14[8], stage1_14[9], stage1_14[10], stage1_14[11], stage1_14[12]},
      {1'b0},
      {stage1_16[7], stage1_16[8], stage1_16[9], stage1_16[10], stage1_16[11], stage1_16[12]},
      {stage2_18[2],stage2_17[3],stage2_16[3],stage2_15[4],stage2_14[7]}
   );
   gpc606_5 gpc562 (
      {stage1_16[13], stage1_16[14], stage1_16[15], stage1_16[16], stage1_16[17], stage1_16[18]},
      {stage1_18[0], stage1_18[1], stage1_18[2], stage1_18[3], stage1_18[4], stage1_18[5]},
      {stage2_20[0],stage2_19[0],stage2_18[3],stage2_17[4],stage2_16[4]}
   );
   gpc606_5 gpc563 (
      {stage1_16[19], stage1_16[20], stage1_16[21], stage1_16[22], stage1_16[23], stage1_16[24]},
      {stage1_18[6], stage1_18[7], stage1_18[8], stage1_18[9], stage1_18[10], 1'b0},
      {stage2_20[1],stage2_19[1],stage2_18[4],stage2_17[5],stage2_16[5]}
   );
   gpc606_5 gpc564 (
      {stage1_17[1], stage1_17[2], stage1_17[3], stage1_17[4], stage1_17[5], stage1_17[6]},
      {stage1_19[0], stage1_19[1], stage1_19[2], stage1_19[3], stage1_19[4], stage1_19[5]},
      {stage2_21[0],stage2_20[2],stage2_19[2],stage2_18[5],stage2_17[6]}
   );
   gpc606_5 gpc565 (
      {stage1_17[7], stage1_17[8], stage1_17[9], stage1_17[10], stage1_17[11], stage1_17[12]},
      {stage1_19[6], stage1_19[7], stage1_19[8], stage1_19[9], stage1_19[10], stage1_19[11]},
      {stage2_21[1],stage2_20[3],stage2_19[3],stage2_18[6],stage2_17[7]}
   );
   gpc606_5 gpc566 (
      {stage1_17[13], stage1_17[14], stage1_17[15], stage1_17[16], stage1_17[17], stage1_17[18]},
      {stage1_19[12], stage1_19[13], stage1_19[14], stage1_19[15], stage1_19[16], stage1_19[17]},
      {stage2_21[2],stage2_20[4],stage2_19[4],stage2_18[7],stage2_17[8]}
   );
   gpc1163_5 gpc567 (
      {stage1_20[0], stage1_20[1], stage1_20[2]},
      {stage1_21[0], stage1_21[1], stage1_21[2], stage1_21[3], stage1_21[4], stage1_21[5]},
      {stage1_22[0]},
      {stage1_23[0]},
      {stage2_24[0],stage2_23[0],stage2_22[0],stage2_21[3],stage2_20[5]}
   );
   gpc1163_5 gpc568 (
      {stage1_20[3], stage1_20[4], stage1_20[5]},
      {stage1_21[6], stage1_21[7], stage1_21[8], stage1_21[9], stage1_21[10], stage1_21[11]},
      {stage1_22[1]},
      {stage1_23[1]},
      {stage2_24[1],stage2_23[1],stage2_22[1],stage2_21[4],stage2_20[6]}
   );
   gpc606_5 gpc569 (
      {stage1_20[6], stage1_20[7], stage1_20[8], stage1_20[9], stage1_20[10], stage1_20[11]},
      {stage1_22[2], stage1_22[3], stage1_22[4], stage1_22[5], stage1_22[6], stage1_22[7]},
      {stage2_24[2],stage2_23[2],stage2_22[2],stage2_21[5],stage2_20[7]}
   );
   gpc606_5 gpc570 (
      {stage1_21[12], stage1_21[13], stage1_21[14], stage1_21[15], stage1_21[16], stage1_21[17]},
      {stage1_23[2], stage1_23[3], stage1_23[4], stage1_23[5], stage1_23[6], stage1_23[7]},
      {stage2_25[0],stage2_24[3],stage2_23[3],stage2_22[3],stage2_21[6]}
   );
   gpc615_5 gpc571 (
      {stage1_23[8], stage1_23[9], stage1_23[10], stage1_23[11], stage1_23[12]},
      {stage1_24[0]},
      {stage1_25[0], stage1_25[1], stage1_25[2], stage1_25[3], stage1_25[4], stage1_25[5]},
      {stage2_27[0],stage2_26[0],stage2_25[1],stage2_24[4],stage2_23[4]}
   );
   gpc615_5 gpc572 (
      {stage1_23[13], stage1_23[14], stage1_23[15], stage1_23[16], stage1_23[17]},
      {stage1_24[1]},
      {stage1_25[6], stage1_25[7], stage1_25[8], stage1_25[9], stage1_25[10], stage1_25[11]},
      {stage2_27[1],stage2_26[1],stage2_25[2],stage2_24[5],stage2_23[5]}
   );
   gpc615_5 gpc573 (
      {stage1_24[2], stage1_24[3], stage1_24[4], stage1_24[5], stage1_24[6]},
      {stage1_25[12]},
      {stage1_26[0], stage1_26[1], stage1_26[2], stage1_26[3], stage1_26[4], stage1_26[5]},
      {stage2_28[0],stage2_27[2],stage2_26[2],stage2_25[3],stage2_24[6]}
   );
   gpc615_5 gpc574 (
      {stage1_24[7], stage1_24[8], stage1_24[9], stage1_24[10], stage1_24[11]},
      {stage1_25[13]},
      {stage1_26[6], stage1_26[7], stage1_26[8], stage1_26[9], stage1_26[10], stage1_26[11]},
      {stage2_28[1],stage2_27[3],stage2_26[3],stage2_25[4],stage2_24[7]}
   );
   gpc606_5 gpc575 (
      {stage1_25[14], stage1_25[15], stage1_25[16], stage1_25[17], 1'b0, 1'b0},
      {stage1_27[0], stage1_27[1], stage1_27[2], stage1_27[3], stage1_27[4], stage1_27[5]},
      {stage2_29[0],stage2_28[2],stage2_27[4],stage2_26[4],stage2_25[5]}
   );
   gpc615_5 gpc576 (
      {stage1_26[12], stage1_26[13], stage1_26[14], stage1_26[15], stage1_26[16]},
      {stage1_27[6]},
      {stage1_28[0], stage1_28[1], stage1_28[2], stage1_28[3], stage1_28[4], stage1_28[5]},
      {stage2_30[0],stage2_29[1],stage2_28[3],stage2_27[5],stage2_26[5]}
   );
   gpc615_5 gpc577 (
      {stage1_27[7], stage1_27[8], stage1_27[9], stage1_27[10], 1'b0},
      {stage1_28[6]},
      {stage1_29[0], stage1_29[1], stage1_29[2], stage1_29[3], stage1_29[4], stage1_29[5]},
      {stage2_31[0],stage2_30[1],stage2_29[2],stage2_28[4],stage2_27[6]}
   );
   gpc606_5 gpc578 (
      {stage1_28[7], stage1_28[8], stage1_28[9], stage1_28[10], stage1_28[11], stage1_28[12]},
      {stage1_30[0], stage1_30[1], stage1_30[2], stage1_30[3], stage1_30[4], stage1_30[5]},
      {stage2_32[0],stage2_31[1],stage2_30[2],stage2_29[3],stage2_28[5]}
   );
   gpc606_5 gpc579 (
      {stage1_29[6], stage1_29[7], stage1_29[8], stage1_29[9], stage1_29[10], stage1_29[11]},
      {stage1_31[0], stage1_31[1], stage1_31[2], stage1_31[3], stage1_31[4], stage1_31[5]},
      {stage2_33[0],stage2_32[1],stage2_31[2],stage2_30[3],stage2_29[4]}
   );
   gpc606_5 gpc580 (
      {stage1_29[12], stage1_29[13], stage1_29[14], stage1_29[15], stage1_29[16], stage1_29[17]},
      {stage1_31[6], stage1_31[7], stage1_31[8], stage1_31[9], stage1_31[10], stage1_31[11]},
      {stage2_33[1],stage2_32[2],stage2_31[3],stage2_30[4],stage2_29[5]}
   );
   gpc615_5 gpc581 (
      {stage1_30[6], stage1_30[7], stage1_30[8], stage1_30[9], stage1_30[10]},
      {stage1_31[12]},
      {stage1_32[0], stage1_32[1], stage1_32[2], stage1_32[3], stage1_32[4], stage1_32[5]},
      {stage2_34[0],stage2_33[2],stage2_32[3],stage2_31[4],stage2_30[5]}
   );
   gpc1406_5 gpc582 (
      {stage1_32[6], stage1_32[7], stage1_32[8], stage1_32[9], stage1_32[10], stage1_32[11]},
      {stage1_34[0], stage1_34[1], stage1_34[2], stage1_34[3]},
      {stage1_35[0]},
      {stage2_36[0],stage2_35[0],stage2_34[1],stage2_33[3],stage2_32[4]}
   );
   gpc1406_5 gpc583 (
      {stage1_32[12], stage1_32[13], stage1_32[14], stage1_32[15], stage1_32[16], stage1_32[17]},
      {stage1_34[4], stage1_34[5], stage1_34[6], stage1_34[7]},
      {stage1_35[1]},
      {stage2_36[1],stage2_35[1],stage2_34[2],stage2_33[4],stage2_32[5]}
   );
   gpc606_5 gpc584 (
      {stage1_32[18], stage1_32[19], stage1_32[20], stage1_32[21], stage1_32[22], stage1_32[23]},
      {stage1_34[8], stage1_34[9], stage1_34[10], stage1_34[11], stage1_34[12], stage1_34[13]},
      {stage2_36[2],stage2_35[2],stage2_34[3],stage2_33[5],stage2_32[6]}
   );
   gpc615_5 gpc585 (
      {stage1_33[0], stage1_33[1], stage1_33[2], stage1_33[3], stage1_33[4]},
      {stage1_34[14]},
      {stage1_35[2], stage1_35[3], stage1_35[4], stage1_35[5], stage1_35[6], stage1_35[7]},
      {stage2_37[0],stage2_36[3],stage2_35[3],stage2_34[4],stage2_33[6]}
   );
   gpc615_5 gpc586 (
      {stage1_33[5], stage1_33[6], stage1_33[7], stage1_33[8], stage1_33[9]},
      {stage1_34[15]},
      {stage1_35[8], stage1_35[9], stage1_35[10], stage1_35[11], stage1_35[12], 1'b0},
      {stage2_37[1],stage2_36[4],stage2_35[4],stage2_34[5],stage2_33[7]}
   );
   gpc615_5 gpc587 (
      {stage1_34[16], stage1_34[17], stage1_34[18], stage1_34[19], stage1_34[20]},
      {1'b0},
      {stage1_36[0], stage1_36[1], stage1_36[2], stage1_36[3], stage1_36[4], stage1_36[5]},
      {stage2_38[0],stage2_37[2],stage2_36[5],stage2_35[5],stage2_34[6]}
   );
   gpc606_5 gpc588 (
      {stage1_36[6], stage1_36[7], stage1_36[8], stage1_36[9], stage1_36[10], stage1_36[11]},
      {stage1_38[0], stage1_38[1], stage1_38[2], stage1_38[3], stage1_38[4], stage1_38[5]},
      {stage2_40[0],stage2_39[0],stage2_38[1],stage2_37[3],stage2_36[6]}
   );
   gpc615_5 gpc589 (
      {stage1_37[0], stage1_37[1], stage1_37[2], stage1_37[3], stage1_37[4]},
      {stage1_38[6]},
      {stage1_39[0], stage1_39[1], stage1_39[2], stage1_39[3], stage1_39[4], stage1_39[5]},
      {stage2_41[0],stage2_40[1],stage2_39[1],stage2_38[2],stage2_37[4]}
   );
   gpc606_5 gpc590 (
      {stage1_38[7], stage1_38[8], stage1_38[9], stage1_38[10], stage1_38[11], stage1_38[12]},
      {stage1_40[0], stage1_40[1], stage1_40[2], stage1_40[3], stage1_40[4], stage1_40[5]},
      {stage2_42[0],stage2_41[1],stage2_40[2],stage2_39[2],stage2_38[3]}
   );
   gpc615_5 gpc591 (
      {stage1_38[13], stage1_38[14], stage1_38[15], stage1_38[16], stage1_38[17]},
      {stage1_39[6]},
      {stage1_40[6], stage1_40[7], stage1_40[8], stage1_40[9], stage1_40[10], stage1_40[11]},
      {stage2_42[1],stage2_41[2],stage2_40[3],stage2_39[3],stage2_38[4]}
   );
   gpc606_5 gpc592 (
      {stage1_39[7], stage1_39[8], stage1_39[9], stage1_39[10], stage1_39[11], stage1_39[12]},
      {stage1_41[0], stage1_41[1], stage1_41[2], stage1_41[3], stage1_41[4], stage1_41[5]},
      {stage2_43[0],stage2_42[2],stage2_41[3],stage2_40[4],stage2_39[4]}
   );
   gpc606_5 gpc593 (
      {stage1_40[12], stage1_40[13], stage1_40[14], stage1_40[15], 1'b0, 1'b0},
      {stage1_42[0], stage1_42[1], stage1_42[2], stage1_42[3], stage1_42[4], stage1_42[5]},
      {stage2_44[0],stage2_43[1],stage2_42[3],stage2_41[4],stage2_40[5]}
   );
   gpc117_4 gpc594 (
      {stage1_41[6], stage1_41[7], stage1_41[8], stage1_41[9], stage1_41[10], stage1_41[11], stage1_41[12]},
      {stage1_42[6]},
      {stage1_43[0]},
      {stage2_44[1],stage2_43[2],stage2_42[4],stage2_41[5]}
   );
   gpc117_4 gpc595 (
      {stage1_41[13], stage1_41[14], stage1_41[15], stage1_41[16], stage1_41[17], stage1_41[18], stage1_41[19]},
      {stage1_42[7]},
      {stage1_43[1]},
      {stage2_44[2],stage2_43[3],stage2_42[5],stage2_41[6]}
   );
   gpc606_5 gpc596 (
      {stage1_43[2], stage1_43[3], stage1_43[4], stage1_43[5], stage1_43[6], stage1_43[7]},
      {stage1_45[0], stage1_45[1], stage1_45[2], stage1_45[3], stage1_45[4], stage1_45[5]},
      {stage2_47[0],stage2_46[0],stage2_45[0],stage2_44[3],stage2_43[4]}
   );
   gpc615_5 gpc597 (
      {stage1_43[8], stage1_43[9], stage1_43[10], stage1_43[11], stage1_43[12]},
      {stage1_44[0]},
      {stage1_45[6], stage1_45[7], stage1_45[8], stage1_45[9], stage1_45[10], stage1_45[11]},
      {stage2_47[1],stage2_46[1],stage2_45[1],stage2_44[4],stage2_43[5]}
   );
   gpc606_5 gpc598 (
      {stage1_45[12], stage1_45[13], stage1_45[14], stage1_45[15], stage1_45[16], stage1_45[17]},
      {stage1_47[0], stage1_47[1], stage1_47[2], stage1_47[3], stage1_47[4], stage1_47[5]},
      {stage2_49[0],stage2_48[0],stage2_47[2],stage2_46[2],stage2_45[2]}
   );
   gpc606_5 gpc599 (
      {stage1_45[18], stage1_45[19], stage1_45[20], stage1_45[21], stage1_45[22], stage1_45[23]},
      {stage1_47[6], stage1_47[7], stage1_47[8], stage1_47[9], stage1_47[10], stage1_47[11]},
      {stage2_49[1],stage2_48[1],stage2_47[3],stage2_46[3],stage2_45[3]}
   );
   gpc615_5 gpc600 (
      {stage1_46[0], stage1_46[1], stage1_46[2], stage1_46[3], stage1_46[4]},
      {stage1_47[12]},
      {stage1_48[0], stage1_48[1], stage1_48[2], stage1_48[3], stage1_48[4], stage1_48[5]},
      {stage2_50[0],stage2_49[2],stage2_48[2],stage2_47[4],stage2_46[4]}
   );
   gpc615_5 gpc601 (
      {stage1_46[5], stage1_46[6], stage1_46[7], stage1_46[8], stage1_46[9]},
      {stage1_47[13]},
      {stage1_48[6], stage1_48[7], stage1_48[8], stage1_48[9], stage1_48[10], stage1_48[11]},
      {stage2_50[1],stage2_49[3],stage2_48[3],stage2_47[5],stage2_46[5]}
   );
   gpc606_5 gpc602 (
      {stage1_48[12], stage1_48[13], stage1_48[14], stage1_48[15], stage1_48[16], stage1_48[17]},
      {stage1_50[0], stage1_50[1], stage1_50[2], stage1_50[3], stage1_50[4], stage1_50[5]},
      {stage2_52[0],stage2_51[0],stage2_50[2],stage2_49[4],stage2_48[4]}
   );
   gpc606_5 gpc603 (
      {stage1_49[0], stage1_49[1], stage1_49[2], stage1_49[3], stage1_49[4], stage1_49[5]},
      {stage1_51[0], stage1_51[1], stage1_51[2], stage1_51[3], stage1_51[4], stage1_51[5]},
      {stage2_53[0],stage2_52[1],stage2_51[1],stage2_50[3],stage2_49[5]}
   );
   gpc615_5 gpc604 (
      {stage1_49[6], stage1_49[7], stage1_49[8], stage1_49[9], stage1_49[10]},
      {stage1_50[6]},
      {stage1_51[6], stage1_51[7], stage1_51[8], stage1_51[9], stage1_51[10], stage1_51[11]},
      {stage2_53[1],stage2_52[2],stage2_51[2],stage2_50[4],stage2_49[6]}
   );
   gpc615_5 gpc605 (
      {stage1_49[11], stage1_49[12], stage1_49[13], stage1_49[14], stage1_49[15]},
      {stage1_50[7]},
      {stage1_51[12], stage1_51[13], stage1_51[14], stage1_51[15], stage1_51[16], stage1_51[17]},
      {stage2_53[2],stage2_52[3],stage2_51[3],stage2_50[5],stage2_49[7]}
   );
   gpc615_5 gpc606 (
      {stage1_50[8], stage1_50[9], stage1_50[10], stage1_50[11], 1'b0},
      {stage1_51[18]},
      {stage1_52[0], stage1_52[1], stage1_52[2], stage1_52[3], stage1_52[4], stage1_52[5]},
      {stage2_54[0],stage2_53[3],stage2_52[4],stage2_51[4],stage2_50[6]}
   );
   gpc1163_5 gpc607 (
      {stage1_51[19], stage1_51[20], 1'b0},
      {stage1_52[6], stage1_52[7], stage1_52[8], stage1_52[9], stage1_52[10], stage1_52[11]},
      {stage1_53[0]},
      {stage1_54[0]},
      {stage2_55[0],stage2_54[1],stage2_53[4],stage2_52[5],stage2_51[5]}
   );
   gpc615_5 gpc608 (
      {stage1_53[1], stage1_53[2], stage1_53[3], stage1_53[4], stage1_53[5]},
      {stage1_54[1]},
      {stage1_55[0], stage1_55[1], stage1_55[2], stage1_55[3], stage1_55[4], stage1_55[5]},
      {stage2_57[0],stage2_56[0],stage2_55[1],stage2_54[2],stage2_53[5]}
   );
   gpc615_5 gpc609 (
      {stage1_53[6], stage1_53[7], stage1_53[8], stage1_53[9], stage1_53[10]},
      {stage1_54[2]},
      {stage1_55[6], stage1_55[7], stage1_55[8], stage1_55[9], stage1_55[10], stage1_55[11]},
      {stage2_57[1],stage2_56[1],stage2_55[2],stage2_54[3],stage2_53[6]}
   );
   gpc615_5 gpc610 (
      {stage1_53[11], stage1_53[12], stage1_53[13], stage1_53[14], stage1_53[15]},
      {stage1_54[3]},
      {stage1_55[12], stage1_55[13], stage1_55[14], stage1_55[15], stage1_55[16], stage1_55[17]},
      {stage2_57[2],stage2_56[2],stage2_55[3],stage2_54[4],stage2_53[7]}
   );
   gpc615_5 gpc611 (
      {stage1_53[16], stage1_53[17], stage1_53[18], stage1_53[19], stage1_53[20]},
      {stage1_54[4]},
      {stage1_55[18], stage1_55[19], stage1_55[20], stage1_55[21], stage1_55[22], stage1_55[23]},
      {stage2_57[3],stage2_56[3],stage2_55[4],stage2_54[5],stage2_53[8]}
   );
   gpc615_5 gpc612 (
      {stage1_54[5], stage1_54[6], stage1_54[7], stage1_54[8], stage1_54[9]},
      {stage1_55[24]},
      {stage1_56[0], stage1_56[1], stage1_56[2], stage1_56[3], stage1_56[4], stage1_56[5]},
      {stage2_58[0],stage2_57[4],stage2_56[4],stage2_55[5],stage2_54[6]}
   );
   gpc615_5 gpc613 (
      {stage1_55[25], stage1_55[26], stage1_55[27], stage1_55[28], stage1_55[29]},
      {stage1_56[6]},
      {stage1_57[0], stage1_57[1], stage1_57[2], stage1_57[3], stage1_57[4], stage1_57[5]},
      {stage2_59[0],stage2_58[1],stage2_57[5],stage2_56[5],stage2_55[6]}
   );
   gpc615_5 gpc614 (
      {stage1_56[7], stage1_56[8], stage1_56[9], stage1_56[10], stage1_56[11]},
      {stage1_57[6]},
      {stage1_58[0], stage1_58[1], stage1_58[2], stage1_58[3], stage1_58[4], stage1_58[5]},
      {stage2_60[0],stage2_59[1],stage2_58[2],stage2_57[6],stage2_56[6]}
   );
   gpc615_5 gpc615 (
      {stage1_57[7], stage1_57[8], stage1_57[9], stage1_57[10], stage1_57[11]},
      {stage1_58[6]},
      {stage1_59[0], stage1_59[1], stage1_59[2], stage1_59[3], stage1_59[4], stage1_59[5]},
      {stage2_61[0],stage2_60[1],stage2_59[2],stage2_58[3],stage2_57[7]}
   );
   gpc615_5 gpc616 (
      {stage1_57[12], stage1_57[13], stage1_57[14], stage1_57[15], stage1_57[16]},
      {stage1_58[7]},
      {stage1_59[6], stage1_59[7], stage1_59[8], stage1_59[9], stage1_59[10], stage1_59[11]},
      {stage2_61[1],stage2_60[2],stage2_59[3],stage2_58[4],stage2_57[8]}
   );
   gpc606_5 gpc617 (
      {stage1_58[8], stage1_58[9], stage1_58[10], stage1_58[11], stage1_58[12], stage1_58[13]},
      {stage1_60[0], stage1_60[1], stage1_60[2], stage1_60[3], stage1_60[4], stage1_60[5]},
      {stage2_62[0],stage2_61[2],stage2_60[3],stage2_59[4],stage2_58[5]}
   );
   gpc606_5 gpc618 (
      {stage1_59[12], stage1_59[13], stage1_59[14], stage1_59[15], stage1_59[16], stage1_59[17]},
      {stage1_61[0], stage1_61[1], stage1_61[2], stage1_61[3], stage1_61[4], stage1_61[5]},
      {stage2_63[0],stage2_62[1],stage2_61[3],stage2_60[4],stage2_59[5]}
   );
   gpc606_5 gpc619 (
      {stage1_60[6], stage1_60[7], stage1_60[8], stage1_60[9], stage1_60[10], stage1_60[11]},
      {stage1_62[0], stage1_62[1], stage1_62[2], stage1_62[3], stage1_62[4], stage1_62[5]},
      {stage2_64[0],stage2_63[1],stage2_62[2],stage2_61[4],stage2_60[5]}
   );
   gpc606_5 gpc620 (
      {stage1_61[6], stage1_61[7], stage1_61[8], stage1_61[9], stage1_61[10], stage1_61[11]},
      {stage1_63[0], stage1_63[1], stage1_63[2], stage1_63[3], stage1_63[4], stage1_63[5]},
      {stage2_65[0],stage2_64[1],stage2_63[2],stage2_62[3],stage2_61[5]}
   );
   gpc207_4 gpc621 (
      {stage1_62[6], stage1_62[7], stage1_62[8], stage1_62[9], stage1_62[10], stage1_62[11], stage1_62[12]},
      {stage1_64[0], stage1_64[1]},
      {stage2_65[1],stage2_64[2],stage2_63[3],stage2_62[4]}
   );
   gpc606_5 gpc622 (
      {stage1_62[13], stage1_62[14], stage1_62[15], stage1_62[16], 1'b0, 1'b0},
      {stage1_64[2], stage1_64[3], stage1_64[4], stage1_64[5], stage1_64[6], stage1_64[7]},
      {stage2_66[0],stage2_65[2],stage2_64[3],stage2_63[4],stage2_62[5]}
   );
   gpc1_1 gpc623 (
      {stage1_0[0]},
      {stage2_0[0]}
   );
   gpc1_1 gpc624 (
      {stage1_0[1]},
      {stage2_0[1]}
   );
   gpc1_1 gpc625 (
      {stage1_0[2]},
      {stage2_0[2]}
   );
   gpc1_1 gpc626 (
      {stage1_0[3]},
      {stage2_0[3]}
   );
   gpc1_1 gpc627 (
      {stage1_0[4]},
      {stage2_0[4]}
   );
   gpc1_1 gpc628 (
      {stage1_0[5]},
      {stage2_0[5]}
   );
   gpc1_1 gpc629 (
      {stage1_0[6]},
      {stage2_0[6]}
   );
   gpc1_1 gpc630 (
      {stage1_0[7]},
      {stage2_0[7]}
   );
   gpc1_1 gpc631 (
      {stage1_0[8]},
      {stage2_0[8]}
   );
   gpc1_1 gpc632 (
      {stage1_0[9]},
      {stage2_0[9]}
   );
   gpc1_1 gpc633 (
      {stage1_0[10]},
      {stage2_0[10]}
   );
   gpc1_1 gpc634 (
      {stage1_1[6]},
      {stage2_1[1]}
   );
   gpc1_1 gpc635 (
      {stage1_1[7]},
      {stage2_1[2]}
   );
   gpc1_1 gpc636 (
      {stage1_2[21]},
      {stage2_2[5]}
   );
   gpc1_1 gpc637 (
      {stage1_2[22]},
      {stage2_2[6]}
   );
   gpc1_1 gpc638 (
      {stage1_2[23]},
      {stage2_2[7]}
   );
   gpc1_1 gpc639 (
      {stage1_2[24]},
      {stage2_2[8]}
   );
   gpc1_1 gpc640 (
      {stage1_3[14]},
      {stage2_3[6]}
   );
   gpc1_1 gpc641 (
      {stage1_3[15]},
      {stage2_3[7]}
   );
   gpc1_1 gpc642 (
      {stage1_3[16]},
      {stage2_3[8]}
   );
   gpc1_1 gpc643 (
      {stage1_5[12]},
      {stage2_5[8]}
   );
   gpc1_1 gpc644 (
      {stage1_5[13]},
      {stage2_5[9]}
   );
   gpc1_1 gpc645 (
      {stage1_6[21]},
      {stage2_6[10]}
   );
   gpc1_1 gpc646 (
      {stage1_6[22]},
      {stage2_6[11]}
   );
   gpc1_1 gpc647 (
      {stage1_6[23]},
      {stage2_6[12]}
   );
   gpc1_1 gpc648 (
      {stage1_6[24]},
      {stage2_6[13]}
   );
   gpc1_1 gpc649 (
      {stage1_6[25]},
      {stage2_6[14]}
   );
   gpc1_1 gpc650 (
      {stage1_6[26]},
      {stage2_6[15]}
   );
   gpc1_1 gpc651 (
      {stage1_6[27]},
      {stage2_6[16]}
   );
   gpc1_1 gpc652 (
      {stage1_6[28]},
      {stage2_6[17]}
   );
   gpc1_1 gpc653 (
      {stage1_8[18]},
      {stage2_8[5]}
   );
   gpc1_1 gpc654 (
      {stage1_9[12]},
      {stage2_9[6]}
   );
   gpc1_1 gpc655 (
      {stage1_9[13]},
      {stage2_9[7]}
   );
   gpc1_1 gpc656 (
      {stage1_9[14]},
      {stage2_9[8]}
   );
   gpc1_1 gpc657 (
      {stage1_9[15]},
      {stage2_9[9]}
   );
   gpc1_1 gpc658 (
      {stage1_13[12]},
      {stage2_13[7]}
   );
   gpc1_1 gpc659 (
      {stage1_13[13]},
      {stage2_13[8]}
   );
   gpc1_1 gpc660 (
      {stage1_14[13]},
      {stage2_14[8]}
   );
   gpc1_1 gpc661 (
      {stage1_14[14]},
      {stage2_14[9]}
   );
   gpc1_1 gpc662 (
      {stage1_14[15]},
      {stage2_14[10]}
   );
   gpc1_1 gpc663 (
      {stage1_14[16]},
      {stage2_14[11]}
   );
   gpc1_1 gpc664 (
      {stage1_16[25]},
      {stage2_16[6]}
   );
   gpc1_1 gpc665 (
      {stage1_16[26]},
      {stage2_16[7]}
   );
   gpc1_1 gpc666 (
      {stage1_16[27]},
      {stage2_16[8]}
   );
   gpc1_1 gpc667 (
      {stage1_16[28]},
      {stage2_16[9]}
   );
   gpc1_1 gpc668 (
      {stage1_16[29]},
      {stage2_16[10]}
   );
   gpc1_1 gpc669 (
      {stage1_16[30]},
      {stage2_16[11]}
   );
   gpc1_1 gpc670 (
      {stage1_17[19]},
      {stage2_17[9]}
   );
   gpc1_1 gpc671 (
      {stage1_17[20]},
      {stage2_17[10]}
   );
   gpc1_1 gpc672 (
      {stage1_17[21]},
      {stage2_17[11]}
   );
   gpc1_1 gpc673 (
      {stage1_19[18]},
      {stage2_19[5]}
   );
   gpc1_1 gpc674 (
      {stage1_22[8]},
      {stage2_22[4]}
   );
   gpc1_1 gpc675 (
      {stage1_22[9]},
      {stage2_22[5]}
   );
   gpc1_1 gpc676 (
      {stage1_22[10]},
      {stage2_22[6]}
   );
   gpc1_1 gpc677 (
      {stage1_22[11]},
      {stage2_22[7]}
   );
   gpc1_1 gpc678 (
      {stage1_22[12]},
      {stage2_22[8]}
   );
   gpc1_1 gpc679 (
      {stage1_22[13]},
      {stage2_22[9]}
   );
   gpc1_1 gpc680 (
      {stage1_28[13]},
      {stage2_28[6]}
   );
   gpc1_1 gpc681 (
      {stage1_28[14]},
      {stage2_28[7]}
   );
   gpc1_1 gpc682 (
      {stage1_28[15]},
      {stage2_28[8]}
   );
   gpc1_1 gpc683 (
      {stage1_31[13]},
      {stage2_31[5]}
   );
   gpc1_1 gpc684 (
      {stage1_31[14]},
      {stage2_31[6]}
   );
   gpc1_1 gpc685 (
      {stage1_31[15]},
      {stage2_31[7]}
   );
   gpc1_1 gpc686 (
      {stage1_31[16]},
      {stage2_31[8]}
   );
   gpc1_1 gpc687 (
      {stage1_32[24]},
      {stage2_32[7]}
   );
   gpc1_1 gpc688 (
      {stage1_33[10]},
      {stage2_33[8]}
   );
   gpc1_1 gpc689 (
      {stage1_33[11]},
      {stage2_33[9]}
   );
   gpc1_1 gpc690 (
      {stage1_33[12]},
      {stage2_33[10]}
   );
   gpc1_1 gpc691 (
      {stage1_33[13]},
      {stage2_33[11]}
   );
   gpc1_1 gpc692 (
      {stage1_33[14]},
      {stage2_33[12]}
   );
   gpc1_1 gpc693 (
      {stage1_33[15]},
      {stage2_33[13]}
   );
   gpc1_1 gpc694 (
      {stage1_33[16]},
      {stage2_33[14]}
   );
   gpc1_1 gpc695 (
      {stage1_33[17]},
      {stage2_33[15]}
   );
   gpc1_1 gpc696 (
      {stage1_33[18]},
      {stage2_33[16]}
   );
   gpc1_1 gpc697 (
      {stage1_36[12]},
      {stage2_36[7]}
   );
   gpc1_1 gpc698 (
      {stage1_37[5]},
      {stage2_37[5]}
   );
   gpc1_1 gpc699 (
      {stage1_37[6]},
      {stage2_37[6]}
   );
   gpc1_1 gpc700 (
      {stage1_37[7]},
      {stage2_37[7]}
   );
   gpc1_1 gpc701 (
      {stage1_37[8]},
      {stage2_37[8]}
   );
   gpc1_1 gpc702 (
      {stage1_37[9]},
      {stage2_37[9]}
   );
   gpc1_1 gpc703 (
      {stage1_37[10]},
      {stage2_37[10]}
   );
   gpc1_1 gpc704 (
      {stage1_37[11]},
      {stage2_37[11]}
   );
   gpc1_1 gpc705 (
      {stage1_37[12]},
      {stage2_37[12]}
   );
   gpc1_1 gpc706 (
      {stage1_37[13]},
      {stage2_37[13]}
   );
   gpc1_1 gpc707 (
      {stage1_39[13]},
      {stage2_39[5]}
   );
   gpc1_1 gpc708 (
      {stage1_39[14]},
      {stage2_39[6]}
   );
   gpc1_1 gpc709 (
      {stage1_42[8]},
      {stage2_42[6]}
   );
   gpc1_1 gpc710 (
      {stage1_42[9]},
      {stage2_42[7]}
   );
   gpc1_1 gpc711 (
      {stage1_42[10]},
      {stage2_42[8]}
   );
   gpc1_1 gpc712 (
      {stage1_42[11]},
      {stage2_42[9]}
   );
   gpc1_1 gpc713 (
      {stage1_42[12]},
      {stage2_42[10]}
   );
   gpc1_1 gpc714 (
      {stage1_43[13]},
      {stage2_43[6]}
   );
   gpc1_1 gpc715 (
      {stage1_44[1]},
      {stage2_44[5]}
   );
   gpc1_1 gpc716 (
      {stage1_44[2]},
      {stage2_44[6]}
   );
   gpc1_1 gpc717 (
      {stage1_44[3]},
      {stage2_44[7]}
   );
   gpc1_1 gpc718 (
      {stage1_44[4]},
      {stage2_44[8]}
   );
   gpc1_1 gpc719 (
      {stage1_44[5]},
      {stage2_44[9]}
   );
   gpc1_1 gpc720 (
      {stage1_44[6]},
      {stage2_44[10]}
   );
   gpc1_1 gpc721 (
      {stage1_44[7]},
      {stage2_44[11]}
   );
   gpc1_1 gpc722 (
      {stage1_44[8]},
      {stage2_44[12]}
   );
   gpc1_1 gpc723 (
      {stage1_44[9]},
      {stage2_44[13]}
   );
   gpc1_1 gpc724 (
      {stage1_44[10]},
      {stage2_44[14]}
   );
   gpc1_1 gpc725 (
      {stage1_44[11]},
      {stage2_44[15]}
   );
   gpc1_1 gpc726 (
      {stage1_44[12]},
      {stage2_44[16]}
   );
   gpc1_1 gpc727 (
      {stage1_44[13]},
      {stage2_44[17]}
   );
   gpc1_1 gpc728 (
      {stage1_45[24]},
      {stage2_45[4]}
   );
   gpc1_1 gpc729 (
      {stage1_46[10]},
      {stage2_46[6]}
   );
   gpc1_1 gpc730 (
      {stage1_46[11]},
      {stage2_46[7]}
   );
   gpc1_1 gpc731 (
      {stage1_47[14]},
      {stage2_47[6]}
   );
   gpc1_1 gpc732 (
      {stage1_47[15]},
      {stage2_47[7]}
   );
   gpc1_1 gpc733 (
      {stage1_47[16]},
      {stage2_47[8]}
   );
   gpc1_1 gpc734 (
      {stage1_47[17]},
      {stage2_47[9]}
   );
   gpc1_1 gpc735 (
      {stage1_48[18]},
      {stage2_48[5]}
   );
   gpc1_1 gpc736 (
      {stage1_48[19]},
      {stage2_48[6]}
   );
   gpc1_1 gpc737 (
      {stage1_49[16]},
      {stage2_49[8]}
   );
   gpc1_1 gpc738 (
      {stage1_49[17]},
      {stage2_49[9]}
   );
   gpc1_1 gpc739 (
      {stage1_49[18]},
      {stage2_49[10]}
   );
   gpc1_1 gpc740 (
      {stage1_49[19]},
      {stage2_49[11]}
   );
   gpc1_1 gpc741 (
      {stage1_53[21]},
      {stage2_53[9]}
   );
   gpc1_1 gpc742 (
      {stage1_53[22]},
      {stage2_53[10]}
   );
   gpc1_1 gpc743 (
      {stage1_56[12]},
      {stage2_56[7]}
   );
   gpc1_1 gpc744 (
      {stage1_56[13]},
      {stage2_56[8]}
   );
   gpc1_1 gpc745 (
      {stage1_56[14]},
      {stage2_56[9]}
   );
   gpc1_1 gpc746 (
      {stage1_59[18]},
      {stage2_59[6]}
   );
   gpc1_1 gpc747 (
      {stage1_59[19]},
      {stage2_59[7]}
   );
   gpc1_1 gpc748 (
      {stage1_59[20]},
      {stage2_59[8]}
   );
   gpc1_1 gpc749 (
      {stage1_59[21]},
      {stage2_59[9]}
   );
   gpc1_1 gpc750 (
      {stage1_59[22]},
      {stage2_59[10]}
   );
   gpc1_1 gpc751 (
      {stage1_59[23]},
      {stage2_59[11]}
   );
   gpc1_1 gpc752 (
      {stage1_60[12]},
      {stage2_60[6]}
   );
   gpc1_1 gpc753 (
      {stage1_61[12]},
      {stage2_61[6]}
   );
   gpc1_1 gpc754 (
      {stage1_63[6]},
      {stage2_63[5]}
   );
   gpc1_1 gpc755 (
      {stage1_63[7]},
      {stage2_63[6]}
   );
   gpc1_1 gpc756 (
      {stage1_63[8]},
      {stage2_63[7]}
   );
   gpc1_1 gpc757 (
      {stage1_63[9]},
      {stage2_63[8]}
   );
   gpc1_1 gpc758 (
      {stage1_63[10]},
      {stage2_63[9]}
   );
   gpc1_1 gpc759 (
      {stage1_64[8]},
      {stage2_64[4]}
   );
   gpc1_1 gpc760 (
      {stage1_65[0]},
      {stage2_65[3]}
   );
   gpc1_1 gpc761 (
      {stage1_65[1]},
      {stage2_65[4]}
   );
   gpc1_1 gpc762 (
      {stage1_65[2]},
      {stage2_65[5]}
   );
   gpc1_1 gpc763 (
      {stage1_65[3]},
      {stage2_65[6]}
   );
   gpc1_1 gpc764 (
      {stage1_65[4]},
      {stage2_65[7]}
   );
   gpc135_4 gpc765 (
      {stage2_0[0], stage2_0[1], stage2_0[2], stage2_0[3], stage2_0[4]},
      {stage2_1[0], stage2_1[1], stage2_1[2]},
      {stage2_2[0]},
      {stage3_3[0],stage3_2[0],stage3_1[0],stage3_0[0]}
   );
   gpc606_5 gpc766 (
      {stage2_0[5], stage2_0[6], stage2_0[7], stage2_0[8], stage2_0[9], stage2_0[10]},
      {stage2_2[1], stage2_2[2], stage2_2[3], stage2_2[4], stage2_2[5], stage2_2[6]},
      {stage3_4[0],stage3_3[1],stage3_2[1],stage3_1[1],stage3_0[1]}
   );
   gpc1343_5 gpc767 (
      {stage2_3[0], stage2_3[1], stage2_3[2]},
      {stage2_4[0], stage2_4[1], stage2_4[2], stage2_4[3]},
      {stage2_5[0], stage2_5[1], stage2_5[2]},
      {stage2_6[0]},
      {stage3_7[0],stage3_6[0],stage3_5[0],stage3_4[1],stage3_3[2]}
   );
   gpc615_5 gpc768 (
      {stage2_3[3], stage2_3[4], stage2_3[5], stage2_3[6], stage2_3[7]},
      {stage2_4[4]},
      {stage2_5[3], stage2_5[4], stage2_5[5], stage2_5[6], stage2_5[7], stage2_5[8]},
      {stage3_7[1],stage3_6[1],stage3_5[1],stage3_4[2],stage3_3[3]}
   );
   gpc2135_5 gpc769 (
      {stage2_6[1], stage2_6[2], stage2_6[3], stage2_6[4], stage2_6[5]},
      {stage2_7[0], stage2_7[1], stage2_7[2]},
      {stage2_8[0]},
      {stage2_9[0], stage2_9[1]},
      {stage3_10[0],stage3_9[0],stage3_8[0],stage3_7[2],stage3_6[2]}
   );
   gpc2135_5 gpc770 (
      {stage2_6[6], stage2_6[7], stage2_6[8], stage2_6[9], stage2_6[10]},
      {stage2_7[3], stage2_7[4], stage2_7[5]},
      {stage2_8[1]},
      {stage2_9[2], stage2_9[3]},
      {stage3_10[1],stage3_9[1],stage3_8[1],stage3_7[3],stage3_6[3]}
   );
   gpc1406_5 gpc771 (
      {stage2_6[11], stage2_6[12], stage2_6[13], stage2_6[14], stage2_6[15], stage2_6[16]},
      {stage2_8[2], stage2_8[3], stage2_8[4], stage2_8[5]},
      {stage2_9[4]},
      {stage3_10[2],stage3_9[2],stage3_8[2],stage3_7[4],stage3_6[4]}
   );
   gpc615_5 gpc772 (
      {stage2_9[5], stage2_9[6], stage2_9[7], stage2_9[8], stage2_9[9]},
      {stage2_10[0]},
      {stage2_11[0], stage2_11[1], stage2_11[2], stage2_11[3], stage2_11[4], stage2_11[5]},
      {stage3_13[0],stage3_12[0],stage3_11[0],stage3_10[3],stage3_9[3]}
   );
   gpc606_5 gpc773 (
      {stage2_10[1], stage2_10[2], stage2_10[3], stage2_10[4], stage2_10[5], stage2_10[6]},
      {stage2_12[0], stage2_12[1], stage2_12[2], stage2_12[3], stage2_12[4], stage2_12[5]},
      {stage3_14[0],stage3_13[1],stage3_12[1],stage3_11[1],stage3_10[4]}
   );
   gpc7_3 gpc774 (
      {stage2_13[0], stage2_13[1], stage2_13[2], stage2_13[3], stage2_13[4], stage2_13[5], stage2_13[6]},
      {stage3_15[0],stage3_14[1],stage3_13[2]}
   );
   gpc606_5 gpc775 (
      {stage2_14[0], stage2_14[1], stage2_14[2], stage2_14[3], stage2_14[4], stage2_14[5]},
      {stage2_16[0], stage2_16[1], stage2_16[2], stage2_16[3], stage2_16[4], stage2_16[5]},
      {stage3_18[0],stage3_17[0],stage3_16[0],stage3_15[1],stage3_14[2]}
   );
   gpc606_5 gpc776 (
      {stage2_14[6], stage2_14[7], stage2_14[8], stage2_14[9], stage2_14[10], stage2_14[11]},
      {stage2_16[6], stage2_16[7], stage2_16[8], stage2_16[9], stage2_16[10], stage2_16[11]},
      {stage3_18[1],stage3_17[1],stage3_16[1],stage3_15[2],stage3_14[3]}
   );
   gpc615_5 gpc777 (
      {stage2_15[0], stage2_15[1], stage2_15[2], stage2_15[3], stage2_15[4]},
      {1'b0},
      {stage2_17[0], stage2_17[1], stage2_17[2], stage2_17[3], stage2_17[4], stage2_17[5]},
      {stage3_19[0],stage3_18[2],stage3_17[2],stage3_16[2],stage3_15[3]}
   );
   gpc606_5 gpc778 (
      {stage2_17[6], stage2_17[7], stage2_17[8], stage2_17[9], stage2_17[10], stage2_17[11]},
      {stage2_19[0], stage2_19[1], stage2_19[2], stage2_19[3], stage2_19[4], stage2_19[5]},
      {stage3_21[0],stage3_20[0],stage3_19[1],stage3_18[3],stage3_17[3]}
   );
   gpc7_3 gpc779 (
      {stage2_18[0], stage2_18[1], stage2_18[2], stage2_18[3], stage2_18[4], stage2_18[5], stage2_18[6]},
      {stage3_20[1],stage3_19[2],stage3_18[4]}
   );
   gpc606_5 gpc780 (
      {stage2_20[0], stage2_20[1], stage2_20[2], stage2_20[3], stage2_20[4], stage2_20[5]},
      {stage2_22[0], stage2_22[1], stage2_22[2], stage2_22[3], stage2_22[4], stage2_22[5]},
      {stage3_24[0],stage3_23[0],stage3_22[0],stage3_21[1],stage3_20[2]}
   );
   gpc117_4 gpc781 (
      {stage2_21[0], stage2_21[1], stage2_21[2], stage2_21[3], stage2_21[4], stage2_21[5], stage2_21[6]},
      {stage2_22[6]},
      {stage2_23[0]},
      {stage3_24[1],stage3_23[1],stage3_22[1],stage3_21[2]}
   );
   gpc615_5 gpc782 (
      {stage2_23[1], stage2_23[2], stage2_23[3], stage2_23[4], stage2_23[5]},
      {stage2_24[0]},
      {stage2_25[0], stage2_25[1], stage2_25[2], stage2_25[3], stage2_25[4], stage2_25[5]},
      {stage3_27[0],stage3_26[0],stage3_25[0],stage3_24[2],stage3_23[2]}
   );
   gpc606_5 gpc783 (
      {stage2_24[1], stage2_24[2], stage2_24[3], stage2_24[4], stage2_24[5], stage2_24[6]},
      {stage2_26[0], stage2_26[1], stage2_26[2], stage2_26[3], stage2_26[4], stage2_26[5]},
      {stage3_28[0],stage3_27[1],stage3_26[1],stage3_25[1],stage3_24[3]}
   );
   gpc615_5 gpc784 (
      {stage2_27[0], stage2_27[1], stage2_27[2], stage2_27[3], stage2_27[4]},
      {stage2_28[0]},
      {stage2_29[0], stage2_29[1], stage2_29[2], stage2_29[3], stage2_29[4], stage2_29[5]},
      {stage3_31[0],stage3_30[0],stage3_29[0],stage3_28[1],stage3_27[2]}
   );
   gpc606_5 gpc785 (
      {stage2_28[1], stage2_28[2], stage2_28[3], stage2_28[4], stage2_28[5], stage2_28[6]},
      {stage2_30[0], stage2_30[1], stage2_30[2], stage2_30[3], stage2_30[4], stage2_30[5]},
      {stage3_32[0],stage3_31[1],stage3_30[1],stage3_29[1],stage3_28[2]}
   );
   gpc615_5 gpc786 (
      {stage2_31[0], stage2_31[1], stage2_31[2], stage2_31[3], stage2_31[4]},
      {stage2_32[0]},
      {stage2_33[0], stage2_33[1], stage2_33[2], stage2_33[3], stage2_33[4], stage2_33[5]},
      {stage3_35[0],stage3_34[0],stage3_33[0],stage3_32[1],stage3_31[2]}
   );
   gpc615_5 gpc787 (
      {stage2_31[5], stage2_31[6], stage2_31[7], stage2_31[8], 1'b0},
      {stage2_32[1]},
      {stage2_33[6], stage2_33[7], stage2_33[8], stage2_33[9], stage2_33[10], stage2_33[11]},
      {stage3_35[1],stage3_34[1],stage3_33[1],stage3_32[2],stage3_31[3]}
   );
   gpc606_5 gpc788 (
      {stage2_32[2], stage2_32[3], stage2_32[4], stage2_32[5], stage2_32[6], stage2_32[7]},
      {stage2_34[0], stage2_34[1], stage2_34[2], stage2_34[3], stage2_34[4], stage2_34[5]},
      {stage3_36[0],stage3_35[2],stage3_34[2],stage3_33[2],stage3_32[3]}
   );
   gpc615_5 gpc789 (
      {stage2_33[12], stage2_33[13], stage2_33[14], stage2_33[15], stage2_33[16]},
      {stage2_34[6]},
      {stage2_35[0], stage2_35[1], stage2_35[2], stage2_35[3], stage2_35[4], stage2_35[5]},
      {stage3_37[0],stage3_36[1],stage3_35[3],stage3_34[3],stage3_33[3]}
   );
   gpc7_3 gpc790 (
      {stage2_36[0], stage2_36[1], stage2_36[2], stage2_36[3], stage2_36[4], stage2_36[5], stage2_36[6]},
      {stage3_38[0],stage3_37[1],stage3_36[2]}
   );
   gpc7_3 gpc791 (
      {stage2_37[0], stage2_37[1], stage2_37[2], stage2_37[3], stage2_37[4], stage2_37[5], stage2_37[6]},
      {stage3_39[0],stage3_38[1],stage3_37[2]}
   );
   gpc7_3 gpc792 (
      {stage2_37[7], stage2_37[8], stage2_37[9], stage2_37[10], stage2_37[11], stage2_37[12], stage2_37[13]},
      {stage3_39[1],stage3_38[2],stage3_37[3]}
   );
   gpc615_5 gpc793 (
      {stage2_38[0], stage2_38[1], stage2_38[2], stage2_38[3], stage2_38[4]},
      {stage2_39[0]},
      {stage2_40[0], stage2_40[1], stage2_40[2], stage2_40[3], stage2_40[4], stage2_40[5]},
      {stage3_42[0],stage3_41[0],stage3_40[0],stage3_39[2],stage3_38[3]}
   );
   gpc606_5 gpc794 (
      {stage2_39[1], stage2_39[2], stage2_39[3], stage2_39[4], stage2_39[5], stage2_39[6]},
      {stage2_41[0], stage2_41[1], stage2_41[2], stage2_41[3], stage2_41[4], stage2_41[5]},
      {stage3_43[0],stage3_42[1],stage3_41[1],stage3_40[1],stage3_39[3]}
   );
   gpc615_5 gpc795 (
      {stage2_42[0], stage2_42[1], stage2_42[2], stage2_42[3], stage2_42[4]},
      {stage2_43[0]},
      {stage2_44[0], stage2_44[1], stage2_44[2], stage2_44[3], stage2_44[4], stage2_44[5]},
      {stage3_46[0],stage3_45[0],stage3_44[0],stage3_43[1],stage3_42[2]}
   );
   gpc615_5 gpc796 (
      {stage2_42[5], stage2_42[6], stage2_42[7], stage2_42[8], stage2_42[9]},
      {stage2_43[1]},
      {stage2_44[6], stage2_44[7], stage2_44[8], stage2_44[9], stage2_44[10], stage2_44[11]},
      {stage3_46[1],stage3_45[1],stage3_44[1],stage3_43[2],stage3_42[3]}
   );
   gpc1325_5 gpc797 (
      {stage2_43[2], stage2_43[3], stage2_43[4], stage2_43[5], stage2_43[6]},
      {stage2_44[12], stage2_44[13]},
      {stage2_45[0], stage2_45[1], stage2_45[2]},
      {stage2_46[0]},
      {stage3_47[0],stage3_46[2],stage3_45[2],stage3_44[2],stage3_43[3]}
   );
   gpc135_4 gpc798 (
      {stage2_44[14], stage2_44[15], stage2_44[16], stage2_44[17], 1'b0},
      {stage2_45[3], stage2_45[4], 1'b0},
      {stage2_46[1]},
      {stage3_47[1],stage3_46[3],stage3_45[3],stage3_44[3]}
   );
   gpc615_5 gpc799 (
      {stage2_46[2], stage2_46[3], stage2_46[4], stage2_46[5], stage2_46[6]},
      {stage2_47[0]},
      {stage2_48[0], stage2_48[1], stage2_48[2], stage2_48[3], stage2_48[4], stage2_48[5]},
      {stage3_50[0],stage3_49[0],stage3_48[0],stage3_47[2],stage3_46[4]}
   );
   gpc615_5 gpc800 (
      {stage2_47[1], stage2_47[2], stage2_47[3], stage2_47[4], stage2_47[5]},
      {stage2_48[6]},
      {stage2_49[0], stage2_49[1], stage2_49[2], stage2_49[3], stage2_49[4], stage2_49[5]},
      {stage3_51[0],stage3_50[1],stage3_49[1],stage3_48[1],stage3_47[3]}
   );
   gpc615_5 gpc801 (
      {stage2_47[6], stage2_47[7], stage2_47[8], stage2_47[9], 1'b0},
      {1'b0},
      {stage2_49[6], stage2_49[7], stage2_49[8], stage2_49[9], stage2_49[10], stage2_49[11]},
      {stage3_51[1],stage3_50[2],stage3_49[2],stage3_48[2],stage3_47[4]}
   );
   gpc15_3 gpc802 (
      {stage2_50[0], stage2_50[1], stage2_50[2], stage2_50[3], stage2_50[4]},
      {stage2_51[0]},
      {stage3_52[0],stage3_51[2],stage3_50[3]}
   );
   gpc615_5 gpc803 (
      {stage2_51[1], stage2_51[2], stage2_51[3], stage2_51[4], stage2_51[5]},
      {stage2_52[0]},
      {stage2_53[0], stage2_53[1], stage2_53[2], stage2_53[3], stage2_53[4], stage2_53[5]},
      {stage3_55[0],stage3_54[0],stage3_53[0],stage3_52[1],stage3_51[3]}
   );
   gpc1406_5 gpc804 (
      {stage2_52[1], stage2_52[2], stage2_52[3], stage2_52[4], stage2_52[5], 1'b0},
      {stage2_54[0], stage2_54[1], stage2_54[2], stage2_54[3]},
      {stage2_55[0]},
      {stage3_56[0],stage3_55[1],stage3_54[1],stage3_53[1],stage3_52[2]}
   );
   gpc606_5 gpc805 (
      {stage2_53[6], stage2_53[7], stage2_53[8], stage2_53[9], stage2_53[10], 1'b0},
      {stage2_55[1], stage2_55[2], stage2_55[3], stage2_55[4], stage2_55[5], stage2_55[6]},
      {stage3_57[0],stage3_56[1],stage3_55[2],stage3_54[2],stage3_53[2]}
   );
   gpc135_4 gpc806 (
      {stage2_56[0], stage2_56[1], stage2_56[2], stage2_56[3], stage2_56[4]},
      {stage2_57[0], stage2_57[1], stage2_57[2]},
      {stage2_58[0]},
      {stage3_59[0],stage3_58[0],stage3_57[1],stage3_56[2]}
   );
   gpc1163_5 gpc807 (
      {stage2_56[5], stage2_56[6], stage2_56[7]},
      {stage2_57[3], stage2_57[4], stage2_57[5], stage2_57[6], stage2_57[7], stage2_57[8]},
      {stage2_58[1]},
      {stage2_59[0]},
      {stage3_60[0],stage3_59[1],stage3_58[1],stage3_57[2],stage3_56[3]}
   );
   gpc1343_5 gpc808 (
      {stage2_58[2], stage2_58[3], stage2_58[4]},
      {stage2_59[1], stage2_59[2], stage2_59[3], stage2_59[4]},
      {stage2_60[0], stage2_60[1], stage2_60[2]},
      {stage2_61[0]},
      {stage3_62[0],stage3_61[0],stage3_60[1],stage3_59[2],stage3_58[2]}
   );
   gpc2135_5 gpc809 (
      {stage2_59[5], stage2_59[6], stage2_59[7], stage2_59[8], stage2_59[9]},
      {stage2_60[3], stage2_60[4], stage2_60[5]},
      {stage2_61[1]},
      {stage2_62[0], stage2_62[1]},
      {stage3_63[0],stage3_62[1],stage3_61[1],stage3_60[2],stage3_59[3]}
   );
   gpc615_5 gpc810 (
      {stage2_61[2], stage2_61[3], stage2_61[4], stage2_61[5], stage2_61[6]},
      {stage2_62[2]},
      {stage2_63[0], stage2_63[1], stage2_63[2], stage2_63[3], stage2_63[4], stage2_63[5]},
      {stage3_65[0],stage3_64[0],stage3_63[1],stage3_62[2],stage3_61[2]}
   );
   gpc615_5 gpc811 (
      {stage2_63[6], stage2_63[7], stage2_63[8], stage2_63[9], 1'b0},
      {stage2_64[0]},
      {stage2_65[0], stage2_65[1], stage2_65[2], stage2_65[3], stage2_65[4], stage2_65[5]},
      {stage3_67[0],stage3_66[0],stage3_65[1],stage3_64[1],stage3_63[2]}
   );
   gpc1_1 gpc812 (
      {stage2_2[7]},
      {stage3_2[2]}
   );
   gpc1_1 gpc813 (
      {stage2_2[8]},
      {stage3_2[3]}
   );
   gpc1_1 gpc814 (
      {stage2_3[8]},
      {stage3_3[4]}
   );
   gpc1_1 gpc815 (
      {stage2_4[5]},
      {stage3_4[3]}
   );
   gpc1_1 gpc816 (
      {stage2_4[6]},
      {stage3_4[4]}
   );
   gpc1_1 gpc817 (
      {stage2_5[9]},
      {stage3_5[2]}
   );
   gpc1_1 gpc818 (
      {stage2_6[17]},
      {stage3_6[5]}
   );
   gpc1_1 gpc819 (
      {stage2_10[7]},
      {stage3_10[5]}
   );
   gpc1_1 gpc820 (
      {stage2_13[7]},
      {stage3_13[3]}
   );
   gpc1_1 gpc821 (
      {stage2_13[8]},
      {stage3_13[4]}
   );
   gpc1_1 gpc822 (
      {stage2_18[7]},
      {stage3_18[5]}
   );
   gpc1_1 gpc823 (
      {stage2_20[6]},
      {stage3_20[3]}
   );
   gpc1_1 gpc824 (
      {stage2_20[7]},
      {stage3_20[4]}
   );
   gpc1_1 gpc825 (
      {stage2_22[7]},
      {stage3_22[2]}
   );
   gpc1_1 gpc826 (
      {stage2_22[8]},
      {stage3_22[3]}
   );
   gpc1_1 gpc827 (
      {stage2_22[9]},
      {stage3_22[4]}
   );
   gpc1_1 gpc828 (
      {stage2_24[7]},
      {stage3_24[4]}
   );
   gpc1_1 gpc829 (
      {stage2_27[5]},
      {stage3_27[3]}
   );
   gpc1_1 gpc830 (
      {stage2_27[6]},
      {stage3_27[4]}
   );
   gpc1_1 gpc831 (
      {stage2_28[7]},
      {stage3_28[3]}
   );
   gpc1_1 gpc832 (
      {stage2_28[8]},
      {stage3_28[4]}
   );
   gpc1_1 gpc833 (
      {stage2_36[7]},
      {stage3_36[3]}
   );
   gpc1_1 gpc834 (
      {stage2_41[6]},
      {stage3_41[2]}
   );
   gpc1_1 gpc835 (
      {stage2_42[10]},
      {stage3_42[4]}
   );
   gpc1_1 gpc836 (
      {stage2_46[7]},
      {stage3_46[5]}
   );
   gpc1_1 gpc837 (
      {stage2_50[5]},
      {stage3_50[4]}
   );
   gpc1_1 gpc838 (
      {stage2_50[6]},
      {stage3_50[5]}
   );
   gpc1_1 gpc839 (
      {stage2_54[4]},
      {stage3_54[3]}
   );
   gpc1_1 gpc840 (
      {stage2_54[5]},
      {stage3_54[4]}
   );
   gpc1_1 gpc841 (
      {stage2_54[6]},
      {stage3_54[5]}
   );
   gpc1_1 gpc842 (
      {stage2_56[8]},
      {stage3_56[4]}
   );
   gpc1_1 gpc843 (
      {stage2_56[9]},
      {stage3_56[5]}
   );
   gpc1_1 gpc844 (
      {stage2_58[5]},
      {stage3_58[3]}
   );
   gpc1_1 gpc845 (
      {stage2_59[10]},
      {stage3_59[4]}
   );
   gpc1_1 gpc846 (
      {stage2_59[11]},
      {stage3_59[5]}
   );
   gpc1_1 gpc847 (
      {stage2_60[6]},
      {stage3_60[3]}
   );
   gpc1_1 gpc848 (
      {stage2_62[3]},
      {stage3_62[3]}
   );
   gpc1_1 gpc849 (
      {stage2_62[4]},
      {stage3_62[4]}
   );
   gpc1_1 gpc850 (
      {stage2_62[5]},
      {stage3_62[5]}
   );
   gpc1_1 gpc851 (
      {stage2_64[1]},
      {stage3_64[2]}
   );
   gpc1_1 gpc852 (
      {stage2_64[2]},
      {stage3_64[3]}
   );
   gpc1_1 gpc853 (
      {stage2_64[3]},
      {stage3_64[4]}
   );
   gpc1_1 gpc854 (
      {stage2_64[4]},
      {stage3_64[5]}
   );
   gpc1_1 gpc855 (
      {stage2_65[6]},
      {stage3_65[2]}
   );
   gpc1_1 gpc856 (
      {stage2_65[7]},
      {stage3_65[3]}
   );
   gpc1_1 gpc857 (
      {stage2_66[0]},
      {stage3_66[1]}
   );
   gpc1343_5 gpc858 (
      {stage3_2[0], stage3_2[1], stage3_2[2]},
      {stage3_3[0], stage3_3[1], stage3_3[2], stage3_3[3]},
      {stage3_4[0], stage3_4[1], stage3_4[2]},
      {stage3_5[0]},
      {stage4_6[0],stage4_5[0],stage4_4[0],stage4_3[0],stage4_2[0]}
   );
   gpc623_5 gpc859 (
      {stage3_4[3], stage3_4[4], 1'b0},
      {stage3_5[1], stage3_5[2]},
      {stage3_6[0], stage3_6[1], stage3_6[2], stage3_6[3], stage3_6[4], stage3_6[5]},
      {stage4_8[0],stage4_7[0],stage4_6[1],stage4_5[1],stage4_4[1]}
   );
   gpc135_4 gpc860 (
      {stage3_7[0], stage3_7[1], stage3_7[2], stage3_7[3], stage3_7[4]},
      {stage3_8[0], stage3_8[1], stage3_8[2]},
      {stage3_9[0]},
      {stage4_10[0],stage4_9[0],stage4_8[1],stage4_7[1]}
   );
   gpc1163_5 gpc861 (
      {stage3_9[1], stage3_9[2], stage3_9[3]},
      {stage3_10[0], stage3_10[1], stage3_10[2], stage3_10[3], stage3_10[4], stage3_10[5]},
      {stage3_11[0]},
      {stage3_12[0]},
      {stage4_13[0],stage4_12[0],stage4_11[0],stage4_10[1],stage4_9[1]}
   );
   gpc1163_5 gpc862 (
      {stage3_12[1], 1'b0, 1'b0},
      {stage3_13[0], stage3_13[1], stage3_13[2], stage3_13[3], stage3_13[4], 1'b0},
      {stage3_14[0]},
      {stage3_15[0]},
      {stage4_16[0],stage4_15[0],stage4_14[0],stage4_13[1],stage4_12[1]}
   );
   gpc1343_5 gpc863 (
      {stage3_14[1], stage3_14[2], stage3_14[3]},
      {stage3_15[1], stage3_15[2], stage3_15[3], 1'b0},
      {stage3_16[0], stage3_16[1], stage3_16[2]},
      {stage3_17[0]},
      {stage4_18[0],stage4_17[0],stage4_16[1],stage4_15[1],stage4_14[1]}
   );
   gpc1163_5 gpc864 (
      {stage3_17[1], stage3_17[2], stage3_17[3]},
      {stage3_18[0], stage3_18[1], stage3_18[2], stage3_18[3], stage3_18[4], stage3_18[5]},
      {stage3_19[0]},
      {stage3_20[0]},
      {stage4_21[0],stage4_20[0],stage4_19[0],stage4_18[1],stage4_17[1]}
   );
   gpc1343_5 gpc865 (
      {stage3_19[1], stage3_19[2], 1'b0},
      {stage3_20[1], stage3_20[2], stage3_20[3], stage3_20[4]},
      {stage3_21[0], stage3_21[1], stage3_21[2]},
      {stage3_22[0]},
      {stage4_23[0],stage4_22[0],stage4_21[1],stage4_20[1],stage4_19[1]}
   );
   gpc2135_5 gpc866 (
      {stage3_22[1], stage3_22[2], stage3_22[3], stage3_22[4], 1'b0},
      {stage3_23[0], stage3_23[1], stage3_23[2]},
      {stage3_24[0]},
      {stage3_25[0], stage3_25[1]},
      {stage4_26[0],stage4_25[0],stage4_24[0],stage4_23[1],stage4_22[1]}
   );
   gpc207_4 gpc867 (
      {stage3_24[1], stage3_24[2], stage3_24[3], stage3_24[4], 1'b0, 1'b0, 1'b0},
      {stage3_26[0], stage3_26[1]},
      {stage4_27[0],stage4_26[1],stage4_25[1],stage4_24[1]}
   );
   gpc207_4 gpc868 (
      {stage3_27[0], stage3_27[1], stage3_27[2], stage3_27[3], stage3_27[4], 1'b0, 1'b0},
      {stage3_29[0], stage3_29[1]},
      {stage4_30[0],stage4_29[0],stage4_28[0],stage4_27[1]}
   );
   gpc1415_5 gpc869 (
      {stage3_28[0], stage3_28[1], stage3_28[2], stage3_28[3], stage3_28[4]},
      {1'b0},
      {stage3_30[0], stage3_30[1], 1'b0, 1'b0},
      {stage3_31[0]},
      {stage4_32[0],stage4_31[0],stage4_30[1],stage4_29[1],stage4_28[1]}
   );
   gpc1343_5 gpc870 (
      {stage3_31[1], stage3_31[2], stage3_31[3]},
      {stage3_32[0], stage3_32[1], stage3_32[2], stage3_32[3]},
      {stage3_33[0], stage3_33[1], stage3_33[2]},
      {stage3_34[0]},
      {stage4_35[0],stage4_34[0],stage4_33[0],stage4_32[1],stage4_31[1]}
   );
   gpc1343_5 gpc871 (
      {stage3_34[1], stage3_34[2], stage3_34[3]},
      {stage3_35[0], stage3_35[1], stage3_35[2], stage3_35[3]},
      {stage3_36[0], stage3_36[1], stage3_36[2]},
      {stage3_37[0]},
      {stage4_38[0],stage4_37[0],stage4_36[0],stage4_35[1],stage4_34[1]}
   );
   gpc1343_5 gpc872 (
      {stage3_37[1], stage3_37[2], stage3_37[3]},
      {stage3_38[0], stage3_38[1], stage3_38[2], stage3_38[3]},
      {stage3_39[0], stage3_39[1], stage3_39[2]},
      {stage3_40[0]},
      {stage4_41[0],stage4_40[0],stage4_39[0],stage4_38[1],stage4_37[1]}
   );
   gpc1343_5 gpc873 (
      {stage3_41[0], stage3_41[1], stage3_41[2]},
      {stage3_42[0], stage3_42[1], stage3_42[2], stage3_42[3]},
      {stage3_43[0], stage3_43[1], stage3_43[2]},
      {stage3_44[0]},
      {stage4_45[0],stage4_44[0],stage4_43[0],stage4_42[0],stage4_41[1]}
   );
   gpc1343_5 gpc874 (
      {stage3_44[1], stage3_44[2], stage3_44[3]},
      {stage3_45[0], stage3_45[1], stage3_45[2], stage3_45[3]},
      {stage3_46[0], stage3_46[1], stage3_46[2]},
      {stage3_47[0]},
      {stage4_48[0],stage4_47[0],stage4_46[0],stage4_45[1],stage4_44[1]}
   );
   gpc1343_5 gpc875 (
      {stage3_46[3], stage3_46[4], stage3_46[5]},
      {stage3_47[1], stage3_47[2], stage3_47[3], stage3_47[4]},
      {stage3_48[0], stage3_48[1], stage3_48[2]},
      {stage3_49[0]},
      {stage4_50[0],stage4_49[0],stage4_48[1],stage4_47[1],stage4_46[1]}
   );
   gpc1163_5 gpc876 (
      {stage3_49[1], stage3_49[2], 1'b0},
      {stage3_50[0], stage3_50[1], stage3_50[2], stage3_50[3], stage3_50[4], stage3_50[5]},
      {stage3_51[0]},
      {stage3_52[0]},
      {stage4_53[0],stage4_52[0],stage4_51[0],stage4_50[1],stage4_49[1]}
   );
   gpc1343_5 gpc877 (
      {stage3_51[1], stage3_51[2], stage3_51[3]},
      {stage3_52[1], stage3_52[2], 1'b0, 1'b0},
      {stage3_53[0], stage3_53[1], stage3_53[2]},
      {stage3_54[0]},
      {stage4_55[0],stage4_54[0],stage4_53[1],stage4_52[1],stage4_51[1]}
   );
   gpc135_4 gpc878 (
      {stage3_54[1], stage3_54[2], stage3_54[3], stage3_54[4], stage3_54[5]},
      {stage3_55[0], stage3_55[1], stage3_55[2]},
      {stage3_56[0]},
      {stage4_57[0],stage4_56[0],stage4_55[1],stage4_54[1]}
   );
   gpc135_4 gpc879 (
      {stage3_56[1], stage3_56[2], stage3_56[3], stage3_56[4], stage3_56[5]},
      {stage3_57[0], stage3_57[1], stage3_57[2]},
      {stage3_58[0]},
      {stage4_59[0],stage4_58[0],stage4_57[1],stage4_56[1]}
   );
   gpc1163_5 gpc880 (
      {stage3_58[1], stage3_58[2], stage3_58[3]},
      {stage3_59[0], stage3_59[1], stage3_59[2], stage3_59[3], stage3_59[4], stage3_59[5]},
      {stage3_60[0]},
      {stage3_61[0]},
      {stage4_62[0],stage4_61[0],stage4_60[0],stage4_59[1],stage4_58[1]}
   );
   gpc623_5 gpc881 (
      {stage3_60[1], stage3_60[2], stage3_60[3]},
      {stage3_61[1], stage3_61[2]},
      {stage3_62[0], stage3_62[1], stage3_62[2], stage3_62[3], stage3_62[4], stage3_62[5]},
      {stage4_64[0],stage4_63[0],stage4_62[1],stage4_61[1],stage4_60[1]}
   );
   gpc1163_5 gpc882 (
      {stage3_63[0], stage3_63[1], stage3_63[2]},
      {stage3_64[0], stage3_64[1], stage3_64[2], stage3_64[3], stage3_64[4], stage3_64[5]},
      {stage3_65[0]},
      {stage3_66[0]},
      {stage4_67[0],stage4_66[0],stage4_65[0],stage4_64[1],stage4_63[1]}
   );
   gpc1415_5 gpc883 (
      {stage3_65[1], stage3_65[2], stage3_65[3], 1'b0, 1'b0},
      {stage3_66[1]},
      {stage3_67[0], 1'b0, 1'b0, 1'b0},
      {1'b0},
      {stage4_68[0],stage4_67[1],stage4_66[1],stage4_65[1]}
   );
   gpc1_1 gpc884 (
      {stage3_0[0]},
      {stage4_0[0]}
   );
   gpc1_1 gpc885 (
      {stage3_0[1]},
      {stage4_0[1]}
   );
   gpc1_1 gpc886 (
      {stage3_1[0]},
      {stage4_1[0]}
   );
   gpc1_1 gpc887 (
      {stage3_1[1]},
      {stage4_1[1]}
   );
   gpc1_1 gpc888 (
      {stage3_2[3]},
      {stage4_2[1]}
   );
   gpc1_1 gpc889 (
      {stage3_3[4]},
      {stage4_3[1]}
   );
   gpc1_1 gpc890 (
      {stage3_11[1]},
      {stage4_11[1]}
   );
   gpc1_1 gpc891 (
      {stage3_33[3]},
      {stage4_33[1]}
   );
   gpc1_1 gpc892 (
      {stage3_36[3]},
      {stage4_36[1]}
   );
   gpc1_1 gpc893 (
      {stage3_39[3]},
      {stage4_39[1]}
   );
   gpc1_1 gpc894 (
      {stage3_40[1]},
      {stage4_40[1]}
   );
   gpc1_1 gpc895 (
      {stage3_42[4]},
      {stage4_42[1]}
   );
   gpc1_1 gpc896 (
      {stage3_43[3]},
      {stage4_43[1]}
   );
endmodule

module testbench();
    reg [31:0] src0;
    reg [31:0] src1;
    reg [31:0] src2;
    reg [31:0] src3;
    reg [31:0] src4;
    reg [31:0] src5;
    reg [31:0] src6;
    reg [31:0] src7;
    reg [31:0] src8;
    reg [31:0] src9;
    reg [31:0] src10;
    reg [31:0] src11;
    reg [31:0] src12;
    reg [31:0] src13;
    reg [31:0] src14;
    reg [31:0] src15;
    reg [31:0] src16;
    reg [31:0] src17;
    reg [31:0] src18;
    reg [31:0] src19;
    reg [31:0] src20;
    reg [31:0] src21;
    reg [31:0] src22;
    reg [31:0] src23;
    reg [31:0] src24;
    reg [31:0] src25;
    reg [31:0] src26;
    reg [31:0] src27;
    reg [31:0] src28;
    reg [31:0] src29;
    reg [31:0] src30;
    reg [31:0] src31;
    reg [31:0] src32;
    reg [31:0] src33;
    reg [31:0] src34;
    reg [31:0] src35;
    reg [31:0] src36;
    reg [31:0] src37;
    reg [31:0] src38;
    reg [31:0] src39;
    reg [31:0] src40;
    reg [31:0] src41;
    reg [31:0] src42;
    reg [31:0] src43;
    reg [31:0] src44;
    reg [31:0] src45;
    reg [31:0] src46;
    reg [31:0] src47;
    reg [31:0] src48;
    reg [31:0] src49;
    reg [31:0] src50;
    reg [31:0] src51;
    reg [31:0] src52;
    reg [31:0] src53;
    reg [31:0] src54;
    reg [31:0] src55;
    reg [31:0] src56;
    reg [31:0] src57;
    reg [31:0] src58;
    reg [31:0] src59;
    reg [31:0] src60;
    reg [31:0] src61;
    reg [31:0] src62;
    reg [31:0] src63;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [0:0] dst35;
    wire [0:0] dst36;
    wire [0:0] dst37;
    wire [0:0] dst38;
    wire [0:0] dst39;
    wire [0:0] dst40;
    wire [0:0] dst41;
    wire [0:0] dst42;
    wire [0:0] dst43;
    wire [0:0] dst44;
    wire [0:0] dst45;
    wire [0:0] dst46;
    wire [0:0] dst47;
    wire [0:0] dst48;
    wire [0:0] dst49;
    wire [0:0] dst50;
    wire [0:0] dst51;
    wire [0:0] dst52;
    wire [0:0] dst53;
    wire [0:0] dst54;
    wire [0:0] dst55;
    wire [0:0] dst56;
    wire [0:0] dst57;
    wire [0:0] dst58;
    wire [0:0] dst59;
    wire [0:0] dst60;
    wire [0:0] dst61;
    wire [0:0] dst62;
    wire [0:0] dst63;
    wire [0:0] dst64;
    wire [0:0] dst65;
    wire [0:0] dst66;
    wire [0:0] dst67;
    wire [0:0] dst68;
    wire [68:0] srcsum;
    wire [68:0] dstsum;
    wire test;
    compressor_CLA32_64 compressor_CLA32_64(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .src30(src30),
        .src31(src31),
        .src32(src32),
        .src33(src33),
        .src34(src34),
        .src35(src35),
        .src36(src36),
        .src37(src37),
        .src38(src38),
        .src39(src39),
        .src40(src40),
        .src41(src41),
        .src42(src42),
        .src43(src43),
        .src44(src44),
        .src45(src45),
        .src46(src46),
        .src47(src47),
        .src48(src48),
        .src49(src49),
        .src50(src50),
        .src51(src51),
        .src52(src52),
        .src53(src53),
        .src54(src54),
        .src55(src55),
        .src56(src56),
        .src57(src57),
        .src58(src58),
        .src59(src59),
        .src60(src60),
        .src61(src61),
        .src62(src62),
        .src63(src63),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34),
        .dst35(dst35),
        .dst36(dst36),
        .dst37(dst37),
        .dst38(dst38),
        .dst39(dst39),
        .dst40(dst40),
        .dst41(dst41),
        .dst42(dst42),
        .dst43(dst43),
        .dst44(dst44),
        .dst45(dst45),
        .dst46(dst46),
        .dst47(dst47),
        .dst48(dst48),
        .dst49(dst49),
        .dst50(dst50),
        .dst51(dst51),
        .dst52(dst52),
        .dst53(dst53),
        .dst54(dst54),
        .dst55(dst55),
        .dst56(dst56),
        .dst57(dst57),
        .dst58(dst58),
        .dst59(dst59),
        .dst60(dst60),
        .dst61(dst61),
        .dst62(dst62),
        .dst63(dst63),
        .dst64(dst64),
        .dst65(dst65),
        .dst66(dst66),
        .dst67(dst67),
        .dst68(dst68));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29] + src0[30] + src0[31])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29] + src1[30] + src1[31])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29] + src2[30] + src2[31])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29] + src3[30] + src3[31])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29] + src4[30] + src4[31])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29] + src5[30] + src5[31])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29] + src6[30] + src6[31])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29] + src7[30] + src7[31])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29] + src8[30] + src8[31])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29] + src9[30] + src9[31])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29] + src10[30] + src10[31])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29] + src11[30] + src11[31])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29] + src12[30] + src12[31])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29] + src13[30] + src13[31])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29] + src14[30] + src14[31])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29] + src15[30] + src15[31])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29] + src16[30] + src16[31])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29] + src17[30] + src17[31])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29] + src18[30] + src18[31])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29] + src19[30] + src19[31])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29] + src20[30] + src20[31])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29] + src21[30] + src21[31])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29] + src22[30] + src22[31])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29] + src23[30] + src23[31])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29] + src24[30] + src24[31])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29] + src25[30] + src25[31])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29] + src26[30] + src26[31])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29] + src27[30] + src27[31])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29] + src28[30] + src28[31])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29] + src29[30] + src29[31])<<29) + ((src30[0] + src30[1] + src30[2] + src30[3] + src30[4] + src30[5] + src30[6] + src30[7] + src30[8] + src30[9] + src30[10] + src30[11] + src30[12] + src30[13] + src30[14] + src30[15] + src30[16] + src30[17] + src30[18] + src30[19] + src30[20] + src30[21] + src30[22] + src30[23] + src30[24] + src30[25] + src30[26] + src30[27] + src30[28] + src30[29] + src30[30] + src30[31])<<30) + ((src31[0] + src31[1] + src31[2] + src31[3] + src31[4] + src31[5] + src31[6] + src31[7] + src31[8] + src31[9] + src31[10] + src31[11] + src31[12] + src31[13] + src31[14] + src31[15] + src31[16] + src31[17] + src31[18] + src31[19] + src31[20] + src31[21] + src31[22] + src31[23] + src31[24] + src31[25] + src31[26] + src31[27] + src31[28] + src31[29] + src31[30] + src31[31])<<31) + ((src32[0] + src32[1] + src32[2] + src32[3] + src32[4] + src32[5] + src32[6] + src32[7] + src32[8] + src32[9] + src32[10] + src32[11] + src32[12] + src32[13] + src32[14] + src32[15] + src32[16] + src32[17] + src32[18] + src32[19] + src32[20] + src32[21] + src32[22] + src32[23] + src32[24] + src32[25] + src32[26] + src32[27] + src32[28] + src32[29] + src32[30] + src32[31])<<32) + ((src33[0] + src33[1] + src33[2] + src33[3] + src33[4] + src33[5] + src33[6] + src33[7] + src33[8] + src33[9] + src33[10] + src33[11] + src33[12] + src33[13] + src33[14] + src33[15] + src33[16] + src33[17] + src33[18] + src33[19] + src33[20] + src33[21] + src33[22] + src33[23] + src33[24] + src33[25] + src33[26] + src33[27] + src33[28] + src33[29] + src33[30] + src33[31])<<33) + ((src34[0] + src34[1] + src34[2] + src34[3] + src34[4] + src34[5] + src34[6] + src34[7] + src34[8] + src34[9] + src34[10] + src34[11] + src34[12] + src34[13] + src34[14] + src34[15] + src34[16] + src34[17] + src34[18] + src34[19] + src34[20] + src34[21] + src34[22] + src34[23] + src34[24] + src34[25] + src34[26] + src34[27] + src34[28] + src34[29] + src34[30] + src34[31])<<34) + ((src35[0] + src35[1] + src35[2] + src35[3] + src35[4] + src35[5] + src35[6] + src35[7] + src35[8] + src35[9] + src35[10] + src35[11] + src35[12] + src35[13] + src35[14] + src35[15] + src35[16] + src35[17] + src35[18] + src35[19] + src35[20] + src35[21] + src35[22] + src35[23] + src35[24] + src35[25] + src35[26] + src35[27] + src35[28] + src35[29] + src35[30] + src35[31])<<35) + ((src36[0] + src36[1] + src36[2] + src36[3] + src36[4] + src36[5] + src36[6] + src36[7] + src36[8] + src36[9] + src36[10] + src36[11] + src36[12] + src36[13] + src36[14] + src36[15] + src36[16] + src36[17] + src36[18] + src36[19] + src36[20] + src36[21] + src36[22] + src36[23] + src36[24] + src36[25] + src36[26] + src36[27] + src36[28] + src36[29] + src36[30] + src36[31])<<36) + ((src37[0] + src37[1] + src37[2] + src37[3] + src37[4] + src37[5] + src37[6] + src37[7] + src37[8] + src37[9] + src37[10] + src37[11] + src37[12] + src37[13] + src37[14] + src37[15] + src37[16] + src37[17] + src37[18] + src37[19] + src37[20] + src37[21] + src37[22] + src37[23] + src37[24] + src37[25] + src37[26] + src37[27] + src37[28] + src37[29] + src37[30] + src37[31])<<37) + ((src38[0] + src38[1] + src38[2] + src38[3] + src38[4] + src38[5] + src38[6] + src38[7] + src38[8] + src38[9] + src38[10] + src38[11] + src38[12] + src38[13] + src38[14] + src38[15] + src38[16] + src38[17] + src38[18] + src38[19] + src38[20] + src38[21] + src38[22] + src38[23] + src38[24] + src38[25] + src38[26] + src38[27] + src38[28] + src38[29] + src38[30] + src38[31])<<38) + ((src39[0] + src39[1] + src39[2] + src39[3] + src39[4] + src39[5] + src39[6] + src39[7] + src39[8] + src39[9] + src39[10] + src39[11] + src39[12] + src39[13] + src39[14] + src39[15] + src39[16] + src39[17] + src39[18] + src39[19] + src39[20] + src39[21] + src39[22] + src39[23] + src39[24] + src39[25] + src39[26] + src39[27] + src39[28] + src39[29] + src39[30] + src39[31])<<39) + ((src40[0] + src40[1] + src40[2] + src40[3] + src40[4] + src40[5] + src40[6] + src40[7] + src40[8] + src40[9] + src40[10] + src40[11] + src40[12] + src40[13] + src40[14] + src40[15] + src40[16] + src40[17] + src40[18] + src40[19] + src40[20] + src40[21] + src40[22] + src40[23] + src40[24] + src40[25] + src40[26] + src40[27] + src40[28] + src40[29] + src40[30] + src40[31])<<40) + ((src41[0] + src41[1] + src41[2] + src41[3] + src41[4] + src41[5] + src41[6] + src41[7] + src41[8] + src41[9] + src41[10] + src41[11] + src41[12] + src41[13] + src41[14] + src41[15] + src41[16] + src41[17] + src41[18] + src41[19] + src41[20] + src41[21] + src41[22] + src41[23] + src41[24] + src41[25] + src41[26] + src41[27] + src41[28] + src41[29] + src41[30] + src41[31])<<41) + ((src42[0] + src42[1] + src42[2] + src42[3] + src42[4] + src42[5] + src42[6] + src42[7] + src42[8] + src42[9] + src42[10] + src42[11] + src42[12] + src42[13] + src42[14] + src42[15] + src42[16] + src42[17] + src42[18] + src42[19] + src42[20] + src42[21] + src42[22] + src42[23] + src42[24] + src42[25] + src42[26] + src42[27] + src42[28] + src42[29] + src42[30] + src42[31])<<42) + ((src43[0] + src43[1] + src43[2] + src43[3] + src43[4] + src43[5] + src43[6] + src43[7] + src43[8] + src43[9] + src43[10] + src43[11] + src43[12] + src43[13] + src43[14] + src43[15] + src43[16] + src43[17] + src43[18] + src43[19] + src43[20] + src43[21] + src43[22] + src43[23] + src43[24] + src43[25] + src43[26] + src43[27] + src43[28] + src43[29] + src43[30] + src43[31])<<43) + ((src44[0] + src44[1] + src44[2] + src44[3] + src44[4] + src44[5] + src44[6] + src44[7] + src44[8] + src44[9] + src44[10] + src44[11] + src44[12] + src44[13] + src44[14] + src44[15] + src44[16] + src44[17] + src44[18] + src44[19] + src44[20] + src44[21] + src44[22] + src44[23] + src44[24] + src44[25] + src44[26] + src44[27] + src44[28] + src44[29] + src44[30] + src44[31])<<44) + ((src45[0] + src45[1] + src45[2] + src45[3] + src45[4] + src45[5] + src45[6] + src45[7] + src45[8] + src45[9] + src45[10] + src45[11] + src45[12] + src45[13] + src45[14] + src45[15] + src45[16] + src45[17] + src45[18] + src45[19] + src45[20] + src45[21] + src45[22] + src45[23] + src45[24] + src45[25] + src45[26] + src45[27] + src45[28] + src45[29] + src45[30] + src45[31])<<45) + ((src46[0] + src46[1] + src46[2] + src46[3] + src46[4] + src46[5] + src46[6] + src46[7] + src46[8] + src46[9] + src46[10] + src46[11] + src46[12] + src46[13] + src46[14] + src46[15] + src46[16] + src46[17] + src46[18] + src46[19] + src46[20] + src46[21] + src46[22] + src46[23] + src46[24] + src46[25] + src46[26] + src46[27] + src46[28] + src46[29] + src46[30] + src46[31])<<46) + ((src47[0] + src47[1] + src47[2] + src47[3] + src47[4] + src47[5] + src47[6] + src47[7] + src47[8] + src47[9] + src47[10] + src47[11] + src47[12] + src47[13] + src47[14] + src47[15] + src47[16] + src47[17] + src47[18] + src47[19] + src47[20] + src47[21] + src47[22] + src47[23] + src47[24] + src47[25] + src47[26] + src47[27] + src47[28] + src47[29] + src47[30] + src47[31])<<47) + ((src48[0] + src48[1] + src48[2] + src48[3] + src48[4] + src48[5] + src48[6] + src48[7] + src48[8] + src48[9] + src48[10] + src48[11] + src48[12] + src48[13] + src48[14] + src48[15] + src48[16] + src48[17] + src48[18] + src48[19] + src48[20] + src48[21] + src48[22] + src48[23] + src48[24] + src48[25] + src48[26] + src48[27] + src48[28] + src48[29] + src48[30] + src48[31])<<48) + ((src49[0] + src49[1] + src49[2] + src49[3] + src49[4] + src49[5] + src49[6] + src49[7] + src49[8] + src49[9] + src49[10] + src49[11] + src49[12] + src49[13] + src49[14] + src49[15] + src49[16] + src49[17] + src49[18] + src49[19] + src49[20] + src49[21] + src49[22] + src49[23] + src49[24] + src49[25] + src49[26] + src49[27] + src49[28] + src49[29] + src49[30] + src49[31])<<49) + ((src50[0] + src50[1] + src50[2] + src50[3] + src50[4] + src50[5] + src50[6] + src50[7] + src50[8] + src50[9] + src50[10] + src50[11] + src50[12] + src50[13] + src50[14] + src50[15] + src50[16] + src50[17] + src50[18] + src50[19] + src50[20] + src50[21] + src50[22] + src50[23] + src50[24] + src50[25] + src50[26] + src50[27] + src50[28] + src50[29] + src50[30] + src50[31])<<50) + ((src51[0] + src51[1] + src51[2] + src51[3] + src51[4] + src51[5] + src51[6] + src51[7] + src51[8] + src51[9] + src51[10] + src51[11] + src51[12] + src51[13] + src51[14] + src51[15] + src51[16] + src51[17] + src51[18] + src51[19] + src51[20] + src51[21] + src51[22] + src51[23] + src51[24] + src51[25] + src51[26] + src51[27] + src51[28] + src51[29] + src51[30] + src51[31])<<51) + ((src52[0] + src52[1] + src52[2] + src52[3] + src52[4] + src52[5] + src52[6] + src52[7] + src52[8] + src52[9] + src52[10] + src52[11] + src52[12] + src52[13] + src52[14] + src52[15] + src52[16] + src52[17] + src52[18] + src52[19] + src52[20] + src52[21] + src52[22] + src52[23] + src52[24] + src52[25] + src52[26] + src52[27] + src52[28] + src52[29] + src52[30] + src52[31])<<52) + ((src53[0] + src53[1] + src53[2] + src53[3] + src53[4] + src53[5] + src53[6] + src53[7] + src53[8] + src53[9] + src53[10] + src53[11] + src53[12] + src53[13] + src53[14] + src53[15] + src53[16] + src53[17] + src53[18] + src53[19] + src53[20] + src53[21] + src53[22] + src53[23] + src53[24] + src53[25] + src53[26] + src53[27] + src53[28] + src53[29] + src53[30] + src53[31])<<53) + ((src54[0] + src54[1] + src54[2] + src54[3] + src54[4] + src54[5] + src54[6] + src54[7] + src54[8] + src54[9] + src54[10] + src54[11] + src54[12] + src54[13] + src54[14] + src54[15] + src54[16] + src54[17] + src54[18] + src54[19] + src54[20] + src54[21] + src54[22] + src54[23] + src54[24] + src54[25] + src54[26] + src54[27] + src54[28] + src54[29] + src54[30] + src54[31])<<54) + ((src55[0] + src55[1] + src55[2] + src55[3] + src55[4] + src55[5] + src55[6] + src55[7] + src55[8] + src55[9] + src55[10] + src55[11] + src55[12] + src55[13] + src55[14] + src55[15] + src55[16] + src55[17] + src55[18] + src55[19] + src55[20] + src55[21] + src55[22] + src55[23] + src55[24] + src55[25] + src55[26] + src55[27] + src55[28] + src55[29] + src55[30] + src55[31])<<55) + ((src56[0] + src56[1] + src56[2] + src56[3] + src56[4] + src56[5] + src56[6] + src56[7] + src56[8] + src56[9] + src56[10] + src56[11] + src56[12] + src56[13] + src56[14] + src56[15] + src56[16] + src56[17] + src56[18] + src56[19] + src56[20] + src56[21] + src56[22] + src56[23] + src56[24] + src56[25] + src56[26] + src56[27] + src56[28] + src56[29] + src56[30] + src56[31])<<56) + ((src57[0] + src57[1] + src57[2] + src57[3] + src57[4] + src57[5] + src57[6] + src57[7] + src57[8] + src57[9] + src57[10] + src57[11] + src57[12] + src57[13] + src57[14] + src57[15] + src57[16] + src57[17] + src57[18] + src57[19] + src57[20] + src57[21] + src57[22] + src57[23] + src57[24] + src57[25] + src57[26] + src57[27] + src57[28] + src57[29] + src57[30] + src57[31])<<57) + ((src58[0] + src58[1] + src58[2] + src58[3] + src58[4] + src58[5] + src58[6] + src58[7] + src58[8] + src58[9] + src58[10] + src58[11] + src58[12] + src58[13] + src58[14] + src58[15] + src58[16] + src58[17] + src58[18] + src58[19] + src58[20] + src58[21] + src58[22] + src58[23] + src58[24] + src58[25] + src58[26] + src58[27] + src58[28] + src58[29] + src58[30] + src58[31])<<58) + ((src59[0] + src59[1] + src59[2] + src59[3] + src59[4] + src59[5] + src59[6] + src59[7] + src59[8] + src59[9] + src59[10] + src59[11] + src59[12] + src59[13] + src59[14] + src59[15] + src59[16] + src59[17] + src59[18] + src59[19] + src59[20] + src59[21] + src59[22] + src59[23] + src59[24] + src59[25] + src59[26] + src59[27] + src59[28] + src59[29] + src59[30] + src59[31])<<59) + ((src60[0] + src60[1] + src60[2] + src60[3] + src60[4] + src60[5] + src60[6] + src60[7] + src60[8] + src60[9] + src60[10] + src60[11] + src60[12] + src60[13] + src60[14] + src60[15] + src60[16] + src60[17] + src60[18] + src60[19] + src60[20] + src60[21] + src60[22] + src60[23] + src60[24] + src60[25] + src60[26] + src60[27] + src60[28] + src60[29] + src60[30] + src60[31])<<60) + ((src61[0] + src61[1] + src61[2] + src61[3] + src61[4] + src61[5] + src61[6] + src61[7] + src61[8] + src61[9] + src61[10] + src61[11] + src61[12] + src61[13] + src61[14] + src61[15] + src61[16] + src61[17] + src61[18] + src61[19] + src61[20] + src61[21] + src61[22] + src61[23] + src61[24] + src61[25] + src61[26] + src61[27] + src61[28] + src61[29] + src61[30] + src61[31])<<61) + ((src62[0] + src62[1] + src62[2] + src62[3] + src62[4] + src62[5] + src62[6] + src62[7] + src62[8] + src62[9] + src62[10] + src62[11] + src62[12] + src62[13] + src62[14] + src62[15] + src62[16] + src62[17] + src62[18] + src62[19] + src62[20] + src62[21] + src62[22] + src62[23] + src62[24] + src62[25] + src62[26] + src62[27] + src62[28] + src62[29] + src62[30] + src62[31])<<62) + ((src63[0] + src63[1] + src63[2] + src63[3] + src63[4] + src63[5] + src63[6] + src63[7] + src63[8] + src63[9] + src63[10] + src63[11] + src63[12] + src63[13] + src63[14] + src63[15] + src63[16] + src63[17] + src63[18] + src63[19] + src63[20] + src63[21] + src63[22] + src63[23] + src63[24] + src63[25] + src63[26] + src63[27] + src63[28] + src63[29] + src63[30] + src63[31])<<63);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34) + ((dst35[0])<<35) + ((dst36[0])<<36) + ((dst37[0])<<37) + ((dst38[0])<<38) + ((dst39[0])<<39) + ((dst40[0])<<40) + ((dst41[0])<<41) + ((dst42[0])<<42) + ((dst43[0])<<43) + ((dst44[0])<<44) + ((dst45[0])<<45) + ((dst46[0])<<46) + ((dst47[0])<<47) + ((dst48[0])<<48) + ((dst49[0])<<49) + ((dst50[0])<<50) + ((dst51[0])<<51) + ((dst52[0])<<52) + ((dst53[0])<<53) + ((dst54[0])<<54) + ((dst55[0])<<55) + ((dst56[0])<<56) + ((dst57[0])<<57) + ((dst58[0])<<58) + ((dst59[0])<<59) + ((dst60[0])<<60) + ((dst61[0])<<61) + ((dst62[0])<<62) + ((dst63[0])<<63) + ((dst64[0])<<64) + ((dst65[0])<<65) + ((dst66[0])<<66) + ((dst67[0])<<67) + ((dst68[0])<<68);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha5f8d4bafea22cc957469750eade12012b4a2e7628a0f5dc1c5a856586ae1cc6075f39d1b96e47295b753ec935deea9601a6e5b4f435dc1e3813bdc1f222c146b3cd293b3132192821cdeccd0d7feee259476a81f221e5cfac69c144dd01254cafafa5664d701134912717c3a43393917868f83670af9c1c0d2b614f44c02b96bb6e49d8f7704a4e515a14cccfe8663b1839dcf42ee6d1087ded0e6a9a3f8161e9f5b44235e8d13198fb09405117099ed483539237c5ae38983f9db851244cc2fd3074a55c73bdfad6b1d6cea7911f553ce1483d801a79f70c2bfe53a62ca5fbd0cf9d8e1b09874a1a898b309af2d523b366918cf191d1d9186cacd369c6c4a2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h571b8953d021249400828d86dbfbe51c1b1cc9fda97bcb1be2e69cf6e76c80f32dec190fe532b1a09e213e7760c7fa84a67eec7b9b7d23ea49a6d2b70a796b8537127796f0517b32c4e0b07f626f61a8f6dd99afe828a40d96cc7a9688a3e1417846aad2e709535d73191c3f21218d8dab708551b522b5228af943e32bf9238a83ad2221bb82f04df1c93ffd5285e524bab6d57b267336fff12477b73bc4ff2491d420e192357efb124368ff7b54f681c420dbb66003ebc52b649a127402a8d0803c6a2359525b14904d5df344e3de84dd486032d1e97ad8dd1bd48b33ba1d25d8beab0d2bd4424d0a0a36c3a5947575c9db11462b3e9e6a8e4c424094912b99;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h515fc4be9e988ba3b54837ded8116098046e0f8c3465d72a46c6fca70c8f1e7f7947f3d9b12bb3460db6cc7f6084e744b4b8a63a68bb4b7d8f8f9a9219e3c3cb853aaa7b68a7bb2f5a5e8360bfc30ea81ceb2bbf10573b28a3d1af03ece377ac6709d60d593dbb5a784dc7ed02fe57948f2e75b226eaa6864ab36f9610e7310782d826ccd97ea474334b5d8bc6d65a61eb9c7a82dab42b320d4aab693f27f541b67f57d9868edf0b93ff9008b4499f83fa38d934f1ddf90306e6e955e07b1ed46baf7255354f1cdae64fbf4d64a9e491f87b2adac3f2b8ecd2e6503693999c592fa3a63d6a8f96cf6cc220c26fa495f2265191142cdd5f9e0968fb1362729c4f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h98f6e600017c927d4b74f7db9747319d1c62a7b4f6792b6221f35aa67c1f3b4a64e8d5f609a86be861f44342596e6ee33b57f6ba48044dabf0dc567c44639e43c1e93dcc23a79cc30271571d5c50a9c35e088dc3b9deb4c2406377bf2a709ca209a6c78d18b48ac291940652cf10e9a1efe70b181c0ec7089752cdf1e30575ce13384a7d8d04ddde502fc9c5b3894928cb299e5d94139151ad2c16e5d3efc09cb9075e91dcac4aa49e54955719c90b9403e3548867f2cc538f9f6156fa442ce2cf161c87ba3f61005172efec265f5f266d6426ad6e94484038a820d5edc5038bd76dcb992acb86102d4c1a37ecb3af94476e48fe231dbeb4ab51c10702767e8c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h439a04e96fb2c4f9601d540d747e8031da729d991fded85f0d383228436d51879b90c9de70bc37f49c4469e424e3de6b26578b4384c5280adbe44177ae158d30e3d872a3d09526d1037a4cc64b4dc33033b89e84afc3b62f89a48524476e446ec97a63c6f78f9122ad2da1103d006b88d30ac7e9b16cf38b0fa085d1702e34da31b6e0093f546e586f8eae746d0482cf72f5baea52fa9c4b2f8a5d1f42d133d585099d6eb4d3813f4070f2961ce3fc0ef5e82022c3c68136a38f9b8b1fe2b7d9f282fca0221e2e3c70b87f71a7c3e88374c6de432705a59f90d9443c1edbf078cd93540628afcef6669a18dc6521b59547a02306d132713915f3ea69d8fa0e6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h40b167aedb43eb31f42e126cdfbd10b5aa0e3622ef1155529898732e45c89b919c72350379e6b47676a7654a7161a84068f11ec74f141a33f43509d281832cd7549edb82084b091509a4ee27101c5fb01a5243007bd40e0f12be54818581b1775a9f8d7aea50f8b3297ab84a29f5d5981189f543ae2b4ae17ae2b9c25af5af99f0087a37d77b9c55009828a788535f936b6162bd6adb2558e3d651ad61c703172c9fbced937d62681632768b910d4afefebc7ed96f17bc7ffaf12eff58d66c227f2d8228d8a8c2f803bc55368b86a1a626a929611fff525dec7ca2bc915b378f4b8ea7591972b5ad77d1e67fa21fdbc272db269350cfbe22fdb286d4982279f3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h65fd0735411b412e0f4f0c1865810115de14155e11465a95498123e77757ae110dfa39582777b4cb79a0943094363d107e274f46037ef8f280da968c5bd7367a323931cbf89592d2b39eaa66b5dd732559abc98827bca30c888ab350d345641a074b0508b98ac2c4f8504fd382e760d3172e52958f9cac48e97a0e7de5a5e34344a2b7a4ecfea759e3012615e6707c8d330f77da2be9dd80aa75042979b75ba1288dd2c1a6dd8867a8e1c80ff78fec23bc6aab91ccea7e3f3b975acc2b04aa1d75275ba4e266c9e9d0761f484acd8ad36e6f41c6916378c29c1c3831e341a59cc51f30def8472cc54d99836c2a95ef2bba2627699b9aa9d2cc7067a7860d10d3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he7af09773b5f9de2761a8c8e309650d0dd2d7987a4bfe01cf1e638734cd70882c259ad3576484e70eec9bc0742f38b03a358fe047801498d9222f555ea8e13b0f3eea1898c8809133b2d98809f903f43982c1a03fec737e3e8a318e741ca7a113cb9be72c34dff99c997cfaf27ad7ee886743841d63c9cf66c124b645b46f4811c7abd8865330d2913d7cd808542cf44b7bf77c321e610ae387049d9b22e6271fb6b5be30cf391852a03a58b866fa598d18fbf21f2f00924ec7a37f82de83ce0f4e45f4d03645de7492555f388d8519091781a2fb8f2f794174d868beb057c69ad653ab27eee41888cab28b74843c4a88e304f363093e84bec70e3f5837e8fce;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7597d0a40f25d45f306f9c4f7cf85b647fc52c3cfee60d54498236d40a91ba00bf18e7e7ae858ce117dd38944614a6c8f82f71d8cef474740260bacd37934acc4440ac9288670a9322e9a0a1a6f8618082409a1a67a8f3572cee18f8456865424b93a22609cc924112a195ec44e3e2fd0a471969549308443bc28d1e05a6acf3e44aa69e2869275b124c5b1cb0f9607827284a7010a6d0b251274c7f0865e65d4759ab322a8b907ce1c5fe371c8aa5a0cd84ba7f805ab2abd58cdcab410c31fb16fc02a7350b7b75e3d4c201d0d6d1daf574d0c5665d82438003c9b6a9067906fa9774f066533a1ab5abc39a18efbd087ca03e97610793f3a4c7333d3b2af6d2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h595976d4d6f51d7349bb6900e13ea3441df57f21aa8bd66e92538a074d07f29067c0cd8728c76f9fb762d67ab802f7de80005a523ae50a7a97dd702a8203a000223a286fdc92d85380a20fdc68c85fc6e39c7df6e40a0c3ad1dd0a24c3e4d42503e3af481c7e0eac1036572ec472ae8dd7f753b5a1da8b7ea78bef5f8b67d582b5b09a576abab7df795efb4de0fa2b195f281f7eb00ff7d9eb3136ea9339307ac9bf6e8d43e25df7d41000c213d5bd5293c87dd82ec7e3aa136e19fd7414b1b8f6ee54b2d3b186c4b44a94f52ee8534a76168fdce32ced51c46c6d3b20677faf27b2f603462c28cc038c08ee39ea0d6092effc7e07a08753560fabd66e5e4d35;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd95f542e9e7d6d543e20a974f60cc05ade3fc040514f1aed4440483342f77bd1ac1408fd509ece54541025dec6a69ac20fcb888705e82fcf643595feef57fd0ed9d9e80694d89a2bb46cbfe3673b98896585c0c2ca97d74d2abc885005b975ce13e1e12fdf96664e5734fb42657777baaa5aaf8ad206571632270926a1a430d6313cb0adf1c587afa72b5bd061b7f27842e5a602693d5c141fb93a2d3bda71ebfa6baaa5581fa2df1661999928c1594d5f06283a6ab36de83d44c14fe950829f479d5617ae646b35e53f46dae4de5a922d6f582066d9d4000d17069c6ebb52330747d243051552a8ab850cb792cd52f3cbf3d704f88913548d049fa5596409fd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha57e581309c378114578d311186388f44cd917b8d053cec6a6efbdad1575d4c5ce5f8f699115947afb599b42a07f8bb3441ff61496a3b571ddac5e59e2f341a0e7d0ad38e881e589f51df51f63cefe323792c2efc24590e3c250a3ac4ff56ee52be889e32a82ee6115805401ddc60953e349fd8dcbc3a54be2ca9340d146a8de9235252766a037b334a583866934f15be53fa5c88d21b61d2fdd3af8817d6648375358f843e24e45256b73d47c8db85c7469bc8a9ef999001c3374c2f127fb4dbd824a4a7e15b4a27fbf040eff673201cb68f24b91ad7f527506845e47b6070c8ff4989e2ba19fa6c4a68761ae7284f1d1f105129654931a711cc1d8d77a08f4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8b3121f292ad7553b9d764106cc17156a2b613a336a4248acbe0d3db43fdab8295b44198fc3cb1ab02caf1ae60437480adccf642dd36fd243892b03385d5c4b1b7795fe825f6038af4eba8a293706ea1d1bc6508ccd28625a35ba50e9ca81c96db8a9599ed565bb75edf154ac5302f0b63e959d8e62c1c79a16772ce7cd196f6462f955312e338a448b0c7b32e8dddec583642f4c5e70d0e382ce7761a1f3a6daeaa59ac2b5129084eb4007746cca1092c975c0f58f3771d11f81ae03355707e87457139a24d7869b25d9011c37c695e6a784f3178594d3a4d4537641c1df37231153c6b84a60acda2d7e111ef6638112cd7d835f340e76c72dd8b7c9d868b1f;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4c9926c8a24e37c2b8b80da46c832cdbda04d2f510cd6dde4c7eca5722a514c4e0acc43d8bedcd33d9f11ce70cab073332b6faf3445e8c4c66fc1e5bd23f61874e8adcdb7b80dfce22aa87bc9a82f20b853105e237eb56766ebc8a8e7338e029d75071ade1aa26c12ca2c7f584243b1a9bf6759f70ca548fbaa448fc8eba255b8466b901d22a3387d9debcebec2e1a32a7e659911ba5a628aaa978923ce17df88faad8c43b5f9da5e8468e21ed59ebae21662ed6ff3b56f8d10a5736d17e2a934891819df9de6e4c24fb0224fe3b4b3393fa36eb7661e9c87e209f97149606ae8c4ee5bb31d1a3d77f618f81e8dce8af92f3bcd509969a5a1d80490244263002;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h85bf21b79d27d11b55774a92134ce0150e843b8b595595da8ecdbb669e3d96bc12a248ca4f3a889ba5d33a5003a7fae746c9d1e6b9b994348cefb43de97a58409089f88e7c5f3a4f02d989591887c8a83a66b75d4298025054267183ebdc86531256ffb7cbef147174f7b8dcda1074dd4665f95ea10f8102c8e5511e8fcbabd763d7842b0dded3c053bae1be405a0d88824391a13e52f482066a31d6602105cbed70c7c9def079ae133abf630377f9f1fbe558125c2aa0c1d37fa14cc6cf1c259a5c95cff756314392016919a21bd38f3fa10d8cd6f8f0c18f6d9d42b2a7d71cc97acd2fcbd27f914809fd8d55ecf59253db2049892d802de0807d8199c455bc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9f68db272e681f42395066b84fd2a6ce8c941560749ffe6fcd05a0480f515b00ed752ea7522d59f3cb3963d4c9af75a1f596d08686cb4efe79fb724592fdbb1319880485cfad1f888dd99ad3962820cc1e5cf62de6021140bc4f7c76b7c6840ea430309f6bc612044cf116f9579feba84bcfa1f3fc23fcb697e167248d1b1f3b0f4148aad3d590cc1463f128b12500640648e762360eb226179f9f83930a72442c9baa44992155f37e97b8edeb590ff3c666bfa29aeb04875e5dd3dbca0d4d655ba3515818e562a18d24bdad15db7617c82b2237664b009730e3054cfd14844bb009e45325036dbc7607406aee828104d4645b7f9e03a13f5ec1a698189dbfb6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h43d79de6482beaf1977cd29de219f7d8d3fbf40c7237858947b00c6e11e3a753dffdb04474dcc817d45d5abeca6930aeef9c601305fb9c18554a1189d0262fe65b8a5a76fedd360d01496c0f75622031398cf3ef65095d9f17c09f9051aafc23861e5ede65c6e737bf20960affcf5266839fa1fdb9bf373e460fabc79602fc6a9adf498eb39663fff73d9f76ba24d55261890dda7b330dbbe0e7bc28d15fd48cb1d60f0181151aa0e12bb725050c602c2cf88517035327b10bcdc2c930dfcbd4a344d0c32c72215b3bf8cf467afa23248f02773730f3df1b8bb74f3642b61b7dcc7ffcfc775f0c841d4bfbb10f5ca932208a152578d62bba24310a99eec34d4b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfd78f7733fab2f1703652f0e9b51ebf053b765b8e4c15235807e7a0bd45ed896ca64ee29940cbba46df204c8902e7d85a7bd37492c04ea20dcb004172b714b8deb862417607f14f8bde103304c2fc47c5837ba81796f88b2e2d904237eeed1eb0f15390fea5be3097738af5fc4a5aebd8fa86627b9e40b23ce6b1153e76370696ee073d9fe429d6eb24d37522031cc5e8448a4b12883ff9a4bb59694c074f034bceceeaab87a1a63058f099a03567e85bd4b59f9956115d83e89f5685a50c5ab44ed2d707a630f5949f6f96ff597ba958eb419440b3be0fbc7d72e2a9a81b31a0630b99d69e7a6cb74b5372e38edfc6685d36265bca2c80ee88968aec0ec2bb6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h5e97dd80bbc6e88bb48c6ec424f8b295f099aacf1493c22fc2227357af8ae76befce743dda86e76bf66f3768fd275afbca4b7db635fb9d05d0a5d859f544c1d365be51fbd2d15ff6695f90bb895080df6986b2fa52918acf60eb54dc45827b6fe7721cc7070bb59d59fcfa096b897c183b6f1269902158bcd1029b66aac4d5049d97a80114f0e190c036516276b75a7b61d7c31dd8dbe8b4e1879c28815264ccfa603b387ccb700365c6d7eb6647295993bb7b9fa87f693039ebac0114fbed3f8c28826e5a2c73c979ce42ce3d7f4ece3363016f0101b88dcfc925d1d3745ae049330083a07c9907c66358450ded259b466174d90ec29fbf8d93ef74f54e49b3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h86204dda68865329d72f04809173c161d624eb7a483acda14d39eda838e85ecbaa7e26ef2bb6a6d08130b9412f7948b1bb5d79345d7becaafd2ff615aa7b6e90fe48ee13497ca30b615a5fa8206165d8701a7524ad18e0267c10726d52d9d1768c89cc3ce5d8bcbe0351e37fd347f0b2d4fdd88f21194b6cad2cbefa78d36a83aedb7feac85283a3946a6a9743c249706a72876fb56d7c248f69c9db0e1670a8f2a570a605bafc27a95b15f24dbe673a84d00a1725b185da8d6adca9b23446c8c1ef321b3573b451be8d94e327e57bd8adc2c4c55bdd4d1c674d74c7c97c0c473b70cf8bf2de90cd7c3eff732cb5fae34fd4c9ef547821039bab962eabfb65c7;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he1c077b12c69f7f8287cd024a18c0439c86e934cd435901c52148846afd61f012caddc1e76192e4e3e3651385f18db5c444dcb5b5a14a1fd32fbd3d45d8cf685fe36066622580c9fcf86412ab3bc76c065eb931c8808f4a4ab58a0eb175ac035d679262312feb23a570343b778f0af982bcfc0699b3ea7989f9dc53540556970929e799cb5a367a156addbbfee1119febe91845dd21e0137afe2fe82ac17e3803014f1e466077a9d5c9080591b618e5d3ed7647d4b42897309938d0333943723a8329c89422fec7d11836e12c569aaa9c87759af03332236cd984abfa9f69d73ad35cbe30de24ce8dcc46c4c817afef0597ec958aaf9826e67d805b7890c807d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb5b47e666115f781eb9920835a9972f9285610a234db6622749ac7939e8f681ece8c6d43c9c47b4224531f6ba18cee29061a6932c1d8ee9d683a204790e2d34684985b4e577f154e864aab9e8d8ae848c3ab5e13c57034ec115650a0528bb22cdb4b4e8da43825f9948a4d68ef26f2a8a7531f1b47d975cec1943b5c1d741214a12c6f36b988a71b2af2180e4c95a05c561f4b41686328277ad059d27ab0ea910c4cdb4dc734edfd69bcc556e78d89a3125a6e5e30dd26330194396034e5df1f6c733dd8df2b466b4e0fc0dc531532dd568766215e38e96b7a07bb797f957b90edc03c8f4fc88618dbce053858c0dca47e82a18466260c8fdd51568a056899a2;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc6e3908dfb648644b903a50162abfaa88a79c22f6433b70d4609ecf909881cad7541fcda5814a44db4688aaa5ef85654f8a2583c5dc1927008e00c86487d406a74c10c90c4c6317850ea7854536eceaa4ff886cf5995a4b2cb91f85f5388fed909f5c10851c2f36e08b37074c7639872628298e81232c9b5ffcb9d78beac4878fa7ff3361fed34b7cc7183ddb0b2006a491b11e95ea65af32495aa18f0925b9f8e28f1d8a401b1a122eb48edee937da2389c6c4cadaa64b0fb41da8b8199eb513b3fcb498b98cbffd87c3b29526ffb100ef040a9912da8c6f62425c84d88d596f219a073c6acb67890ec31c0fcf59077092e4db391d5cdbe88bf1c2ecab59f07;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'habd54d4471e4472272ce4a1811308b2dcb24fcfded5b934ccbeebae21364df2594a938a2e88a2ef950c25f90512ed4078316679b5eacaf09aa5a58ddb03531c538eec9247d51e3585d95a6748834ba60545fb19854b92e22fe6fa41db32abf9cf845adf1ed1c8a8957d7bdc4b2dd9967d878d5c27057d0679f888236ddaef06c7d358038a116150f961c73165cb4571c7d588cd0fb4adbf1b97d1c186f7391936391c06a135a99d266abd1e70c39163bc30bcb9cbc2e11983164610f19ff23f0ef5b7b86125a2bcea9086eb732c3cd503d92aaed2b6948428620d7b2707dcce7a4c27756c67050a883fb387c88fc44e0bbac51ce42c1fb630502991cbefb1712;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h309bf6a24ce026389771ffcd5fce352492a1b1836b35fff390ce54f684648ef545212ee79b41bf7880d669d0b4d50912d1cc7506b83e5014c31f1f87a98df93b4a8b74f595b20362e704ac5082e206f69b76846612e32345b114f6e4a68d55d91df9accaefabbe4901d0f4613ceca0336e10b1534af411effca6a0c098f1ccb574714b57a5ed35c3d746723940e4c06e1ae7af801ff1f93fe1a18faf4a72276a4af7cc78030366c7e33714fe383ac717d4744d088ae011327cc75b22d2d2135e42273ff4fcaaa78b1ae2d54564db183b42677991668aa54ecfb703e9726e611ed8f2e5c85a780e6f882dedb864d9b1524002734f3bbaa68f2b3714c6f59d14ed;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb349db1a40391d57a05cfd76ec355653cd1bf29b48712213ed095eb2cf46aa914f2fe8b5a4b8ff461439c64d6a4481382f0830b22d4a776da1a614a8b63f26274e2aee2a9e21e2c9ed5762b9c42ac4d1530cdfb21ed16cd64b4869a015cefe1c719538bcf944c44d07685b37114b6c89024f1d8b5f6be9d7934930419b7edf5f1995e11080fd719d0a43ff94f981b899bbf09c1ffa846e28dd3866546bf0246ca89d89077bac31542632958c610977ed6ca91793f0940e9aabe2b63597a9d24694fbfd363c843e8bac43a3fdc872d02ed81dbb72171f6d695aacd09ac47963a54b76c4c3008042dfeb7ea2952442d329212d6788ecf3fc5bc1be11d22921f9a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h510fc55f1bd88f32d7413a3fd946977c969146c57c349cdec500cff3f0656239c2b606042493c972c89c497fc85f9761e3b90cc932529448dfc33a526664649bc20e7eedcfba4d1656572ae54a9da620a3c39f05715237b6c684bad63284ac0711c930cabab0d6fcebe83468804185bf869b55b8f0189402fa85a21c34561ab00a6e8f4ab1d663a2de8f3d74be15e2e4a1fd97b81b552501e58baff958647f863ed2d7edf1a62ea2ca5a58482e1fb21f24517c72404a1561b096aa62deeb668f6b09a742270a8de65db116ecf2f1f58b710ef4ffb9767d0a1fda3cfb1fc382bf70e20b175825d4615f09e885d1d44bd70e1e94737d9d9069f4154ee29f4a26d8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h26734823afd5fd2f776b30f779cbefe64661a5a3a641ecedb065b621a666679175c6af364bd12e2b8c6e2fa70c5767a299541dd6bde2a3ac6ef837b651f5e7682f87592034318223d2195d0149124b479caf4c6629c2f9410a1fddab8ce4eab40f0ab2be164e1b657e3a3d250eaedc805adcdc6f58db89209613a6dfdd0fd13bce8354148bf8b6914b4084df2c8b2b648a7416e6cdeb219fe45dc305c4986334c170b1e39684508c25e7cd288bbff4f109be0b90da2efdf68a577ee4a9008a046956af5ede8bde16f2d26b2d29aeed8e5092d158099d7dffb012374e740d54ada921792a6eda69a82a2d2b18e80f8cef8e32e14640594ef257c9f7ddd1e588d0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h767bd01e7151bf3040647d549b8a685c69a65c29b8685ad6a456ec4a21c49a925849cfb15e04121614681688d89701d24e1c5c8cdaf250146437f7f53bfdefae7db500119ffa8b346aa0b85f21b414f346a54c37c1751a37d9b1cc2b1f34b38074c9df211ad104f2f854356ba9ca246364e6bbbe190b69264e420208cda05961efae7f921896b5ced95d44f0db23c33e6e1db530c0fdfc8c7ac8e423f4bfc54590dd52f901d783c2a2c5998f9cda64d5641dac770778fea763594de20ffc85dc3e25038270c1043ed6ed2edf4e570c911a204ae2de92207128f9f65691abe3cf74e60301e6f050b1e7aba48c0de75b8c3faf93f7d0fd7a0d5f101d75daa4bca9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h171dfb734e19b69b723eff6a957654c94d8a92da01ba9e130250cff8c974080ce610decb6ea56e56b501c75d549baa2e9f15bd57f0a191893c5e488d0d67f084fc31148b528ac4baeb86549a0e3688571a5e11a39375b381f8b29b7e9c99376a5813db45b40356b890e0fe6793395c01a083a4fea90c4b66b523138746e48438c2f2a403e3aa81e4eb623730e669531f58dfeb6af42e96658ea95651682b85eaa29a1a348bb54b67d5850ecc16d09b2d3b260a39855ac0c44d3973984f86850e84d2fdc2e9cf16c343ecb7614051f9f7f8896ae579bc665a708c5e24bc05414a2d3bfbc5c132d98c469b273cd652b7bc3419d50e43b318ecf06dd374d3588508;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h366f05ce38135e9ecfcbfefffcf9bd082f06e3854e6e51cd8d572f608bb0fd4d9764fd31b78e6ab1aee16300af88bdc0f20f7d8586dc580e165f49b47917379c026eefa09807815bc14d519e069c37d8cd461961538bb4ffa3e2660709d4f2ebfda02b79653ababcba1ff88bfd273c5169a56d2c20d1f0bdbb820308474f89a12506ff95703e6690b29aa8c874cb711674e4ae2bc472fe1c8319dcd40cdd55755c2c90af29187aa7fbd1fac21e212f8fa8bbbd566da1494b0abba3a2704d62bd2901d52d3c5e9be37fa694b27b13c499fba554f9085a42309eb4e8410a7e4b7def10d659a5b2d11c31358b54591d39db5acf86f8c81d92f1d0b11100c8bccc5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hdb00249a88e6573d2c54e76d0468664f1d40bb586bd16f1561c4686cf46624faad22d488af0f51fb41fbc04ddd9325752abb45d99a8f99407f048f452dc00ec1bf3cbc372c99f0f7ff16d9b263660a18f4e4c0297f86dcbaa19d176b6c798b228e2237898f1ac5e1094e8cbae06b259a17b9d6998eab026a8a9d535415ec345897139cff41835930ca39970c6faa3de01bd54ddd265b5143d9a1be5cf049461bb3750b2529e186212145cb2beb65e0cf565fe6cf74355da9c61a79e773fd0bee64a43d5383712ee7cbf026fea6868d2c43740f0122851455bd786950a55adda01d530a03792f6a1c45eb579d0a16213bf3c1818b78521c790f2be24e2af6c38b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h541e278f82e6ada9323446bb2a1e8780dcb23d073c0ed845933c4d21720af0c16ae620c9016a6394c6f1d2a05c28ba841b1957ed0de97a2d9fe48086edfe1459ecfd3fae7b39686c880c972f56deb10f89492af9e663ed486520d68f2c182c66ea320c6190f19c1f2825b0204734b79b93522135937afb7f0ffe3cd212cb3e515d557666995da28eb06db52bfb07c00a4df7c33e1808dab8ed73894a7079602604e6c5173d56c51b28097ff05d2988622a3c9f7c04b5f72ca608e14a527f60e6572acac962ba2f1651cc668acbd84f5da704a23c085bec837c2ce4c1f5a9ffdeb875507e1fee24876a59d79f73c1284a9fbd0d95568429a0f7cf876564776c7a;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h83d0fde699b9f1da5744d5cefe4bddf10cef2e5ae3ec38aa3b0bffb49e17d1df8775e99562842a80e6e500fecd9ab672d031e2db2c6fc213994e2927f05fe133c8abaeb326299fb898f2460626cc361a5924ca8d9ef4775dc5f171b887d038e1b24734887ae723e144e23539b7998b0819f3c529baf29a589a7d3f82b9c5d93d9b397f49c8999edf357ae14221b9e6c32aeefc74929977d408a93f11ebaee4c6d02fb46d564ca7f43bab91a68474c9d8133795de907dc26b41dada2621e0fbf75f4e33cfdddef1d0aecd5b9ab8dd3deac03d6a14b7c8132e4e9f56ca92933bdb9e7ad10b595725380288de8d1ff305a88afece035a3df8c971c401987602e1bc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h60ead5fbacc73db7ac19b44c228b62abe6ff2fa6772f6394d2d52c5347bf1a0e32cad5ecb2657c005823b462841581b55f0015d8b9a3ecdcef3876a2a7e15478201a2cf240af6d4a12110e9f24b886673fe71e4ae8223bad400e8841ea16e3b3e3096b21cf2139e00761517a59c5e8813d9fa6b4e0fe8d48a2b77ba935b6b73db0dcfc4557a921f05032da94a3ed1a2375300c6eedd6a8b8cc3d89266917b7f1fbd722dff790826e1508983d03646d491ed119cc9fc931e2e24386f798c5cf57b72da59d1495c6369eb46ca09a0f058770e34221c8a33fc90c1917d943578bb20f55846491ad2ab9b2134acef910a8fdc5dd88ffc208332eef07ae95c26c0e8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h24a62a97e1f4eebc92c2e85fa28be7f83c6fd08b4585cf16a904791c655abb73cf88bfa332163ce4ba78e6843b8ba1db7b6ab2c7bf9c7908870e9a40f8e3c8dff5fe82d67583acfc52f74598d8f5f9a9d921d7eb45203d9e401a492e320fa5e3e16354330ae67abdcc06c931fa6a0941920f4ee795e1985e4e39bf9a863685d072e7dee1d69f88c8dccabaa6fd6bcac22e20584fc05a39eb9dc1e8ad34dfb2b236a8bfe81bd10774e94684314000f2157c7f455720a58ab6b7dfb1609901981c3e719865eb52ec1597481e2795dbb782f7eed086d84f1a7e8e12588a779c7edfabc8f7d0190c4efe771c31f727853d5bc395eea6903cfeaae637f62d614578fa;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hc85177c04228f47e48fc11df55e0dcf0e8afa490a75c922ebba56b37e802b836aaa8b6bc18ae5b848db5b29c2f0d9d929e10695fdbb7839f33c86905ee957b50bc34fcdf5bbe97b3a5247f42ed18723980ae15cab0a9bbe0bf961dbcb5230a418df19162acd33142722dbe3630929eed9a2868cd131e9174d3fd49a994d7b1236b1a36aa65cf41e69d627c4f35a1d961811974531d025b910deba086b70be46c537f3d47cd80fa48a055a4c8541a2f23c74f60fbb182f7b1edc8dbf914b5ac4cea10e9893975a1711ad0459213c43769ae8940680417fce79644d3032e945f66d2f780a75f9b46e239836785b5feaab2fbd39b46f835e30bd067d56b17ba60e8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hfa992abf8ae5e5cfc9f081da34679636e2a01947cdb237918f3d1c4408dcba64205c88564e76c929642230ef62f62ddccbe7b88aa92962cf507ed525626400cdc6e66fb1e8141c1799d107a182deb86158508eb84d0a5a61b1c8974b88cf3e64d08bf8be141df83f65c64b020b552e13892863196f34cdcb88c1258fcca4baccbf0480173b3fce930f68805f2657c66a0ac58487a8f6c385f72e459b51913f699b0d82e11179701d6ed7b245bff0f60e0257f96044c05c55a8eb2f5b4b02273c4bef0ffb4bf185aa3ba7888ca7ecb6c8833f90fc100187f035ec661208d703c308a22e94167df9bf4b415fd9659d8d3b9651a69bfc289b5746efb6da3085f8a8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he3942ae759af2282a5cce6d2aea4950381278aea06e02530c5d8736743b0d32201f9e8ab31d498545b4db96dc99e9f83b704938d4f3b1b8520152ee3074bb16a48ff8703175cf3822a8cce55a13b5e366a5170aefc4ea89e901622b5f840689c73388db7a69b1ea9baf349cfc8a778cde2319242c5b5c474a9d14ffe595a96fd1f48097f2ce3852ab70237ce501ebbdae9c4ff5109e0a386287b4f721e042e53905163054ae6cac6413a5f877f8b18ffe8f4b6bcf44d5857f4fab435c81d4e92558c873267cc1be7dfa2e6b9175ca060738dff7662a38927f27fbb8ed54269ee78b79c0ef99485e00b5425705e07d3f2957b639328a80b65c0837a69b93c579c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h373d7700785eefb3bcdc9ddac7d2814b164035dc015b0f7d05d9a45b683087fc5d404aa85c37704663200222ee36ddb166e81effce6e2ce8bf73e4ed1152bcb87f06662eb10bbb7f60f8619e48b031a4d9df88f9a1390cf728782a0411cac5befb438a2c48d5359b285df2d866529f91c02b26c87f652c07885b53fe352d8292c5bf4801ae8da4063667afc9831a650ed9eabc01e2fbed741ac9e83181b66f2003266290aa7681fe92796c51ca2d98b459aea6002d516a732d80fb40a34e85cb28eafdaab0e87731ec30fe780211ad04522bbec1d7c8416422cdc2f136a4579eb206b6e50468c88396a4a0a533196d421ee19f774a371cd20edfc62da0532a37;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6bcfbce7cb154085757d20047507a619443a84089adf9dd2df7459b4327c299b0603f1c6b8c2dc0ff0a89a9bcd864806c01a39865f562ca578f9d6a8d2b8f35814b3154909b78c281948d28fa4092fc62eaee815669d2c8a03eb3767298f35d5430511ff818f1f30ed41651640e9abac539ab626c3bf8e97f9397022a5f65bf34d53b5387859f9c12062cdbb719279642f916e12b932bbfb9058c8bdcb35e243f33e987aeac5b046fbb231e74055b9b226c01838def19abf9968fc82acfe28904f112f2dfefc98b9e81ca1340ee869749e554d389c94ff2c0974c12c7b396b20002a27ac681bb2f6d2233e6ffff71024318dbcec124d3e7f3a2c1793792d48b4;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h486ff46f886d6061b043f69b6f1a993a01e3bdec159dbdfc0150fa85daf3cec26bca0b7de9f16109680da3439968c2ecbd0c69dac41de91c68d259158bd9dbff74488a1dd28150fdf622324667f40a059fc4dd6ef093d11160c39dc431d8fe4c1d5775192f9090a47c6e25629b612308a3cbcbee3b8a71c141e1c091f5575013c24e0160de45e865e3a126e136544b5cc51f65e1adf6231b8733296d659442e3d9bd0f1beb683d98c6a3f171ef6c3e74b9460ff45dd2f9e5f62a756dddeaa3298700895cc1d7d8f83d6324e6d2d23011c045d935a336a403d13b2f490e24b779482ab0b43bfd8684cc916b65ba25ee0c2e8f92d356217044993d3ece3362c2de;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h99c348372080cfccbb36e6fb07d553ab273295b410c8c5196a5894084d79fd460ed06c4e69ebab234ee1d5ea7849caddc5160206e3b85571ae15c3eb579322748a944dd7e660f9666c8e5090884ffda7e6544f8af65933fa925df4fe98cca3a8e3798cc986352352215b8dfc34b8e06a031c59d070456220a0617aeb6ad8865104cce4b911afb671b370580ab7ee1f2a12833875b5a779b589b710cd219c445eb56b2e8b61a707c4f8dc62ad0246838e3c4c7e1f773f551622eed4b1165f4a0539a81c5859b809c9530ebfc69ea02723ee801fb5e6ca4540522a4390d018f995b86f99c6b68cca05fd91eea5fca4fc2c10e48c4fb926d7f4ec9658c251569830;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h240d88addd771482bfd434573beddd3647334180b06383f0ecb1fed2779b2a7a64448e119de1300b076ebdd4bcf6851083440b1439a1247a65001c7bf828299931bede64e5d9b426f90bc9adca3e676cb473bb675e82f87c2fc2acdd6e3f313a0a8b5736c9a79a0c0204ed0fb40c1518c37a554998e5358c124af89faacee7dca0e51ba1a6246e72700909af2bc8ffc1dd90d0dcff42196d52f35556263658fdde96070c801ea7739bb867dd15959f0e98e8b621b2d917a32d4419a5b0be7e69f00a35efe5e95fa55517245a281492497cb753b7e7ff6790e2e671157b44a6c08415a24b08d9dc2be236278db522479f1a9b89af53c3a6369e4b45c3ca1e27ae;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb2d3e8ad5f7c06c2dd81f2e8b69e20ac8ad770aa952bfb284243e4c69ed7af96946e65a22c1f9effb54173abd33436aad6cd9a128acbaf6706abf6bb053f4cc22b1ef68be8fc5c3b3e20bfec1a36be4d93cc6bef6ec54155a7d5bdfe15880f9c73be19ec8a285546af1c7c6847a872bc20e40504f13fa119d04b2196eed82647517d2ba3fb2b55c5968e27612ad523a98e07138f1b5cf5b9809ccefe486e07ea603642f0f7342d8d67d25cf120ac9caeb0cab697e1828191a2b1e20f5763442b73aaf4b529bc9f0c8961e8e046b1bbaa0844f2ab5be9af9c98a1b436b716194bfcadf1350af164ee95c7ba72eadcb10b312f228624c989eb135aad00cd249e63;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'ha2e32d71fdd9aaed9e07fdf342102d1e777dedffa1bce05022affaa69f4d35bc52306aae337238810802aa6ae88dbfc15e8e36b1550d3a5ef95fb3fe30477b08f6071c6a0c191432589336c78596aeec1fe093cf7e42ecbefb6d8b8da0770b948b9ad0e7988cb767bb621dd911f7c89d3606fe5d44ed0520ab6d6b7aca57a9b1cbc644055fd02d8c127115bb91c5b8669fa1e209ead15f0d9bc5f70721dcbf6b52ed8517a0cce3a22f44ac9d67891593bf51f66e368da7ffde5eb9083aab201f3390856b8651325b96bdb919c337205c84258ebd350e769f791293daa9b0e3e975f8dba4b90ebb2394a0cba8ad9ff697edd658b5357278aac857a60d1ad6560c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb3e084c22754f56679228feaca5f42e33e4a86a70c01677444842ef63921cd9b28955875e92e68ce1b867fe9a6406cac2448a47c6d195144d174cdc3567f791457cd92269d9a7e9c8eb56571e40d778bb733b0acad0a5ef87a07de0fdf440320ec9b38231adb55838a9b588147660a88ecd162ea4b961b1634c494c8ad8deb5ba37ef9b787ff3750463ebc7672b73196ed2ca3bc8a2d5484a1d7a150e730f417cb4da256a6fcfeb97e4d6154ef815182400ea8acbc958bdc7267633307dba19730a1d655d6ac0e4d0479e6b3e442e4efb1c735ad028b44a8aa6914782ea004c1d17424ff00fd620ee1b552d5377ef45256ce71beeb7fc6c45b367871706acf24;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h580a2c66753633f56d84b1c5b7c84ca609c362be409ca09d16bb70b1deb0fc3274d832645218b4b7e1ff9e52e442ff645129583a44161bcd84e89cd97e1b23e5d65a0c738336d558c8ac82a89984ed1d6b7a0310115dc1be5a6d1cfa3c6b8d15bb3340effdd86953dd8fa011316e208043c1004bd43955f7fbb89e38ee38b9bcdc55235f33549492ca02647c3aa5d729a39a35a58e04a6862f7ab5cb7f9652afe5bdc98f863446f229bcef023daa8599f547e2feffde9aa20a445cd6cda0ab77a60423b9cf67eb5f92a407bfb577436f62866eb28dd85428dcf91c8acff8c5a0a0a43a9ab0cdf88f8df1d2392c273a50580edb3426b0efa3a04bc87abc715508;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hcec4ff8e1bd3ea0bf9e17890950fe279a29dacf489bc529d3472dfc4a77a49177822da92c3b26f30938d4971a4bcd03a0d8ef4ca9a680ba077f9c1740b03d9619e43b5379064519e3cc7bc004dab625f4f88ff382a218834730690b120c8168fef0dac18cdc55050f55926cf1f9a651599d824fe514b4e8f15638cd6dfd9ca970d59330cbc0430bd89d62dcaf4b332ba091ededfadd980a397e36f627f489c2d1e156210927b4e30c4cc4937d405f27988353ace0e6612a7232e155a6e1bfcd7b150dee9d4cb6293cb27b8776574a04af97ae479824e17a67ef298ed49ce9bb693f7561d1c4864e7a4fc2db932b564cfc155f689610c4e76e952ebc6d2bdf335;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf977d4075f2619a2044c2a1bab737ba432439386cf0d8dcc546fa82e74fdf26608e68e2cbc39e2efc3dece509619fb662f521bb5dbb7ec2f1ad8cffe9942ef8743ccb8ec1346be65a74de89ba192055531cc0952ee6fa478028b4e433c43151ac33f01beb573259e25de714b4760f8c1d863b36c46024f3f931e103fabac9f78b9d33d2cbd805f328bd127cb161971eb036496f4e910f004bfcb3657733a2d7337b982b0199392229860c920d7570f742b805e3c8a75ccdacef94b47852d6b5577dd237afe023cb3d0198cc011dbae76bbec08f583332e45040dfc27bdba874d29ab99b60022e4247bcb82e9a1c942cc0e08506448ecc116adb15dccc6eb5bf9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h36968b9a0b009e8d4ce5f9f1002117be5a7689c7a886caf6cc0d3d8b469047aa768840ef79a955b42df632969534050d621c1c519eca37467d48561e308c6e417c65212b2b2eb3e45a91abdc98cfedc43ffcafd02ea0c10a0b59d6e8ac39a3aec11ab6842f2fa362095eba1d25722c8d7dd40c50495c8d242bd13995fb91ef2b0c98ce54a1cd0f52c34725cb240f9d7c2a2a205082379163ef7755b362b0bd194474ad6f8afc48ffa6c3dbf5930f2ca97ea8bb0399aaa489596886865db8aea09a423a60cc36f64e7d807f117e26bedfb4db767912a8e5c4d4f078bdeee0b92ad03342c54b9d2a0374a6b6430d442bf62fcc66581a1fd45a9d64fb7220c41d8d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8f7ca5fc6ddca0e2c4b695c47261497d5e70565ed1ca444ae8b2769dd3cc10291951cb85a5fef26a4f7c2ca9058136aff0818b27fa4a5cddb0f4ee1ef80d3cf3b98333a2b156dfad37a9e2c126f4b10d38b67f63f97aa22fc7468d1551eefb23e3b3b075a56a3c2317b1a7bb7f0cb33157ab2bc27db39bcc512404ac4345f65dcd5b58cb118ff2beb8d5fb529bf599400103a4cf664b2e7c15e898327716508d8f90d0877b4490ca98014b13292eddb6254c170d56b7a33681e161229b0098c4ded5ad2f9fd95f9400df4d4f1c57032c1309ea58ba7fa05279a8f8fde8f408da082f52d4639164fdd3870578464f3dbd9ccc918773f0fadc3f2e84989ca13721;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4c389f324da2c13161147bc34da98ad9756d572a59e2780912461c3ee598b213c016db7505b13dd1cb33b70442c6b4f2b444581ae1c1e409e61881e27f5f9aa1f41e74679cf172820e1a0d3209ada241bf79b7298d415397e811921adbba2fd3d048f8cf20f3aa76dfc7ebdad356c980fbe9b3129b29bcb8fe480422c9a9a384881c8b8cf891b21d461f8d85c3cf99125986a8c6b6304880e8857185c51850bfb9214d22d7be6e93c576dc72a5785507f93a21845b0a4a9595a0d86b1a99e7c43aa5033673d64afe22e251509cca059be42af0af78d7292337f9c5f1134a8138851105d8160433e19e57c2a503a3f74ed83cbb74edefeb69f60c2e3097c668f1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h15afc8a3dfa38f34fd81442d6e853508d6e48147fd29d1f6cfad8d375157ab93ceb79b0ab454c9cee98f1ba6f061348bee94d566834ff7c5679b3f107771568714135aee69c98607435ea0c2f667132fe6ce0fd30f51c704594ae6a86ecd53f0c83b373b99ab98d6be96b037af820b30d07a4be6d2377209fb8c6e2171da0ed1c56fde679cc0338cd73c6950213810c516b403bd5f7268d6654e3d59a0e8e294caec0da26bef2fecd559166a04b27dbc92b47e9ddf6307066ecd0e2ecffa1d3717d8ffe9f645a8ed12b00508bd824b42db917a2c15d03dc20b5f2cb2d128b93246ac3db4906628e27d5353f9eeb9dfc657468fe66812c2a4b7e62d61503b274c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h305a600f78a9c78d4b33c9a805e7733bbd80aa5bd539c5528af7a33efede4de40e6bc0ccfee0110273bb6fc7003ac4470465f330884dab44a88010ed313dbf60fc075045a0f102e6b73d1d80476a4865b5aedb4a4cc369b0e00b7537911da17ba1764ad8cc2455c1748925e05f317efc810a46864a3759eb8e779f33316b62fa5c50e16139b8317323d979d68944b1f620b95d89d5e2135415c221a44858e9fb5b90cea6e4a3557cf2df4fe1bb271503513caae5f9607b222b00332968fa028f3c0434beee24859b82635c23737ce61a7fa7a0314c8808035381e19201cc67eda85497272fcc30492ee3d8efac3bb10ea5e73b9dc73c64e2a16fedd5c040d604;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hbfe0a32da1a6eeed99d4dbe081dc934e926994a3128c89496f84eca4ed0ca92e11ce84c0a01f9a5cb01fe3ea89c7f3d73c773b479563c445faf44ce03165208f7a9ed7011b335453bf2bd83d5986df40f682fe89923212f1b31c10d32fccd76d4655c808e991424dcb28fc5551fc11bab707880355369869335c2dba7cf5a674af904626602ff2a468659ee50947d7d40438f3440a593e7419e4bf785d773f82868977366748c60632c701270d3d22017f651e89f3452c379c9681844fe6c14de2a22aef867e0286541acd3db48e12266079d99ce00991ebfe408ad2821ac26b40dbfeddb7e412114a61aedbc035e4c3ddcae68e0b546062fdb3f3212bcb5314;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hea8ed272013e9cbf6ae6bfa159073362d7f7b21329e81ae85c232973fbcf1a93caabcb8cd897d13aa274674f7799829d3ec54ba7e7d7d2d32acae0967e46d106488d5f17e1a05380c889f3361aba66276ac079e47264982f54f296148c93eae39b3daa949c1b61b12ff47965491a33d02a5467170adb47b62d95fdf91095f91c96bc2981f017637c02302eae292c289f963649634c54b1f8b835149aa4ab1e1508d6fedc2aada7f1c6426a38a4137beb4a9e21b6e13c5d31837e2df2aae781cc3667bcdc831dfdf87b3f957f309784bed9d511e52da80d57ceb0ba524db834b10ae1fb84bf0fc079849d5ca76da926e830ae53793618331d1edd3a32ea8988fd;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hbc2892da606ecb2ad3b0fb1b3d918ea8bc7d284acaa864c8d7314939408f15dd21792e444aa41ef46df855a59d47972899e5911cef90fde2e917d72470aa68ae42292969eb5e03edaef4ed6caba33bb96faa0840c60963815ba0fef8f2c110c7774d3b2f552d7d87dc3555ed92fb9ba14523d83e3f872762c625db3ff89b37a10562d18aff22ac805133eb06f88557ed8b288d0b2a79cd9ea490131f2659e71f403262b855799fd9674d5f581488886aea15fb3067d37488ebbe16a9c20a6368eaa92eb467a0cc87adb0221a6efd3eb56c4334534694d6266113083dbfcb209a03cbbad714c57686358fb9ed6e93d3e8d56bb244b001d9b7accaf2ca573f7ae6;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h979232fa818a2ab4b1cc7dbcf2a7aa2ee01e9e112586d4298143ee3acc1d70616be6728ab426a0aad859fd1b6f18d4796beb67d427ca5e1f8a5c98b5fd02883841027f655b8d0c7903b13a556b28257d8459a14324f0248b66d8bc5d4e4058a85a8c88cad8188c9080003c4cf03f6a14d4893a19d37d446245c79dd99d18045ef25f6e71664ef4d5d8cd923940c449d8ff6f5cafb161cc1bd973442fac494f2cff961cb0001b695b664ab4ff9e76c1b64e844b852a7764d1af691869783125931000b67d4c755aef68ea100cbcb29d1621b47c087e566f5dc1ff6a6aff8bd777b2f6e18af7b01526fd011dc9ea2f895fb164e793372e7b814fb6da5d630a6d84;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h6d5581aec4a2738bb70f480cb165837d319415c7e4add47b2f6f0b82f65d03aa0f6d39c3e89e819f17f748042359e3ea2b43397117a537fcaf4ccc2f0cb368152cda5999b0e667078d937b858bcc6adea78512cafec3fead9cbb9b9396d6463b552f1c1a5b8abfd468e0705cff03ad5e7086dceaf63902896e82ee01868b6ca5af76faee1a7398f373061b5b90a145ee206909983028459a531acbaa37bbefa9ef85072c641cf5b2d173ef4455a68fc52aff9e04c339167c5dc270d9fd3ceab1d7de6567c6113340bec8314dff9cfbc61586fbb95870cb1407eb6ae5d0616988864355c0a4c18c444f2306f9bc6e3f466e816edf4d08ed4d569ba02526eaad3d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3e08b4ed0b1a6e2fa333d7c576f08bf63a6c5bed51be350be3524b469c92f2e9ea5d42d2b06d011c67555912e5d5aa92f46725e0dca327a6e91d89b586a043cae7d754e08ce902fe5c5df2943ced0fbce9697597ee9245c296976a4e59cb173550840e70a729013aab2a5140001374d5d0fc8faf159b12d7700aa95a262987d8073d727e9ef1b208cd0c0d6f3ca7a95c88624baf193ba423c353ca31f240a836d4277dff81901ba39be9468fe2e746bcf7a110663882c0224f2cdbf7d187478ed28adc9c52e57ea80dcb6ba66b88161e62384508eae3da18963e4979316368f063732fb974fc8384eff6f8dea69405b409ff1d02a4d9a0db10201251db16cafe;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he1941b06252b8400fb0fd212c8d58aefa5a945caf63d3356c0d9f17ccf3f42e0df79e8cfb64d63573a48e89f61e818de2794646e10eaa98e1b80c3fd2d284fa72c4be4b9270dcae2e9852ffd96b1000323d9693a59c6854704bc8d89ade82d9b76f526f10970c1b07b1a6b471fa0772de6f743a092be3b9883964a3c71880f855add75a66830d7106b3f5c10d45488d8dcbd920b94e643e2cda9f6729e91f6c43b2bb984a87cdcaaba0ecd8f0fbc5250e9bcf995069ebb3f1b793ff157af1205cb730c36efaef3bf9a4979e4e5ce728e9550a0b53ecc1c47678f0883736e3f42e47d79903fd9cd7c16103d3e315f2b341422687d3000cdfc88f2f06bbc0b48b3;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he66dfc7670c4936307268001a00e06536fdad3e701b4c3e16348066fd61efd797f46cc1cce491cab008b5e11be4f05233d3f8135ca1966bf29e8a31279c14866f5fd4fcd21d0237b492c2d835f477c868dfb68dd55b2226e02ee6dbb33f4d8bcc46378f0b8bca2b3f4881e595b537fb84d104eda2e006612e668214e05e930403c5c1c615170a985489088a7d68d172c4316a96b67bb571a688684f7cc6a937277f5c51ac2e8ff3728cfb274b2f29d9468790be893c8c15bfd4f714f2c590468a88221d53fbb599932b4d0940f763d66d75360b1ee2d82ec2fc291bb3febdb178c2a90eeece1f2f5c56925b93bbf5bdd7c06a15259677c9088c11caccb513266;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb58002872828ab514b4040710f79a24eebf8ae1a079251ce8f2a9cf6330eb9b0d110ec732df2ea62437050d734f66eaa82c19b0c94c74f7e56cf31dac5923a7c6dd7227d7ff7200e70c990e481493bfc82177eb517b09a49e4cf43d4427fc605d6cd4d8339e7e5abbae0f54cd055b3737fb90255214cbdbc1fe92375f9dae1cad388ae008f759bda4ad920dd4f27a975b2b63134041ea1ce63eb00f11405d47d1d3c1dbcdffab778f785dda6a9d2d9b0f3ba8515c181c9e83ae57b4b7ad7b8610e4db1f2adc47cbb691b1f09ef1ade0ee41e4716b52ee7c33b6d3a3d195eabc8c5e08c5d4f9ab1a1b4c904df302a6bcfea3ffa3e7cd6454faecc089a3bbcf6ea;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h9f843b55adf9fbbd91850bd4f52e2472cf7efb56c4da60eaf63513ab70fb7bde43842f5a72ff47bf6493c39238e1730cb6cc54e2db9f1b696ca9e54adc2b3b2d04813347665d1cc70d1bc8a316fba194eb00f4ed30cfb266bafe62685036cd120bc6848fbf58e53a406acdcb3e7def2b4c20240c974ca6fee2a4fd18cd77661758494c3032c1bee73b14b740da01225952e6883c8f37ab0250192461e24a0db4d337a77dbe079653eae68a9573bf78e17f49b9047f0f4b051c1173e4e6085c0c88b290a8a0001120b66a0f1239f807b1acfff0515596b7a404a69e3ca1c26cc8eb1b173d9fe615305513cea46f78803ad02d1c2982586430f72c04b39e460322;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h185a6f853b2674723fd8eda7c8956524d8f0e0cb93b23384e0bd7136d39573e317288de778f6c34d238718a042c4da551bc46b3230a0bd8d17385d4b96d073c2eb6747e8d999c53e4bbd3d730a100f6f770d0b8f3494cca3af6591cf3426880cf6d6b2d6e3f99555b156ee04e0d2d1a61f2f508dd19aeca60d6238c80785eef25e646f4810677d81b9b221f25a26d96f354eaffe95d96fa64a17673b7ff4d87650fbc123c70791fc94ca8092ea825eeef4b64d282224135b9eb032b4a28bf54f7280661f838e3f7a7db005869059b0e1bd7ced86ae241250d8f3b9219c24df65e03296cb4abad337cceceacf3524066901c80f5e02f5b2223b76fcb89d3d7d51;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf6f83f841965e2bc9e1bddab8941cb308b4db8d44f9f9cea925ea452b59f0531ebc34de3ab6450db07b329bf5305333dbec21de9ea7132d39998e08cb3e65467850cf3503d7d36b9f7a3d2b91e3a26dfef3fbeee4227cf49e60edd77612d450316f2c47ceb665799d70c736879418e51cdda61b2780e46e08c575ac435a90c33e48c1e35718bca6def44d9450f6970d0ab10c75b380df38845f57b2cbe43e25f38e630cb02f65d933c23c7f507a3faa71eec569efb52b9efc2f9c2044d1c6f379634a2013dd0814a44cc9a6b7f107fae59617b88e2887cd867ec604c5481b85e37d3c6c70ed81f7b35da848db5b3155e67d13804db13e5a4cd83c5f962d7344b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8d49eb813854c743e0a3c80cf529920182eef635bf4b12ebb134a68807d68ceac054108587e11cfc0f66e234b9abff88226fe681f947b90de6281d3ee72a42b477e1266de761f3ec2c103ad7c53fea83ad8082bb2c03cb96188fb8b431c591be35c5afb8cd2c9833847cddc0527f3b1b3c749bb6bf5039f8556b399099ed98987df19ad7edd950fb9be605bd00750fa32f38725a897b77703cbc74564f5354391902125333fe8866fad49807001d859f10e86fd0ca6030bf435bb451a4379c99d6c138c7008a0b938b438be86db13d4d07596f7394828b58ffa613d9a98adb3b0848d55e30426f5062d6b44aa8a2690b2864e927d2bafb20e4bd7168d1323a8b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h301aab168cad51029004b708d3f65fb6ca144a6c9de5c492cc43e14ef887468689a1391166a8669074fbd468802dbaa6b9b106df3efd71d4d7591bc290ef7e3719e77a6bc69de2c01011792c316045d54531e994bea11f5462b5382e96b57b0e66de668b547e0cf38fdfab1e45fde42ab3ff5ad16257ba7d4fcf569412662d07fb07bbac7852d74704d9bdd6ce809ca904a1b79f6dedc0c0704087b925c6cce3ba23289fb64816f2b7b7ceb738a1c289ca30c57e0f78905f227536cf06c55b54ada63d4d0c6fc199f546eca246eb5ceaecfd96ef3cda24d7d4bde6b277163b095df6b55e17e563941fbf8b81c644c83c181e9b788fa2c2a2e21e2ba946f24353;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hff76e4542767d073a78966e6bba4600d5a1f826fc6f8afffe7bce0423c4e17d8b0c0847c93951cc484262a3d149402e47800b60cb3ec111e81f790866402edcb89c4240b6668ddfd0869808690f0418fefb524b7ab4a2f7aa02931329601a871e54fc45c267002e6ce520a27668fbaebac2efbdf9414023c662b5bdbdd3268c0d69970e0b3ea29f227dc078d18f8d450786a8251662b66e483422a5f87bf93592178fd476f5d8a4f60cd59c9e078d10fc583580d87021fa641a22020dd8eb36b6235a16e3e3fb659617f576d7200e25aa66849327ec7094303e252eeb34fb607909478ceab01ecf2a32dc923e64fd48a494c4a81bd28846ad2b0a8c532f9d828;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h2e301aa8786e6d5f08d7b71a17c3a4c2505302d185aa3b50d02b980b8f4e3b0bcc5888ba25c15b446285795fbfe8c9caaac59553f3497302140952dfcf3e86689e8551024bb3ed0f001069b6647dd0ce51ad90557ab40db54bf0a3774796dbcdda11d84219e8b8557cda8f6a0e6200a670e04b2d67a635a82636d18edd203d9536695fb357eb784a5bd9cec2265853e7acb7fe44840a8978872f560bdb41b420ca10c90625743698774f6763ca327156991b3698eb3c3476ffee8fa7dc8491d7613407425e26f2e7b3d700f0bbde60c9be04ccb8e9a979d2214e9e71f500b2a3b6266b07f2e66c08223351e5803264e80417018826c0a78673eeaab130543abc;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hafcdda24c9297d43e441f561e15d3f3757e427110eeb6b868fb95eace93fb1778a9c7389d0b2894213e84aabbb3c63b7deb5f11bfdeff9dd1bf98c9bfd8624a44f422f3e0d22cf96c8b2fcabb527bc746ffe23dfdeeafde04e7689d8e25b15893df938a86bbdb75225d56afda42ec3e4e2f80c81274fed43807b6dde56759f9d37a011ec08216436c8fc301f781f2de69bf80da4378cdcce2c69b526b4d6c7db370b2c6ecc07769b6991dc25405f7d80d1a6364bde24b2b1e3791cfad620a33d3883fb79d8149c64b8f3129c1294adf910b7dd4a7aeac354006ef9dd17cedf4f9e018888089cfac267f09dcaa4e3d99fa4cae286e3fc664ece6a0e0d55375a88;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h67e05ea806dff2f3ac04aab50d59f92f1a9fa03c02b35c651c07c1856edbd0690b2cb95eee1cc8e0a9658e75ac8e5cf7a32174507dfc23ebf99fae4ac52528a44664dffd5b811f497a32c25472c1c6e6c28e94b8f8c8b0197705014100e7932b4c8e0fba8c5798e11e750ce63fbac1adb9775b677752b9270db1ffd946d4a1271b3c7a857fd4f33fc47088c5343718508e13a54fbf9a97d4aa823ad1cbbc7d10aabba54e96580c96c966e2b00c75bff17490846828304b4416ff740874fa7d7ce0a85d05186749a0df61edf0f780cb3e8850e2a65a9ad4d6fe92d2026eac61aaed2a4d3f76904c00e6820f20a0a1055008e81b846ae9a45f1673395820370268;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8157083e18265de4206a47735497676f6202b23c0ea037fd86fd701c07e96158168b5f9f9a5ff8e6ccfa145846fae7cd2fd0831484e848c773fe7ae95ee24947ef212ffca8df3bf81bf180c47cc7f6c93c7bd791711a9be66d4e1a0d7f95d454c277b9e4bc93003640b24085f3cc306d5291f676aee711c61d13718fdfa4ca993c0fa2d5654a6b55f05479ced8ab9ead82a975dc7b41f3b2f890c37bf5557d7505900a3e7e61d6936b981e947722a46bea372a4ab5f429634d32efaecbd1f438798d8759177ecab8c55fbd83453df7ffec9a8ce4f31b25dbbc73c96aef4c64f5294e3c979472c3a37a2863f7708335e678b6d2c95be60033e4072d9c9c216c29;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h7a555ab040c13dd9e6e9a7c439405cc0d8ceec74ad6d1884bcdb7529392cfd2a54f22b337c3aa4ce38c56f15dd4a3e8a879d3a6f9a942ee02837c9a89497dc4feacfacb26092cb75bf09399fb153f7e68610a059bfa0cf7614499f405f75b63762841f565c31d26c8c287c401061177595afbcd53aba4e44edf729df279d977b9ec9b6430dd9375d7acd6a29829b0382ea9fa2c27ffa0f331698b51ae1e33bbd9898f9874956585b9c397c18d3032a6184dbd71fd17951be5832a22934cf61e3777356f4c0439b5dafc474cf6417e42a9250544225de12192f91b7aa3ec72d0e99d79200a01ae8b107bc7b9e67dbbed1f936fe26ee084a3062daccfe6288e9ab;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb945870001d753e04fcc48e44919160d8cabaa21dcc41fd2ecda0b9f098091bae2c13bce12068f8e105f511d9eea3772f856c5cbccba7cdd832ec47d3f4e7ee6063e61777ed1fdf0baf8419640c11919a793c39b97057b593c2424df62658f66082c42bb1b432fa4506710b6042a3f44da77be648f43c99756a9911bc68e8bff50a87792955f0ee9fa40f2859dc4af643f0b82df244f0ef1584293cf7fd6ee178006e879b7da04b79998905efdada15a85b624bd47c7b317d4b6d709740e673598897c0f27ebdbe63ce770c6e174985eda3861f39501d9a9ac84f6a5e706b10dea877d6c9fa16cba020b768616cae077236515548cdb33ed3d71985a4937031c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h28bba9ecba6d10d82802b0e705b011330f278020eefabde88c7c2cc78add170aaae219aef5b7b3f6c35e61715bf20167153b20ab356ef8b4f55b78f67840e931f7642d0cf72ca3e4cdffc6b5d99b0b0f8e7b4b9cd95f77e284f2c651c34e6eaa1b0deac59486174dd3decb5a0d5f73a3f4e7bde8cb98205db4d8bbfb01f93db08dce52842b0dd2778beb65b2ec293145954fe349fe0908edfdca58878c41f2fcbc3c081f6a235141eb868e35eacbd720b9af83ebaaf14612ca73f03197fd4d8deaff0e9465a418886446472f7e2ad3bcd7b1852970b494bb60f51e398a43abed631c79e31771cc8470a97dfed1af97e1a326b39a5e39eee19775ba5cc34bedb5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hb5eaaff3e161bc90568766446de2c7ed7db7370dddf102a132b6419d16d684f3c813da2ef5e0e1d12e1a33a0802055a56e34fb4947d528b5c0d29ec903ff07f1c80b777cc8b7fd712068a4d6408a24ba895e9b23dbc0d5ecb210451655795ba0589a2bc08521d66806ca6a478ce6be9ef5f3e7358d4a3cb80e489a6da2f51898f60e3f7fb24453dc69676b6591fedb164f6d933526ab15cc71728076a8536b99d21a0d34bea2389cc6cd0398a508bad855144f7298888e601c2d7fd9454ac6e7f314b402add8145cd7f7c0aa8780d9d6c515a420e8da6a2f56fb4cdefc609295d55e42f5e3843cbfa72929aaae64ae984d24bebb1e4e4274b11dad1d544d469c;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h42893668dd04d1332c72bcb86a18190af11d963d447bfc2a71d4c2bf3fcc96b7de38cf92713057ab0ce9b7ce7e4ad471ce3c3e79d77611682a800917c0e1a49af046406e067f953392e2834772a819db96b220f9146814c89fa732823607d971dbb01bedde5c0d810f39a68c36dc0cdcbf67c96147b110106b60916c12c00e5a1589a00188509c4e8a65c123cec2a564b3e1fd8938a7897dd3b187acb96494bc87de5c2e62202fe933208738bd5e046fff9736f00dc9a2c0b8a59971d402723269cfd1da2b86c45931d1b670318ebc0edaea4a20ef60fd9317320cb5b0d424b7679f15e8bb74483ef57d68e2f234c3ce941d88e59841a6458752e134cc68640e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hd6957ef92f386d297440575266d2a8fd559bd6eee79489e71abeef98407d9942dc87b46b84388cb52ed4374ab123989ba95323630f9a4848d49134ce3e7ebba347afd1b7e3524c9dc964dce10ab4b1d1f3583924e1498ca1ea238a5716af94d8d8d326edb662dac29c3deadd9fdaa1094f221fd51e690d723fc166b521f6273753e0d157bf73980d3efd13a68945d1ea52fcce1b1194b37f3e687dbe50d3f03da29dc05f42ae1b43c06ede0ddf8f88df4631684fcc77c98c36a7695cce3c70f5b175d5ca78fedb27adfc98f2867ae0e78f92113c6cb7824d99ce33e9e38b41d06f4a209a15eb933926520945ec1af398f282b9c48d325a61404b0f32f7415314;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4c7d16f3475ddfda0854c4657937f563b6a86f87a919b02370d4bfa766dbcd7375085f0c19db86d2e26a1ec089af84ace359891e391498d6bcf5fca14798a851df2111ecef0795fae9456f58fdb69a719fd935073ce048dd40f58a4b5553b545f160382a8bba128d93294d409f5b8585d7645a5b489b5a7ec5571b0c17e62dd10f86c6ad3232692cb5df756a88e2d695314866d5b2c2247a56bd78e8f6d6b30ebe7fb876c1021990d1bfd8957a526ce1b0a3e428082254f61b662843efcd440806cbf685ece42e39b529cb01cb00fecf819475267383705ff3606d24d33d11361b65f00fa947312df2b55cf935c60e46bc54a3232612d56fa98d4ce891abe56b;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h652f6717405a3631cde778e82e79d8c8cc3d538827a0f9f21c2dc3ef2557a7c2eea2ee0fcf0e90926bc94631927dc313f7cd66af1a0242c30b7eaf0824312bbd2a91a4787fffb650a16be24567f46828ed7419264427ec65a0ab04d9bafcd2fa42faa476e53aed37375beb803c11b23b3d4bb3f5720cf8ac15087dce53e6de78d42fa7aef973f292f662d7a80dccff5d5cc39d12e68598bad8a2d3726cfbc391a947176a0184f5b0b469bd92dade88fdbd05428a74d51eb567608216630956c794f4900a3b2add9419c51c3ebf4c29f716dd9fed5c4b9f57992148dcc49eef0923be8f2d0aa8341e84e975d3efbb4df97fada2d0f040c046f9ac7e72ecf67c4d;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf68c98ec59c685a7b122412a50a5755af7e3533dae809c52c925fa4130721ff35b572a8c55219a1256a3ccc053dec2ec32197b423c562c1be6b4fc1e454f3a5e9b3b2b47db8908319540ef850d2012971346cf9a77810d1f05205312d8a942054feadc1b5920809ed1e6e8dc6dd46c6a4fafe575dd477a40dc97b908e8b8629ba0c3be81c302dd393ce46b096363dbd8f5509ad987dda32c91160e03a0820aa5168c7a80d6827c3a5430ab67e6dccd2b0dc6d175ff64bc8b01c5ad2bd87683769ffbab11e27ff235f5ec8f07e406f5734076a357e1240b2df6430c19a54398eee607ad6f752982fc2c7ac66a15b878ce8e5b64335bd83c06a62697868f0d7842;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h8fabe7b8445c625805beeeb8b047be8069f389cffb15d645c7de4f76c9ef7a773ea9ab69e8a37edce4595750b1707050009b8e2337e076c79333f0645fd527358d243aefc8c0b8eda4a234be44a8bc479f55fe33b11e8a455c87a07b01e4112a16aa1ff3d3b6e06dc2ba897f69e2b68fa2030da53ba2eabe2f0f3512626cbe4973ef2d601a0fb6b9b3bac546eac61df5d49d5d034b7a092315387283a4bf0c25d2708c53078c068606603a82da8e19f8822058abb10b4fb31b6563e052e3b326d8c8a81689fdb4bc73697bf24e2339f721d909c4272896265083f896c15074e2f687e582b0ea22c48a84003a3bd588d72766bc72b93f3d8b743efd450fb25897;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he2b1f2b7702986e0c249468156b07c2e0c20e5ab69b8ab01592ed56fb2cd7fd41b332b14ebd665afbd443fdf8746fffb88acc09f5804f0d054e571e78154532cb6108f474bae7dc8428a9291707e8253a9603f524c415ab8cfe781fbf26ec38e9673ab32d1fe6df88016fc46dd1b3c4a75a53575e570217e5e8c1c234a7255e98abe81413810faf4679f2262425bf740430d6aef8e54a4682557c47e85449ecefdd65bb1cf87aa5d6f265a496ab290d9d3db302c25e68953b7ddc205d02d3b7f04715fc43705842155efbfe5e1a184b7569d7cf98880827aa711acdd2394fb4a5a86c253ecca726998b71ae8277090b2ec5fcd85c03d11f519f09c39e6d4d5c1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h93421ef62d55789e33a179e9e5e245d7b7d29a15e346339f81cfe39b63ee0cee072af21b6d7eddab0cc64cea126901e0359f59ca33b3c3e81af4ab035171b357e49f7836a8745e25ab1cf6282b8ee0b599eed3b12f6a84cab00b3bebd532020c788de11e1f0dc82272c7eef351ad9eca3f8027597ad886b9c0f7637dd8b646b93cf4837a3959b9097493071f46ddeb0650afceb004d87ed6892c209e5216b668e06df835c29605a48574a986a18cbabbbc82f3ab088d1bdbb755aae8beba81834d495bf5f6b577d660147732cca2ad7bec134e902651fee3c1d52b7e5fe665a27c95fe079f6bda319d3dc53ff4736f8474d27658fb415a5a82fac23b3df5126e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hf21b75a925f186cc3a3d939eec0893a87af59ba2fad4de1b2abbd651930fc43b05e61f6095461901d69da2673a7f1baaecc9d9a93df68a5a10129edbf3a510327fde52317da4aea29d5da56159f2c847343e7374f49a5fcdff38a6bdef34a65bd363c5756370318d5513bba60513fee84c278b4f51734ff69c2ebf050ac38d914130022ed743b306169dcf8d02c3f54f8705d030fec3e27cce458a08e20b2840d3c24c5c8cfdad482f42b990744bc78e9a60ba483e57d6035c3dbdc097e09edd069ae212ddf5a952c642bd303bce937aa824822330a65f47d49af27259737425387cb488a7096c44b046a6e0cd75ff2418bdeaaa2523d956b8baa765022f2bc5;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1a9532eab3e54fb8c77fdce1a715f29298293fbf024692f8cb22b83dfd59ce5430be9dad6e7a13ab1a45838ad22bd239b346d9af4a671454c83d416d5ce18c36452d60b5d2d6194496d24f3c5c3069968bf7edaaa321302486325485602c11d9ae31401e4679fee930688c2b4a6d86b09af8e378d6293b556745385af079b90866bb4f992684f4e3515f199d4499c007b3218de538c064f6545136c34104ee1ab87df67c32f2b868010c36910ba51bdb5bdb5a9ef41c15f7f603d441855ecca67c158e6764cb01557cd5d404b39834eb5456b6b3cbf2c752ad48f0de9ab25509310cac6ae35863188b358066d1e143d08aac6bcaa8e2798ff362bb5bc14f3ee9;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'he0d8c200cd181e11ca39cba877d4f4faa1baf1b39adf719d26f46ea077a39b905ebdd59df3e82ba37085c13b6bfc9e8b93082fe8b9c8aefdfee222be843d3356be0428d87cc06293d41a6abc34f4ab4816ca7bcbba8bf13512fc6fa2f91123e55ccdede6a0ce83c5968f2da198cc3ff895039dbe0386cf82658ebe2eb311b5e53ef55b54dc9462e509fa386d6e1d19daef05fa9b8568f0769efbebf41591e6ad2852f373d70a999b2ebc50a1450ed55595626e04310f6e1f6ff0813e6c16bbf37f21ebd51d2831c1a135298f53774f1800d7c7f6c0ba9b48f911ac0a7ed1dab0b06a6bc869c89353e3dcd076f3776c20b2326ff0524323e01cd967a4f01f4969;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h4fec356e207e550456df4beef9e921a6b808e380aa856965adf2eff940cea9be2b6e73bb9c1835c7bbf3c191b45ae44871fcb1dbdc04defa652010ea35d8fef954b1388dbf690dfb0276a8cd1d8c6a15e83b3d6bba2a7624e90e343e86a3567cdd908d47e699be77dc5b7d92296e5d20ff1f6ef210bbd577bc3ca3b939d3f686da7070735dd205734125fcf353a6255c9834d577133393be1df22a1e485a450ecf06d4dcf14b423c51373fc19d661467d51fa256f52ba3b96de0d4dbd35692b153dd056bf31d6142a28714bb0f5fea06eec07e517912b88d3cea27327c77b87b40c62e91661dd615357fcd6cc500af020752c60582c736817eb57b141fc96dfa;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h938231fa6303b8cbefd72908f83757b00cc0c8c185e59e10c5287a0836a66c0bca073222fedb219e10366fb97b9973fb7ed3097f87cc2e14e4406b23e0a45a72f16c50f5809f19c9b686f4ece0a22243582c9e471270233017728e966c3184cd4d3a99b56363be78f836460e52df950825d248eb82d04b8adcb759aa763928f78845e6845cbf74edaf7a29c3ef38ef40deee80ced8279cf9163059d2be82ebaba15edde4400f3c276228bc960dd9cfed4f4d74f2f34a9506866f14f682dd37d426261858d9a1e28530d93a35d573f838e9f7f6f1d2c6762078c8d9fc2f85ada92e91ae8b2db9dd523baf6d1e6a19b02eb3159b616d940246b8fe1044309897af;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hae60fa145028ac38d5da40aef52ba4ee464536cce7c9c704ab0a6d4712e2dbbf089c908281c216844cf4a5de7a303d39ba2a140022da2a0262554b2cc75905d92a081ffee32c2f5bae70d5557517be064077cda12589403368e5a0c8ad2c42c8117cfd2a4166622f44dc2a780d5c434e12189a57ddaa8b3c1313882b98091ea707d914c00998170b25e7c2361f7d08a6cd4344c5b28fde0c0097a43f35e3dd4662d11b8fc1624dd5c429aed3acc2884e3e9830569be6516eaf484c59b0f65ea5f6a188670ac6bd98504d2adb88b0114e96e2722719035c3a7ce6ccda6171507101d8c94fcd0c5870e5072be57b65abc19d0331dd45c0d7e123db9d33f3bba279;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'hba9ffb50ed53137b03b10349f6dc8653b3836135812c9febb74fcfb9d2b2d8df4552950e343e0b937142287d9af08a9daf9e1057aa95ae3787952cdb9aed228f7e16d7db3c49ab6ddef8aca0222b4cc03225199043168180c594aa5bf3962bff0d7f7038f47f95b7215732cba4d3f20dc50bc4142c882c9fc9911f435d621ff7f1f62b177c91ca967c1cfc1ce969e140c4572822faef13edf662476f53f10b2746295cf3d3af8ab0fd3228c16b19e90dd3e5de057f282042851677c7eae80c472643a789fa98c99db96094e4370c5c4ec54f56abfc581690457a3a43c95e1d17e22b14f6ad4e8dae2bd15dd33bff00c7c2ebdfea36c2347071536ffe7c955f9e;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h385df3b12329180435b989303be3dce20bfab3b8e75c8343b92b811fdef61cc70276a8a27a1030531de80503e6b4dedd391ee02235c3cb157672435d9769501700795934e3046b1e92b74efa51e0e4850752b31f1a7b77be1a89744d262336d7a133a80ae94cec44591174672fc1b22a1dd5bbbe299c6a104a8ab9701b477e61c283201e21cc31a3822d709843f3395c365528473e66ea05421526dd9160cce6fd11df8779b14d9f63b89a9e41aec7fd1869af9b97bb625678ec97f641b09832b0881c55bba055b50a3830cc530c886e33bc354498173deb82094b5ea6cb08a27cc348b944d21724b61a3f3d486b7721ed08be9327671ef44249cb3cf2ca7da1;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h3cc3b8409fe56eb88ae661b83e7bda17d7dc91dc078308cc91afbe747480bb70a0686ce3c265cd3108efc6ac900357ed982947b937cc2e5afc3189ea831564d79b53936bb1a80e23c2c2676603b3a0e61480de43b570a6229a804a6bbee486f90ba50ebe1492002f64f207c500338a26c5c3d7d75333407549eebccedf4b0b20bbe9d4a36a30fa10f4bcda84bd273571f3075dc474fdf1d49ecaa97166eda3f6b614abefd1d4f6dd887cc4385b6b276cff66b51b00d97f55e873e2c907b1a444cb67100ad851142c078c6cf01d90e396859e7746fe91ee206bf23999eb459dc2dc1f63d6641ea9d9786dd78b358f4561b5956f515a51e64bfd5c64d7ea87950;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h2a453a942052eae99f3fad20e9daf83bfb6d518faab26615c4771a7296ceb2c946e52ff2777f9d5b50b8b05bbf193a4474511182e804143f28ef4c0a2a7022c8543d80ffad85179cc73d5dfa39b909b4c215cb7d526e846906cac9c6648f819afd8ab9be3ae4a434fe45faa46c5a77eb72ed1cba7e2646484f4f6daf63f5bf00c4017d06897cfa9eb858012d367798ddd82bfaed9b78d97880433ba6a19931a0c513ae442883a190a1fe53c3a53c2581a0b05904969492c56a9fd9a2169078b7167100bb7278069772728d422ca73d02367e0a22ae0d3e04a1f82b65167b8bdf156fb70957081a4bde719e502f12b33b82876f213373676933ee17761717b791;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h948a0bff3ecb3692f28ac5b7c2ec369e4d9d49eee8760b2b309207afead37625c47a5f5b8bafe5fd3d052617cc6b0e13deb36f935ed454cef2718b34f4ea2967f15a2bc4d6f88b5f6c67cbbfebc97c6eef7a79954cfe4832d9d5ec98ff27ae7b953e8e51e08bcf59a830c82d3f32ec0327210bdd70e17cdf799a28c94b6ea166fa414c649d9de63d9f9e7dd0b66b2a200fde22eaeec2b9a00f81126d925afa1b667f01655e64a1f05afc623b4783b77febe53276200dee69bb0e5a03b1e3493ce7cca0957b4392ac3e031352b3c186d418d2dfd4a499f66b542b30bfcef9ee7a0f4a6213aea854bfc516eac5e7b5ddb2495af89ce12844857f5ed6ade0e1a7f8;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h36fefabbefc7589c19825cffb2a3bebb19367182bd149e0980ecad160a82f24dd8be3ec84c95ce1a53c8eee1cd1cbe7d9d3f314aa5fc0daecd09e33fd10592685b32c451c66112df8483e24e6c179ec35bd953989f444586dfaebf28263e5fef21d2a8de64976f04bb95a8ddef7a63614c38c3e3cdb128233dd1927aa5a968938c6b97be8b060ba547852e34f096691ca288efec543aa96a16ba90c80e41a6148f17c433cfc73ac6e58c1281f434abf055ca0e3d57691e1870de03b0efa95c8ba4eb693d3bacde175b07f5c294758bd1f67d5a9dddd8afb5acb75ea2df0af097cd665d071bf5b04a8dd6048e2bbe812af0dcdeb4723ff8dabfb7327d28f2ebf0;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h1ab8dae8c9bbf2b6ff24102d7e3c88f4f6bb6c5a5d21226cc513f1da063805e9f670806eeb0da6d5a012907a7413c9eeb87c2dff3a43035013ad8feb632c65ff68f54f902fa0c867f2138be3603f0f4cd45f9cfd469b1741bcedf81ace342f3eef1a9b972a1b5c263796e88d653e98b0af5392cb5cfefbcea98b6d3df2387ff5587c63cb39026d6e455a2753eb3587e1b77101e7078bfd1c88bff27362a3dbc89ee183938f7575439e9fbd52b87d860f3bec4b5373e78c96416961f5eb7ce961d6d419a010df73f839ecbb627471e1feffa51ba47b60dbbb6f62bcbb82208221097cd2ab1a39308072e7f51abb8b32778e31dc5031052b0eed7fcbb76d8d5372;
        #1
        {src63, src62, src61, src60, src59, src58, src57, src56, src55, src54, src53, src52, src51, src50, src49, src48, src47, src46, src45, src44, src43, src42, src41, src40, src39, src38, src37, src36, src35, src34, src33, src32, src31, src30, src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 2048'h77e843a5687602e04d47b3b996917a60748fc53f0e438ce92834e0fbefbb92b1001f88d07ad64d1e9cd330dcf3a67791dc180a0c5541232f06513b076642051d00107e10d4ba61e74c495319cd205b7ed80081aadaa2238ea946f9e810a5d007f7c3d41cb9ae411f5d91cebf8525f3be48852e0ed288f09301d5cac5e1076ec8cf7991f267ef2c794760b7993359a81eab883ca1da41e10577e23e14af6fd2fe8071b02eb5c5e1b5a41efe436994278e86b1754e79f9a2c09f2b446fe851e284a40b78de35f54b6362d22de178acf979de4532ac54b2c23a61f304dd11ea8fa60eddb8458da7ed883941d608557eb92a17f7fe970882372e1d5c5aa8dd6db118;
        #1
        $finish();
    end
endmodule
