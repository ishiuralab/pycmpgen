module testbench();
    reg [8:0] src0;
    reg [8:0] src1;
    reg [8:0] src2;
    reg [8:0] src3;
    reg [8:0] src4;
    reg [8:0] src5;
    reg [8:0] src6;
    reg [8:0] src7;
    reg [8:0] src8;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [12:0] srcsum;
    wire [12:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8])<<8);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ffffffffffffffffffff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19f21385539b7112503be;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hadcc6ce7dc4541a2917c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h167c6ede0b578e2fd7dd7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd66d7b013dd83e281ada;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h98b6053023d68855fbda;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb60eca14ca6b23f2d83d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha54213863267a756fe0d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h208d62ae0d1eae94e4c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18858707c8c4160a9d33e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf1dc2582baac5aebf8c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14f338ec21818f6f52c98;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h150c3670331abec7aa9c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9fd60e41bff909ba83f8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h187d6e06dee919263413f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha73914d474b6b7c8312d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h98fbbd970f43bac3496a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcee7f42fbda2f936685c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d895e37c414356c647a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h151d5a8d3d75995095664;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd2448d9f1cab307c05ad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15189c61dc4df9919708b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h39db23b4a7e9a1a4321f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbc2430a9ab8804be86f2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4bdfc0f335251ce098f4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf96e695c72f9999f6b20;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15d9a8bab84df11f036d4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he1b5fa3ea2c50f2e6304;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc4d1ae9aec4ac41c1b7c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11db3a421db82a4274378;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17a125ef88c616db4f220;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h62e7fcceaa5cf6d71958;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11586cec90d5786268be8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c39f9d81d9835a679e78;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4775487ff9899ad9e4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15a4298be3b5ac7912e01;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h94279a8599052531a58e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15ab4c6fdab571f5348a9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a3ace7caefc2e21b3298;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d7837b8dbdc7b458b23;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5abd3499d4c3b2f06498;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h908af521a11324cf2a89;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4a340e92544a5e534cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9b0fd03018196530fdaf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha3dc06fd502f4e01a26e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cb28b35dfc1ec8045345;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cac22b853b689119d8e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h82bda40b8d813c6b0358;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18469821b61ed4388f377;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h190e1ff8cec2a299bf141;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha408abbbe6a5751e94f5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11603cb2b2c5757f673d0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf94cf7b332d1cb819afe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcb83e53f379e5c0d2b55;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ba836fbe438a759e4a6f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he459da4c268c2c189525;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1de410b135b64db334e28;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b1a74a64dc32cee52094;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7505e57c0a40df725659;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h751d089816ed8581d6fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb058f0eb75e9c242afa5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1780ae8f53e438e5d2466;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc99ac195ee81ee37df92;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10c6d139fa2d60d564218;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1baaad6eb5e32d451c3c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h21256fafc398e2f59d67;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h27854da78fa302952ab5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12cc026cb43b00967c39b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf8dfa7abd51b5eea59;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1600ff45960e1fdec42bc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h148f394556ccc355a71a2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h53816177f60484b4b9c7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1098bcbc54165ec72ff0b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h151faea84e09d716ec560;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb9519fb776aa3aff3db5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dbf4e79ce8a72f0d6a85;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h78db62f6d1187c6464a3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fa9fa3bd375c3bf4d9e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cb26dede1bbcd0f35fe6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h58034781aea9a455ef04;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcff8635a3971f380fec1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h451dab66495fbd05274d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h89331db1f4d6b616b44f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e1b1db63d9ebfd6dfb7f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12afba072105f978f2ebd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h100c4856005381c7ad4fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e3b5959cad02663f1edd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d09d1cecd13895367625;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e53b4f9fbb2372504a1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h640dc2df746193fb91ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5eacd4d5a52b1272a7f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12b47f8fb2d24d62cc107;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12c522459aa8f38462f69;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8896e58f824fca4b176;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17d6d1cb4d187933b6ff4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h906a342631e34066dea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbdfdf9e022f2d40faf59;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18ab6cc9c4916386f9a27;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1750591f242c303919a87;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e97ad966a34954edd49a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a6f6bc2bc19a6f7731ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d9e4cdb941622c2ef88c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h204b0867b658d5fac49a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h563a387c31a0c4174b4d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf76f3fbfd3fd7dbb79d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c87ee525b3382358e95;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h143062879203b9444fa8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1361a2eb6aeb55e89c4ab;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1efde587d29997d1a6fda;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eba6d1e1dfedae20a78f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a72221ea5ce118f3f91a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf84489fb9129395cfa4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a1d9d9d0e05448ed36d7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10b646709e624527f7316;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19e5880f82a891af2dcb8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b996eebd7fab0a667fac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1baf6f014fe07be5ce2bd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14329f338563195ea9a84;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9ecb3dd1b574693d2caa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18b4bfff45b6fcb0fd4be;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c7af2ebe4fce2e9913d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfe13986259aa563be529;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15b73dd2a67ce8f3b12d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d124788b88fb7720720d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16b843d912f883ca0d38d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h94c919f65d3844b8ff43;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h64ca69faeeabd914f636;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha12aa03b873fecf38cd2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h161bf05207161ca1f5707;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9c21383386b111832660;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7f590dd3a8311ed3e7fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hba134e3b39221630406;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12c0c7baec62d05de079d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb1cc79011f535ce38a52;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h81fe9dc8a6b83ce0cbe6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eadee7974760062a2e05;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h102af5e0bb69c6dc69629;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h89360c78d3484ba65a00;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11b50111bce49bae02ea1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e33b01692cf9ddd8dacd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e0b027be62cb5cb4eb47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19a4e8c1bf6aea82ace49;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf2126260abc10fa74fec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h25bac1b897787bdb8264;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcbf763f416f59411eb60;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f20aa4b74aa0895d71ba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f33810dfbc10dc2bd1e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hef8d2dc37dc1ab70bd8b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b332762b36afa0701d94;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a69147835cf948ef116e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h272f99c94e535844a2c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ab476b2870d67dfaaaf2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h52e0b22f3af27c01d06;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h42503831f7cd839db5a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h36644ae6c1801dffef2d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ce464199fbea2c7991f3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he78dfdc59084c522e00d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4132157278e636b3977a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eb55e10030254c39d53d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h241ef4a154e9351513e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ddc4c387b1fff5f49f2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he546b9ce6ffc1f4b65f4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h102ad3b6fdf5041c5deae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h136b5fb39538cd279e534;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h31cc57a2a6d3d991c198;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14a2af47e35243e256636;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ea5407a7f7c1417d1aa2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h56208cf4326110f30e0c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f6248898716b08c2693;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bcfdd67800e6a8436deb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc70b4b86dc62d8df51f2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1907b8438dd61027b838c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h658e58ccb3a00d277b58;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h72d11ed5f92d7a5b522f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1076e8f1ada6dd32edf6a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h605abdb411c5c4598c76;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ecb5ae856a7667611dd4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h60fce713bcae7d370d50;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e2da7c63f72924775a0a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb9dbf84980f9ac7da8b2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h187fdbce7d666a03d2106;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e2d3c334d6bb79d3a025;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf4fd6afe2ba16d9c93cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6e50c9c9db0eb0998e59;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1aab0c970a31971be398b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc862cfd5f80e26b13d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h184ac79920e1d67604290;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ad8557ddd1f9a12b1334;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10c03606f55f52bc8c5c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1596b6bf494ad4fa05eeb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h41c075680e3b959952f3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a59403421ed3af7ba0c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b3df5817689a7d5da0c7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ba800b5d9302505275f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h143f81f36b861c57e53b1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6eb2376577eed841049f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1af1b2d1847d3326c4849;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11fd88af92f23c5f4beeb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10f815151b022dcecb455;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2f67ef70c10a69e79262;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h100c1590af9b43ab54d1f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ea2dffc7ff2f3dc17be8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd6ca9bfd554a78b5e0a0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11281ede915741969c458;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5249dc0107010fc3e62;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h92b79fdc4d8b86d381db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h178de81ccc9c7a996c08;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1121c34fbffe6400f34d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c678cce659bf0331c8b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f9ce8682e05da805ecf5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1929e3793948b2e2e7c1b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13f27c999c4b60d7966fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc5542da253bd2393d3c1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc5c4e8ce651409737f25;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hde331fd8b84411ded824;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he6972279e0abba5120f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14fd85302544d0dbc2bc8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h59e7148d38389806db81;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd97987aa36ac96e34bb3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19af7c82c900f4d458672;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12040a492b9b39b8e79c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1517e796a2aab4d91540;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1148a905909732d860084;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2aa771183e155bd67e55;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha929fcd5ef69f5ed33ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c21a375261e6c548fd44;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1495a15b2ced53873ebef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h332dc2a1ff2b2b314a5e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f617d08ef3db70e56fe0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14963518564d0fdd064b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h83e90351e9ac0ad9910f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h95af33849025e88c9c6e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2665cce3b175f0456eec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h73f02f150f9073917526;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19f6bf3d9fd2f4a87b0cb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f036584f9796f0cbe0b6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h137c51e4826c11dfdc200;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1db52ee0ba2f229fc659d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h186cb27c25000328f26c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h22b451da9195f64858b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5a8b595869de7804a899;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3a3b77cbca34b21ef8c7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h39d3719658fff714a456;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h199876b47771dea373c31;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf03d7707baf404476950;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h150706dea6a592a1e3d61;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc32dfbdc94efe0b5bb46;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h375db283550dc718bd23;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h86b88c771b30a4776031;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1187810b0c73332954dbe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h51b48cd20506ce3902ae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcca4ccf432e404130249;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h177a3e9a3e8ffaada82a4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha0119e339ef54c89d01;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h130ae891df8c041be53a2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bdda6947218c03f2191f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fb4303fe6e4cb5a4d72b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd10bdb3ae0394c421c3f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d2b4d645a0affd78960;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f18c2a73b11a230726a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b39e0f773bb5fd92d442;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h31759454b376dcc938fa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h100fb68cc94ee2aa0d159;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1192f86a11acdc156eabd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6b62c6b75132a06b5b18;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8eb3ce7945be5714fdec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4747165a83d4b9eb2716;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f2fd19d2f5d2d430f4af;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha688f26529f9f9d583e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c92627249757c115a475;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h57e0b85a1932b3623508;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1079f29595a782bf5864f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10c8aa4a82ea0848a32ad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha82a17f972470d30743c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1babc2a90237f6959a5b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h908ba916ccb946f18bb1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hda3e2595b9a4583cec7e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'habae508053b7c9e56ac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b2d2a56f23bebd551b2f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h197437ea6a322ea4c0b79;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h127096bb1c956c3e0f976;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haa51ffab480f58c7ef54;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18f06eee979c66c0a5b4d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19e67a2572842d681d2c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he90aea0ad66a98602af9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h142072aa124712f48a3f1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13a080ce5a316fcdb7e2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12036cadf5c7a56acf19c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8d123b132fadb6c890e3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdfa1aecf21a3b5fbeea0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he399fcd38b20ff15d394;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h68b197543cb00bdac9d5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bc7a921437aac22d4ec4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h847e80220745d2149375;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4d2c8f426b45bdd38846;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h932be76bbb919c199340;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h455a9a86588ef3eec708;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bda390c8301697dc987d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hddff5ee09aa5dc26b704;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c36d59b1611d98c9915;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h171ac09e15bea69886a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16e3dcf7aaa3c7e4480c9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10b838098eb3c6886fbc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h144b19a6d3dae7279084c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1722ac49c893c4fb1869b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h141681224be22eadd6945;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1556b0e2035cf6cdcc8f2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d753fccc3b65a509c7ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h120cafd6a0f3044acfe5a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ed4be68fff99aeb5098;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h104e13ad043fada82c7d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf0786b980ca047c5036e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12ab5f073ddd8e22f1ad7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd0d406205dd8f67e0fbb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16f2bb822daa4407fe0b7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h29b2ef690b0ec79b17d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h256088ebbe9ee88b703;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd96fb8fe23298e9e75e2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12ca8ef6ec6d903680fa7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h901e79264d95f3fc567;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e20f3f68a6734e582a43;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16012683b761066c9ab85;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ad5f338168360bf7589f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1236e2b0b6c0e45032377;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18572c0a56c8bb8128d7a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bb62800ac934b2baaff1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h307bb0e965f615480b86;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a33af9a4df1b52b15437;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2d82db8b0d24ba301633;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h62d064ff5c95ab973cdc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h156292d3d4176b08c912;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf778c0d5079414eb49e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1727de22c2175303e6750;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h143e43f9e72e16ad4fa9c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7a23b6a9c0220b2f505;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13d7c23a5ec978aa9421a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2dd981eaeb7ee3913491;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd4adc8200737925de4d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6260de42ef941fb1928c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19e18a9e7037632af07d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb3e28ce37512487dd58b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b24c8c295cb474bca5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18cdf9e4f069edcf5de3b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha96c35f9b4f8d69c5c88;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h41c66691c7ebf72128c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb9c54bc74036793dfeac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fd8ea7653d26be6caaad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19275430f1bc06e211fbb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h116d2f06466b09017ed73;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5fa41ce59b61180c5359;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2f1efd14e6698c830b4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e8bb9f8d9a22df8c6de;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h54df1dcb05b0bb09f1b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he9d24713990996bb12ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e6e5f1057dd0d39edb55;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfdabb85677b33166d478;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17216d4ce5c24e61aaf06;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ee1ee949248c8f3af34b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f70d2664588cfe4f07bc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c8a73b460062e29714ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h131132c65d1cdf6bcc4f8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12e059f37a5f77a7a3fb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cc92c5b3baba7d009ac4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h964bc20b73c7633e3f35;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hab547ae48c3897ebdaef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h124cc0ef4832392bb7d7d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13f471f353003b7ad1bb0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f9325836ac1e93ba0cc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h58695a8a5ef8d8b93ae3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14910ea566916a7c969c7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a886b140ca58d24aeb1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b3ebcee17ec714ccfedd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h104e18ad2ed1a4f42915b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h100c74af0b5e1e6e374e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h67cd2c8d3625f43383e1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b831ded35495ebec4655;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfefb44b215fadabb8d48;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10f2fe5da9793c59df88f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h89f2da2b90e9ecd4ee43;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h42d59f0443504251c1f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e4d1fd80155df654a296;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f62c9a52d3054c06ae11;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf7a424fcf080d8a9a373;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10805783cc573a272e581;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a1ce1e8356c89b85cfcc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1da24f7db8fc790f071ad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e4f8b6c6ead9cc2ff5df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19922c17a8faad9399bda;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h165cf5cd581f4ed00835b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h185733716312984faf3fd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hda413ff0a958ffe0607d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h72fa211e372fd6bcac2a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a537ff28cbc7d7444985;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h174fc4bc1725bdf9d8f1f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h782df1e6b32f6b84413d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb0c56a4452f4c9d384a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf0e513d7086c5015247;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18024d94ac9faa613de30;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b56fc520b87e2d19d467;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h139bdd234200580c1c153;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15cb76ff31a37fa527e76;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2a42abae6e55f3e3368c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d0e4fdb5404aee066d44;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4e12688c996d01fdf6d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17822e9141d72b0acb319;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e99f80fd45c1201b6eaa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bc8690d3b1a879682b77;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4514709d6593ec72927e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8ad225c16fa78175461c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he86e61ba8f432674728c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9ffa1686f019a8aa09d9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ebd37f9570caa7d11c46;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1523b43f9dd780107ba5c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bba605d4cfdebe100dc4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ffc67c6a5451603f3f8e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19431bf3fdbc8a5b1733b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eef4563a10a7a50db5c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hce89e133f03ce631c411;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11c2c9ffbcf2ed9b07278;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12253c1fd9628a230a33a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h88b24a6bbd450aef1320;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd4d38ebb2ae3ea6ac55b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8562ca62da1c0f0ea6a3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19f0c3223d776f1bcff06;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19849602aa1e1a914c72d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h85ab619083378ecf55fd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf35aefc833e86c30e317;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ed3cf5a1b6c50f7e482e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15125574740656f438a4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f5a1b23e6d051db5da24;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h115a36ccf398cd23315a1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4dcbda0237ef7648d762;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5a2ef6a9f9fad2a01754;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a0e694f47d8ed5a1059b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h106a650a08b94a9fa2e47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h851bfbcab52028ed51be;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h100c5ae34666f48bffe80;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cc6873bb9dccb039c25a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb62b254f09e5418e5094;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12cd289d7e6fd7bfedc94;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e48d7ed9c95c8ce04304;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he6d00d75862190837fad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d66d16efbfc437c8f54c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1724041c8bd9d77b5e2d4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ccd9560ab006565d0348;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h76965b411c5cc50bf3ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ac192ff392c58c788f1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3bcf520a36b08b4083cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h87428382bc39f197e922;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9cda6f10f916ce23ad61;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h79fb4d0ceb825e0a303a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d8e9d5f8c68e3019aacb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h100366ed813f506f4f81e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haf8aa999bc9e757a5a81;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd080d7f8f258e66e14aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha16fee5ab02aaae0dca8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbc810d3c8e1a91fe6ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9b21dc22d1f645ef60ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha26e1b95a8be52c8a184;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1da9e70294aa444abd7e8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2739a9b79dbe65b7a0e9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6f126b926df783449c22;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h167462cd346aa3ab458f6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4454e7a73bf51b29c33e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ddfcf7d875fc39ef680;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1469eb1ff5063bdbc9555;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h183ef550d9e4b6b7b50cd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b2bc35f4587400248c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11ff6cd9cd939614881b4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13ee7ec8611c750d72b01;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he9b897cee788d7c91e7d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1401d527df7548ed4ebb2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3b49eb65c7e4ae4bcec0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h87a154add7385d6433d5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16c477572146f8a402492;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd6316feb4c5b4d9708fe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7faa3d3928a0c8cd7896;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he3a5062dac86ba4bf232;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h105db02bd7eb9ffcaafd8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e1e53390e1af5ffbeb67;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd67236325ef5b6aece76;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16b6edfa34cad4d7da330;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb57b7aaf24ea5920580d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h94e36202de95dbebf7d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h142fe7955a78e39d622f9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19b3ce186b91ad4e1a975;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7366ccec57d71dc11516;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3321e4a4b7847a588571;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h748e7152b9a9f3ade391;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2df7777b312b62f7adf5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18757c9bb2c26834d0a3e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5fd9d35d7199e5c0158c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a04f31a5bd42bd27b5eb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14b6c21b180812425a9f8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb3c6b1e4465d296814e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd836b479592e73b8e5f2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha8b674610bd31d62edf8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d83f6388826b02387680;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c6c572e241ac790898ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10bc409b4582cbfb47a3f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18ebdfad566ac95ce9e90;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16511ad73dee45c0c55;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17e8e2239a90fae4076c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a14c3d63541bc989f01e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc19ad9e8f1e7472f6f57;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10a065ae93b1652c6ba0f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d71005d888bf691af574;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1757d79becd24e19d8224;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b194d5fadf7e25bf8e64;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfb4e8abafa29149656ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h162bc563e7312e5d53471;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e985dcb3f77a0e6db9f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ae4377bb39cf0486f6b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1631e3ef85137c6d74046;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb3c5633e0600fa442adf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c00f5dee099e6e2ad12c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4f157d7359dac1750506;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h207247a5f0b7ca7318b9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h194fb704db535550d4624;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18608181a6fbd3c8ab568;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b6efc01b4af6d1dc621d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1588d1b609131f4a14051;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c6f7147c8d3b0f97ea5d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14269f8fedbd6d3e6573e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h409b4af44e029a790e46;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b2181e144d681c93da49;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1837e07f7a9efe8865e75;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha5129c9138775dc75f32;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c774e03d94031d33bfd3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16b8254e0b2e0e96b3bd6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14c7add6a5c6b210c69ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15d0e46c600699e488e22;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17d570a20156971822435;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h62645185640aec8ac5eb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hee6c8d14a208547703ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hed018bdbed612b9a3e14;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h52fae46b10d626e32ece;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e7995af2036eb65c7ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3809ca83497a571783b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb86e055da727322920f4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h199ca4e5b28a42f838caa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8560cb82babd00f7da53;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h89afbab7fdd528f5b72;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h198b341f63ad28ade767a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1341c5b3675bbde8f9e7a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf4ab008be014a6c50902;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1411552ac4ada69dd0b78;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he9cb7fb06830b5d61480;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e37e4c5415df4867f38f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1638679c5eabfec28f3b1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5b372efd1b7d1d6c2069;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcc0dc23b6193b41586f9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c17ccb2b2080e1f45b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9341085523dbe871a6f5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16ae519bfe42b152ee646;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10e2cd805471b9561b1d8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4e5efa79cabb91e43fa2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfe2a9d3a7de38023299;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a32cee96aed1d1d3f7c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1351761b1a1804e2ffb05;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h98cfda12aa2f254988f3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c2bd0ffe1caaeff09889;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13adc344544750697f275;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h30307162ae28d9f8085b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he91761789d5ec4620e32;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h123cefb2dbeb15306e800;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6a2d5b9c94cfa3007eb5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1644844c777fd448faedb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h20b69571e6b4520921de;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc78e10ad5ef59a5b0038;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10f7210193b2653e13e19;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd3313bfac446dbdcbb35;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbbfb96e595ba4c494070;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c47fde09a692b1ec70e6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd60b593b021fc4d3340b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h36c6696537ec67b4537f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f6765764ec26ab80e42a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc031c39b8f30dfbd3c80;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h184a66dd645971f639533;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ed3e819843176b68e62;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15a42bc24ce9de89c9eb9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16aad732651d7d395f4ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1275ea1c1ea3c36961162;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfac9d1630cbeffe11204;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1349105ca651f4f7ad4a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a06aaa2a792e5a698b65;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h174ed91c1ec1fc141297b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6ce0dc95c9e89fec8c25;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19d64f0d19409d8d92b27;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b5ef5eb0a9fed8e4a935;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbfb2f7b03567e5251c98;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10608ae0b6caa892d6dc8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he0f28e669e319050062a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfcc2d0f6b07b0a3dcfd3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dabea971b2e8cf891f37;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d252ca9f05b564314bbd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h146c39d96dfa783466674;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd7ec2b7777530802961e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d0dc3981a39169efe879;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ef46c46a41e8cbc9ff76;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16395931ed0fb5edd3f20;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ca0ed97a8513c0c53da4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c842d5e15ee353d4dcfb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha12b6bf8cd9aabb40409;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h141f17ee7fad65590bb3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h163c85ff99ce61c450ec7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3cb580e1610ae5f5a467;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18fb400063cba5967c974;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heee7de8e9b67d07593ef;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he70fb78c83cefd3cdb8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h841fb8be08498985e9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ef663162e5f7fcfb60ec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bf3f8587f16dfde221cd;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd77bccbdb5e4a5d992f9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8600c4dae7249a9fb87a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e5188e4757fe1008d633;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18f504be7f557ccae3772;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he5173c4bd31b552179a0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15198799ab029bbf4416f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h135adcf781ad9a72e1b7a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfdf3e0ab646a92c16b4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c6d4c5c99818fe931377;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11a5d8407bfa2fb2df438;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h411d8330ece779880548;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e1e9b5fd3c48a7872c1b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12e1f3da7db094fd30ea3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h150c4a94b3aa1f19f2b69;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c0f47779c3006289f093;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdc0e41082b139962ff3d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c793440a43942e8668d7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcee1615e5cb165381557;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5ee99af101d5f9090093;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ca672218d2855187c40c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15f3e6284ae0597397c98;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'habed8f0a811f4d16f2b1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h197b31e853ff3b71eba66;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5392e42aff60a0cdfcd8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd4d7d13f473fffee9066;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5abd21a30e4940bfc7f1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h152e7d2f73fa3a33f802c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e259d53599440b1ee6d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h62ecb09d2677027f25d1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17e15e0b20f93902162db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e6054ae982026b791c07;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17f7053fb96f5a2db4ba6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c4e10311e089de0aa7a9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5a40842ebdc2b019af61;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h140981f93a2bf491c1e23;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h166d12cf3e9004301c0e3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h192b1e6df9740960d5ed3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12b7f6d8ed37b2f8d77ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a1200ca02b7cd211db68;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d59de0d36b4f498871df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h379011707aaf8373b346;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h131ede13848d79fa0a107;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc0eb71ea86897aab18c2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h101f5f287dfd39ea76ee1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hda7dbd9b0ebb05f5ddf3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9ed3d216b4292664bc59;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h155660a70721ad07f294b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h196bf67dd443a0654a918;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd3a28b5b4718f4339228;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdecaef730ecc89b43529;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10356c367d7efc6bc489d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ff2de77e7d88ca8faac1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4eb523bbba495d55847a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h192b6dcad11a6b3c25db9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ac1915fcf8444996534e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h98e5933ee76645259520;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16bf6dde6defa7708fc74;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc440c356b9b64d920212;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h103687e6fd887035befe8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h443dee081048aa8579d3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfdc47cea67fd9b76c55d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6a8da7ab9cae3f186e1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h101add41fc7adfb742071;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3794a1dc828d2e56bdd9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h660ff62ca2606a723b8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h101adc03686eb3030cbc8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1823833eb41212a8d148e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h952d2ee407d64932945a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a2f2ff0e4558eae83185;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a65cd7791548dd491060;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hec801c140e173920990e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb1ea89d1317f1165d40e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h623181c1184cf055422;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f30f039569e3c61ba8c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h110ede90ad5428a1dc38c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a4980c8f80d9d95d4809;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b34103dd45b02fee06c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17b4cede0e3f718ba158a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h80258442d948ac1bce04;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha9e72f3d55a44870d71d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fde11d9f7bf52bf798aa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12f6aa66173e07bdddf83;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h587767e7973727d675e7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h126a121e6fe21150db16a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1022edbc290cf77afb490;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdf934a0b54890c36217b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb376ec7c2099fc23fdf3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h958df3723124a6637845;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha8c6391e822ebe9d7181;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2d8f3a79ec370f66a80e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1807bb8360c48c2922d06;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ceeca538bb23bcb42155;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e0132c3c0e1241029cf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1acbb228c40cb4a7eb357;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hae3a006c6e43a0194ddc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha467caf1ec6c35c853ad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb4fa2eee7c3eb944f7c3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'habe215a3b946f586f1c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12b9913ff7f32db3f5fdb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h143d6384d8b8b4e90dbfc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f0ce127a7c5718afc1ad;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7efc4653c25b4834b338;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdc6e7e1cc9c4fb931c0f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h630c8d1a7a58313a6573;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d789c2a3a86623187b27;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcfe015bfd3ab21e2055a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h126e318c767a52d5b10ce;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dacbc432b6d68ddc0398;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha0390f24f9b0a6cce3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haf04531eebe005ec21e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1484c8eed22633b496214;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hccfe36d9a1f2464aaead;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1eefc59001e8e106f5087;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc5baaf4ca5e412b80ee;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c20c3ac0001c53e452ec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfc0559250daa5200bfca;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb7cef0a84f34a259e4b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h127f92f2159b79bf65b8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h751681f8e0d3dc956cc3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2741579c9e287adc151f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h28b403dbf3ac5f2d94f5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f7388705ed6ded12c752;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bbbe28b47b471073ef8c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fc15634209d5aabf235;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17aa7ede3a3163579077f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19a5117185ea3f321417a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e6834984ee5dd86ff67;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hedaf428972ccbcc361bc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb6841350fb7792afb81b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h103daf03042f6eeb525b6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19efbb1df19cf738a68b8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7a198352a16e096c8a2e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14c587db11a516e100bd1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c64c075a932c5b6a18b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14598afeb8084f0a10b6b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a942841a61b12cc87707;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15691f5a99bd04a730824;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h143fe36f67446c317c2eb;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h149ebfc4b2850043eff7e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h173e3d98a122aa0f95c58;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bbf530d4f480043a61b6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19acb9a69b47d3772d13;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ac09fb94f0281d905345;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10f73b73f4cbd1d087cbf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1267d784ed1756243906c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d94139fb235e48f039fa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h127774cbf34b743eef25d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3b9c404a1d5c819e8cc7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18003614d5b6d6d03f710;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16938c1323c689f55cd84;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b81b755317c043dac6f0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he0dcf621d7389cb004a8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1db5079e919062021b6d6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2b31242e8e0b067919d2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1091b9280b7e8515351c0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h120299dac6ce8cc40c072;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13346ff4837537be8af2e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1442616cff1a7aa0acfba;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h161fe997cb0e28730cb9d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c2b58e47c5d6897aba0c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h68ae4eabae2f91b3239e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h73724d468b1608fee996;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16826478500ef389678e3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha02e6e673f82c7c2114b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h752fe35e5f76c424565c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4dab5e166e8441f87b3a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbac1db31ff693aa87d1f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bc2cbc61678f9c2af187;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b08c843b27e01ee1e6e3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfd608d6666e4aeb37b45;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12a283786f8ee6d18fa57;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h48e2ff6ed06c56a619c6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3789ff3d051921fbb5a1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h58bc8e8ee13b745d2fe7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9dcee410a49762f798f5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14a073eef9bd4f3fa776b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbc481a2ab4b9f8e6b9f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h28644feefd54b4362126;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb505e8d7bc811f37a487;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13ec59b736db709d8a55d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'haf6af0b4470b6de01284;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h119fc133ea7840ae5ba45;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e71fb4f228e3b94420df;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbb57bc820e0241477f75;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19040d7ea8792c87b392f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb4ac9b34dfca99b16369;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c1e0e17504e37b643287;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ca278873396b1a9dadfa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4b805d2f6c333d2c1da2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19e356541f72aaad94b11;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h140c94670926076898207;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h31974004f09ecb8bac4b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h146e7541423b624052c5b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16248da5ac57c4f06eaec;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3beb43c39a155b1a9dc1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10a7cd3cc26b1291f08ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h27c5121971d9acae6a2a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h57c6231cbd9da5be2b6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he0467cc23384755cfe26;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8b7cb1c7f7d62a32d59b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1296f4b0b604bac29af82;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'heb64725ad3de647c0216;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha4daf2f95937fd482800;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h182d11c36280dba2eabb5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h124d04c9a61989feb0d72;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf5e5327dbe12bcd7e122;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha77467b7ad44298b885e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f17db005c06897190b53;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h146eecba0becddc3b11a1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hfb0339fe0d6cba078eae;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14a0913227615c91b4fed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf895eebe2e5d486d59f8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb5f8a7c4522adc93e86c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he212dc9bebc19562a7c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4540f2fe9eaee88a5ace;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h189851b71d91c91f4c89d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10261cd0885e6d089b31a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h84f7ad516e98f8891244;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11f10c7248442c3b1e178;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9d0f4d2ea7d777e2ce72;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h52839bc942de9be15ac9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a70b22d50ee0ad3a4cfe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14b7a5905a379b5424d47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb05d4ff9130d7a445157;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h9f558f63f6b1dc50bf5b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ee67b52b0fc24ec96b5f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15d4494761bdd7a7eac51;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f721c7b9104b11089aa6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c806836310cb23cde950;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11f9351c01a191bf937e9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15b40522761c6854df82d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha2779ac1b785dd58cb3c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ee99f3cfed1be327c37f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19eadc621e0d6bbe06c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f4c16e91d9611a8c7231;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h50cef55a3c1d31e3a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13a988ae165e3cbdc8b4f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c2eb77213f8e154f148e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4b7bdd5755435a90ceac;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1299444646d1cf0c32bde;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ab56238d1bc0ffbd35a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8843abba17ab94d6e1dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c1425d310586c7adba8f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11e02cbe2ab9b222d5331;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ed4bf26be3dba10ae272;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3a6e09f94a829e5a657;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h913ad71036639601b588;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fe09285c060f1120958;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19630c2abae4d841889c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a9b2f624c1d0ba7f588f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1208a744e4f032426f014;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15df1882d41f917d01bf1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a20a1a8f89f72e0d151d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a7c393fdc814ab5cd99;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h140749d599661d841167;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18ed605ef8ad0ec2a9b4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1145550121ba948bb9a7c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b3f9d16f50f1532c4f46;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7d1beca618456a61099d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb592e299a8b8fb38abc5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h359ff420cb910bc71cff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h74e85d4589344a0f585;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d8a82ed22a82dd6e7f78;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h102e8c00eb672330d2346;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h27a461ad53c18afee77;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2d5d8407b55808b4f8c1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13618b51e99f7bde94b74;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h657b9b95a9464477e84d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h164ee018317d387ed499;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8ebc679b0b072a96e623;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17001e41a3e48e660e224;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d37e8e09149af2e9b33;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f39c1d34942286032b88;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h73451df3c9a9f5de6bc2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12853e818608318946a0e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hadb6aa900e74e31076b1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h229ac239ac05090bd838;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he213a6aed74ab0cd15ff;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1824af99bb93a47f3f5fe;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8da07babf1ab88a82a80;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17e44b971b8d17c952a59;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14063be7fd820c386133;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h77c30968fb11c5d909a2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e000be7a821923932389;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h333e689e234600ce0b16;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8248860c528a2240762a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbbf8e408ab0a1d9834db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16474b10c05a19aaa62db;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8b31715b33aa21775468;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15327ee193e4692f8c30b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h127f6db7965b4230c511f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h75755009f60e5e1815ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f04bf863d9de41d40c32;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1bbd4b4ed5fba634b9e8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd913654afaa497f3daf7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1affa4987fbdbc0729e33;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10fc772b8da4808c6e7a0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h18c026a117673436879c4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14a0caa49d34270412e47;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h422c94d1e320f5650b4c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13249ee0695e46c46d80d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c1f9d6053ca28a367a3c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ad0a171c150da1cf275;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16cfd8205d4d94f237942;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b5d31817e4ee9f43b255;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h31b7533b75f7b92e1253;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h883924351defca64cbe8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1ce93910aaec36aeea9b1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h147aa571568c209734871;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5ef4fa79b93789269928;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11cc645722681075991b9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15c88ee76e92e444d80a0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf120e8a5040d813c4d65;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h172abd300b604f387ff8e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1152ae88486b1c4a0d918;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h149d666a66f4be12b973a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha0fc9dfe07be1fe5f859;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16d8304d3bda05269cf2b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h298e900b5122baa3003b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdd5ffa94982be005a8dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h105a6423e5ed7f36aacb7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h25a989ffc617e6cf3ff2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha70953dbfba7e08ba6ea;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h34a176f135c90425a4dc;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h227e7fe0903e3dae0597;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1718eb00f8494f8a79e89;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19146b466fbc0936cca40;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hef7abdf6c02cf2cbc645;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1a6ea7174e327e3c1f1a1;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hd911a4c65feef7c32235;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3ac217d4a539bc65a30e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdcbe5e292053caada1b0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hea1e4d721a53c4ae0de4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h496890e3da96b697517d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc306b3064e99029bddaa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1b0b8b9ae31432ce0f108;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d4e8dd17d2c30db35a22;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h176cd7985876bfe5a799d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19aa4de66dab13934a3ed;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h10eb7e95111b05d451789;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h97769bff91a6daf63186;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17c010c5bd78b3a6c6490;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf02a640890b9764cbe8d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5700b2e778c9c2c1edb5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h14de69c8d2c68e6abb4e5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fe918ef4ddb0626e312f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3aaff8d600bf677540bf;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1213146a8475523d6df91;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c35fe7dd6f927396775c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcaf9ad3a5770a640ac9b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d855210b0cfaaa66521b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1f3289f397f80fe8f6a1a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h45838c709e3f62de43c8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h11dd97bf326310df1357a;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8548da36579f3569a9fa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17ad760cfd676b9d91f77;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1cf94c14cc30380f23baa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1e2701503d52ea55ddaa5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hdb6522c89cc0e4cc9fc0;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h15ae4bca2c119edca44c5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h123ca9a8c9c139a955494;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h481490413cf3d0abc92b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1c1ae5d488c1281f57704;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12f3a078a6826e08e2ab3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hb5c87ee2d9420fb2b786;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbd832bec541898385ae4;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he25ac0d0f72503907807;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h20a093be602a5d00ecb5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h7c645cd9696ab4555234;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1906f4fb8bd92861f2004;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1fc3b032865f3cfff33b6;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h2e0c4fbb69ae6d47cc64;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1654b9db5f81dc89729b5;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h6abeb88e6b6a9b913134;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf4b4e0a9b589f56fd731;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h106f25770f6de2cc0e632;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13675f2be58a7914d50f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha549653d19be4415c762;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc2d02d24d5736256dc8;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'he6b93c75cdef9e981087;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19f4aac04775827016f24;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha7718ddfa5df568224f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1093bdad8890c16fa8915;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h120ce9ba030f396fd76fa;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hcf3e2bbb93752fa34529;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha3685d7aaab4efadeb21;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1dfd537200a7e2f7dab3f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc393b5e1645beb188e16;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h4c1e6d1b57b9fe09c486;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h5205e112cc692c193b5b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hca50fa648d7f0f4b5fd3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h135321a03d8b19df50cd9;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hc9910384cb5efd980019;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h13150c22a78a54442e0e2;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h646b89134b016603ea4b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h168349f777c5c64cdd137;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hf02048bec963417b9226;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1470ca6d876931c0c1f7e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'ha7996eb8f3c1d1191a0e;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h844caa3349ffa44b9ee3;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h80ffbf152eac1cedba7f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h8e48b00034916398567c;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h16fa676faf5432c985073;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1d9cdd0e08fb058595e1d;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h22041e964b73c2809a49;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h12afec1cd6ecb4938d39b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3eb6531d10564592680b;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h3dbecca9d976b5b72e5f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'hbe16d79ce984634162a7;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h19f1c1542876192f82717;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h17384b1f883bcec15038f;
        #1
        {src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 81'h1550cb02dde74082f863d;
        #1
        $finish();
    end
endmodule
