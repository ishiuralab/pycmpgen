module testbench();
    reg [29:0] src0;
    reg [29:0] src1;
    reg [29:0] src2;
    reg [29:0] src3;
    reg [29:0] src4;
    reg [29:0] src5;
    reg [29:0] src6;
    reg [29:0] src7;
    reg [29:0] src8;
    reg [29:0] src9;
    reg [29:0] src10;
    reg [29:0] src11;
    reg [29:0] src12;
    reg [29:0] src13;
    reg [29:0] src14;
    reg [29:0] src15;
    reg [29:0] src16;
    reg [29:0] src17;
    reg [29:0] src18;
    reg [29:0] src19;
    reg [29:0] src20;
    reg [29:0] src21;
    reg [29:0] src22;
    reg [29:0] src23;
    reg [29:0] src24;
    reg [29:0] src25;
    reg [29:0] src26;
    reg [29:0] src27;
    reg [29:0] src28;
    reg [29:0] src29;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [0:0] dst18;
    wire [0:0] dst19;
    wire [0:0] dst20;
    wire [0:0] dst21;
    wire [0:0] dst22;
    wire [0:0] dst23;
    wire [0:0] dst24;
    wire [0:0] dst25;
    wire [0:0] dst26;
    wire [0:0] dst27;
    wire [0:0] dst28;
    wire [0:0] dst29;
    wire [0:0] dst30;
    wire [0:0] dst31;
    wire [0:0] dst32;
    wire [0:0] dst33;
    wire [0:0] dst34;
    wire [34:0] srcsum;
    wire [34:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .src14(src14),
        .src15(src15),
        .src16(src16),
        .src17(src17),
        .src18(src18),
        .src19(src19),
        .src20(src20),
        .src21(src21),
        .src22(src22),
        .src23(src23),
        .src24(src24),
        .src25(src25),
        .src26(src26),
        .src27(src27),
        .src28(src28),
        .src29(src29),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17),
        .dst18(dst18),
        .dst19(dst19),
        .dst20(dst20),
        .dst21(dst21),
        .dst22(dst22),
        .dst23(dst23),
        .dst24(dst24),
        .dst25(dst25),
        .dst26(dst26),
        .dst27(dst27),
        .dst28(dst28),
        .dst29(dst29),
        .dst30(dst30),
        .dst31(dst31),
        .dst32(dst32),
        .dst33(dst33),
        .dst34(dst34));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13] + src0[14] + src0[15] + src0[16] + src0[17] + src0[18] + src0[19] + src0[20] + src0[21] + src0[22] + src0[23] + src0[24] + src0[25] + src0[26] + src0[27] + src0[28] + src0[29])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13] + src1[14] + src1[15] + src1[16] + src1[17] + src1[18] + src1[19] + src1[20] + src1[21] + src1[22] + src1[23] + src1[24] + src1[25] + src1[26] + src1[27] + src1[28] + src1[29])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13] + src2[14] + src2[15] + src2[16] + src2[17] + src2[18] + src2[19] + src2[20] + src2[21] + src2[22] + src2[23] + src2[24] + src2[25] + src2[26] + src2[27] + src2[28] + src2[29])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13] + src3[14] + src3[15] + src3[16] + src3[17] + src3[18] + src3[19] + src3[20] + src3[21] + src3[22] + src3[23] + src3[24] + src3[25] + src3[26] + src3[27] + src3[28] + src3[29])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13] + src4[14] + src4[15] + src4[16] + src4[17] + src4[18] + src4[19] + src4[20] + src4[21] + src4[22] + src4[23] + src4[24] + src4[25] + src4[26] + src4[27] + src4[28] + src4[29])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13] + src5[14] + src5[15] + src5[16] + src5[17] + src5[18] + src5[19] + src5[20] + src5[21] + src5[22] + src5[23] + src5[24] + src5[25] + src5[26] + src5[27] + src5[28] + src5[29])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13] + src6[14] + src6[15] + src6[16] + src6[17] + src6[18] + src6[19] + src6[20] + src6[21] + src6[22] + src6[23] + src6[24] + src6[25] + src6[26] + src6[27] + src6[28] + src6[29])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13] + src7[14] + src7[15] + src7[16] + src7[17] + src7[18] + src7[19] + src7[20] + src7[21] + src7[22] + src7[23] + src7[24] + src7[25] + src7[26] + src7[27] + src7[28] + src7[29])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13] + src8[14] + src8[15] + src8[16] + src8[17] + src8[18] + src8[19] + src8[20] + src8[21] + src8[22] + src8[23] + src8[24] + src8[25] + src8[26] + src8[27] + src8[28] + src8[29])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13] + src9[14] + src9[15] + src9[16] + src9[17] + src9[18] + src9[19] + src9[20] + src9[21] + src9[22] + src9[23] + src9[24] + src9[25] + src9[26] + src9[27] + src9[28] + src9[29])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13] + src10[14] + src10[15] + src10[16] + src10[17] + src10[18] + src10[19] + src10[20] + src10[21] + src10[22] + src10[23] + src10[24] + src10[25] + src10[26] + src10[27] + src10[28] + src10[29])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13] + src11[14] + src11[15] + src11[16] + src11[17] + src11[18] + src11[19] + src11[20] + src11[21] + src11[22] + src11[23] + src11[24] + src11[25] + src11[26] + src11[27] + src11[28] + src11[29])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13] + src12[14] + src12[15] + src12[16] + src12[17] + src12[18] + src12[19] + src12[20] + src12[21] + src12[22] + src12[23] + src12[24] + src12[25] + src12[26] + src12[27] + src12[28] + src12[29])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13] + src13[14] + src13[15] + src13[16] + src13[17] + src13[18] + src13[19] + src13[20] + src13[21] + src13[22] + src13[23] + src13[24] + src13[25] + src13[26] + src13[27] + src13[28] + src13[29])<<13) + ((src14[0] + src14[1] + src14[2] + src14[3] + src14[4] + src14[5] + src14[6] + src14[7] + src14[8] + src14[9] + src14[10] + src14[11] + src14[12] + src14[13] + src14[14] + src14[15] + src14[16] + src14[17] + src14[18] + src14[19] + src14[20] + src14[21] + src14[22] + src14[23] + src14[24] + src14[25] + src14[26] + src14[27] + src14[28] + src14[29])<<14) + ((src15[0] + src15[1] + src15[2] + src15[3] + src15[4] + src15[5] + src15[6] + src15[7] + src15[8] + src15[9] + src15[10] + src15[11] + src15[12] + src15[13] + src15[14] + src15[15] + src15[16] + src15[17] + src15[18] + src15[19] + src15[20] + src15[21] + src15[22] + src15[23] + src15[24] + src15[25] + src15[26] + src15[27] + src15[28] + src15[29])<<15) + ((src16[0] + src16[1] + src16[2] + src16[3] + src16[4] + src16[5] + src16[6] + src16[7] + src16[8] + src16[9] + src16[10] + src16[11] + src16[12] + src16[13] + src16[14] + src16[15] + src16[16] + src16[17] + src16[18] + src16[19] + src16[20] + src16[21] + src16[22] + src16[23] + src16[24] + src16[25] + src16[26] + src16[27] + src16[28] + src16[29])<<16) + ((src17[0] + src17[1] + src17[2] + src17[3] + src17[4] + src17[5] + src17[6] + src17[7] + src17[8] + src17[9] + src17[10] + src17[11] + src17[12] + src17[13] + src17[14] + src17[15] + src17[16] + src17[17] + src17[18] + src17[19] + src17[20] + src17[21] + src17[22] + src17[23] + src17[24] + src17[25] + src17[26] + src17[27] + src17[28] + src17[29])<<17) + ((src18[0] + src18[1] + src18[2] + src18[3] + src18[4] + src18[5] + src18[6] + src18[7] + src18[8] + src18[9] + src18[10] + src18[11] + src18[12] + src18[13] + src18[14] + src18[15] + src18[16] + src18[17] + src18[18] + src18[19] + src18[20] + src18[21] + src18[22] + src18[23] + src18[24] + src18[25] + src18[26] + src18[27] + src18[28] + src18[29])<<18) + ((src19[0] + src19[1] + src19[2] + src19[3] + src19[4] + src19[5] + src19[6] + src19[7] + src19[8] + src19[9] + src19[10] + src19[11] + src19[12] + src19[13] + src19[14] + src19[15] + src19[16] + src19[17] + src19[18] + src19[19] + src19[20] + src19[21] + src19[22] + src19[23] + src19[24] + src19[25] + src19[26] + src19[27] + src19[28] + src19[29])<<19) + ((src20[0] + src20[1] + src20[2] + src20[3] + src20[4] + src20[5] + src20[6] + src20[7] + src20[8] + src20[9] + src20[10] + src20[11] + src20[12] + src20[13] + src20[14] + src20[15] + src20[16] + src20[17] + src20[18] + src20[19] + src20[20] + src20[21] + src20[22] + src20[23] + src20[24] + src20[25] + src20[26] + src20[27] + src20[28] + src20[29])<<20) + ((src21[0] + src21[1] + src21[2] + src21[3] + src21[4] + src21[5] + src21[6] + src21[7] + src21[8] + src21[9] + src21[10] + src21[11] + src21[12] + src21[13] + src21[14] + src21[15] + src21[16] + src21[17] + src21[18] + src21[19] + src21[20] + src21[21] + src21[22] + src21[23] + src21[24] + src21[25] + src21[26] + src21[27] + src21[28] + src21[29])<<21) + ((src22[0] + src22[1] + src22[2] + src22[3] + src22[4] + src22[5] + src22[6] + src22[7] + src22[8] + src22[9] + src22[10] + src22[11] + src22[12] + src22[13] + src22[14] + src22[15] + src22[16] + src22[17] + src22[18] + src22[19] + src22[20] + src22[21] + src22[22] + src22[23] + src22[24] + src22[25] + src22[26] + src22[27] + src22[28] + src22[29])<<22) + ((src23[0] + src23[1] + src23[2] + src23[3] + src23[4] + src23[5] + src23[6] + src23[7] + src23[8] + src23[9] + src23[10] + src23[11] + src23[12] + src23[13] + src23[14] + src23[15] + src23[16] + src23[17] + src23[18] + src23[19] + src23[20] + src23[21] + src23[22] + src23[23] + src23[24] + src23[25] + src23[26] + src23[27] + src23[28] + src23[29])<<23) + ((src24[0] + src24[1] + src24[2] + src24[3] + src24[4] + src24[5] + src24[6] + src24[7] + src24[8] + src24[9] + src24[10] + src24[11] + src24[12] + src24[13] + src24[14] + src24[15] + src24[16] + src24[17] + src24[18] + src24[19] + src24[20] + src24[21] + src24[22] + src24[23] + src24[24] + src24[25] + src24[26] + src24[27] + src24[28] + src24[29])<<24) + ((src25[0] + src25[1] + src25[2] + src25[3] + src25[4] + src25[5] + src25[6] + src25[7] + src25[8] + src25[9] + src25[10] + src25[11] + src25[12] + src25[13] + src25[14] + src25[15] + src25[16] + src25[17] + src25[18] + src25[19] + src25[20] + src25[21] + src25[22] + src25[23] + src25[24] + src25[25] + src25[26] + src25[27] + src25[28] + src25[29])<<25) + ((src26[0] + src26[1] + src26[2] + src26[3] + src26[4] + src26[5] + src26[6] + src26[7] + src26[8] + src26[9] + src26[10] + src26[11] + src26[12] + src26[13] + src26[14] + src26[15] + src26[16] + src26[17] + src26[18] + src26[19] + src26[20] + src26[21] + src26[22] + src26[23] + src26[24] + src26[25] + src26[26] + src26[27] + src26[28] + src26[29])<<26) + ((src27[0] + src27[1] + src27[2] + src27[3] + src27[4] + src27[5] + src27[6] + src27[7] + src27[8] + src27[9] + src27[10] + src27[11] + src27[12] + src27[13] + src27[14] + src27[15] + src27[16] + src27[17] + src27[18] + src27[19] + src27[20] + src27[21] + src27[22] + src27[23] + src27[24] + src27[25] + src27[26] + src27[27] + src27[28] + src27[29])<<27) + ((src28[0] + src28[1] + src28[2] + src28[3] + src28[4] + src28[5] + src28[6] + src28[7] + src28[8] + src28[9] + src28[10] + src28[11] + src28[12] + src28[13] + src28[14] + src28[15] + src28[16] + src28[17] + src28[18] + src28[19] + src28[20] + src28[21] + src28[22] + src28[23] + src28[24] + src28[25] + src28[26] + src28[27] + src28[28] + src28[29])<<28) + ((src29[0] + src29[1] + src29[2] + src29[3] + src29[4] + src29[5] + src29[6] + src29[7] + src29[8] + src29[9] + src29[10] + src29[11] + src29[12] + src29[13] + src29[14] + src29[15] + src29[16] + src29[17] + src29[18] + src29[19] + src29[20] + src29[21] + src29[22] + src29[23] + src29[24] + src29[25] + src29[26] + src29[27] + src29[28] + src29[29])<<29);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17) + ((dst18[0])<<18) + ((dst19[0])<<19) + ((dst20[0])<<20) + ((dst21[0])<<21) + ((dst22[0])<<22) + ((dst23[0])<<23) + ((dst24[0])<<24) + ((dst25[0])<<25) + ((dst26[0])<<26) + ((dst27[0])<<27) + ((dst28[0])<<28) + ((dst29[0])<<29) + ((dst30[0])<<30) + ((dst31[0])<<31) + ((dst32[0])<<32) + ((dst33[0])<<33) + ((dst34[0])<<34);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h707ddbd8cc86a7ac8c26458173fec596a8148708831389e7169c83e0269f815f4a072b655be5c9622d4fe95d6256f1900c8cca7aa7cce64cb07804050200eeda863a68753175dd27d0ce2f550726578ce14fbd8705f8f85d1ff499624c203e3947cd3d9729665b00608b62e13ee837c1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h379d0b6018368b5fa385a38202d85b31350ecfbff90b6cbd0ad2986f2bbde71871590f7de420766f0d34ded1fdaed570a630c250af7bc3cd64a96b6f3a13a41499c432940c0ff1813c0d3cbafc5f704d4228aa8d19ebcacda8eeaaabdcac895f40cbd648e1da2cd253702009f6f06732f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h417409866afbbf9ac35da2f7db4690dc4d7986050df6eff4bdeb5152b1d68b4370037d2489ce19d4a7c17a056392ac45eb32153bf92b97bfa8c7066e2809d1f1dcf4c3c106de6c553708da17e49f7f625108b990c2080ded5fdffb2538c27919a6701ddb83f6927a117033943347bbe8f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd26d6ed2ba6ae42fc93c9b90c2f28c7236b0d8a388fc02095e70f7512548e506039ede00b3088f48a99f933835e853776d988b6852ac885b306261b1a7d36153f4af24485c143b4259cc4d203c860e1819a73ab775ca8eb7e44dd1e79b7a5f2f432a44c3ff487f386acb6d5fbe6b85a41;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22f3df5cc86b648aa9646af6325d0bba72d19f0a538855ae1756b64ba9c714d9c65ca9855f299c90e0d3d9d422b8bbc784bcf0a134ec8779293a828be6fbd4d556e7f1cd6da42e85d7a81bc63a3209d8b8755312186b5d1522db997ab04962494a3b2cd1d08fb29cf291889ff8d149a35;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78e08a9233c058b45db1036f8e78ab764dfe4efa1b2aa23d9d7dfd966ca4b9093a6329c393ad86aa7b78c0376fce8335b40f94df1b5445cb140508cf65b4ae25d4903ae6765b3e1eda16e945d3151939a0574b48f35bb24fc5460cd5edf5a65a5dfd29827be420d2be06011d7a0779b42;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee84cd5661a7c57581dd949bc18b9cc149ee4566d41890b3208721e4e0df07265627e18fdc9d14286dbfbbdedde972bb3c01f03bac4c4387faf0fe6bb14278e859ad5aca2e8bc39a5f20c02475cc0ee1371f2f03c8e220a03854c8d4f24c61751e3efcf001a55a76ad3018cb5cca596eb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6191320d000e9dc1c643f8415631a7bac1f57959e651508cc5a49c032a04c01ccaae706b4ee44165d5cd66355bbe40d48ec70fc91336068aead8b4b76aea8149ab4018bf4b2bf3f52edebd912dfad4740295f70331c726d5e89627a91f9d8eb86697ccb3ed13458381b2a2501ef1b0b7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h521745f0d43da8151a40266280ef3697111257ae6c2896918e3a93239d5e3f9d9bf868f1c9c2136c149e6d14a701c7e84cc505cc0db68e9e709f0be1b7aca6908bf0142c213f91581b993a930a33e05a824ce1af1da93224d9a41c4a059264e7243dc4e34eb0c050b92a715eeb78bac0f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h13e8607cd27aba7407a4701d6ecef3e9e302d92da307d19b9a00c30d7cf8a340a31700a5c057024298645cf29a6a903d50b396ca6e3c78cbb3b86eb028353e21af7c36e27ae3f4cdfbfcfd05d7e98c3d04992684d5e8a0bf43fa09bdbf667c0d315e7850a454fb7d56d0ff9bd7f6389d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d10f9a30cba812dc7533774d689ab792a8a9b058f4559ebcb4d48142ed8a475b04038d4ca80ccaa2f5a1e9b7f8163832fa3bbd3c7fbba03d2e3d2fadfb3666a5df2c8e1214d6eea1571e48202f321b0ac1a48f8707ed196fcfabfd504cff9032922763f297e1be6742d2c8b5ae573784;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c93a3498fecef0197ee1b23e884095c577f9c3cc7fb6535c31bd5505d9182cb1f130ea8c95eb3aa5ce5d87389a7988a3433923bcd02373f3e6ab3c1e5b9a845d40bfb8fd35ee7f9d8bb354e54f1601c86c2055230c84fb7cd185864e2e0b7fd64ca58fd950ac9178b07fddd629d19942;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc98348ecaec9625bdb025c17a6be2e8e2a4a5693977d9d5a1a7097fd4d132a5678f8523b9ca89284dee61cb448541fca75c44d228c429d988c00a3cefa4044b71ff6086c7c7e509cd8c8a731bb009c4e240821c93de650218e02b01528f9f1f8c90198fddec4e33caffd74e0bbea52572;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3aec3ee880c6679d2aec9f42adb2999bea9ff0b0de97ac0bdaed0d2b02a394e39f86c5d09ce5984c5642c2727ddb33435f70a63e7d24e2d8cb9b7b0991c2095439f2f8b00f9fe7378f25ebf05a7a807d11c448afeed241e8d5f35821253c218dc1a7ddfa9bd703a0edcf2b1db37f6c2f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc85c2c5b359022311efa0143aad8b1e3a5fa0930585265c04b5fb600c6fd33cf0f0801681aab88d9fe030e0449ae9d72fb1986a7ac1923a9dd124fcf559b7795632ec146d5de72676896c398fec701a9b22de1c2abfc26fa74a0a3057657bb9f5e61981225d96cb06de0a30747f95b4b9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6302d625a42b1a1ab67916a8cd764d590c692b0d3ff8f55f18bee9f85e3dbf64d21991eb8a2ed2ee38bb7d99d5465d38cb559dfdce621a3dc383770e99306acaeb3defda92b6aa015ba5cff9ccf16f3249bd317e2c5d40c62f4311047e8255dd3a52081af8d246995e14e42897a41474;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51c5acccc61d478a0a33ec63fb7d3e6d64c342bc7710b7c49f278a63052f68dfe481a947fed5339884fe72cc190b8fb04ac9b71e2ff96260f041447f4592dd46e88f5b5f8b0814389e4e53f981b64e06c8f4b652f3ff33775d4ffff47de61535950213d593d5eeca4f7fc3d951c0fa0fb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9cc20cd403054ab5226fb49443e5a13b894f311671940d5358556f403a56f7f8c77411f5f39f1d46352999aeefc142c2f6588b7716579225affe6d3f05c700c0b1ca9aed675ff6cd0c3cc8cebec25e72884e3cb00abb515370e6e1be139017f8f08c5007b7a76e730d6f2eb6b5590121a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h403a6a625d670fc6b45687d5c6fe88824c6438af253bb179b20e5250a3fbaf7ebb261503d0696fc2c5dca3f870203c8b5f49f7a3b400efec6d48377642b1d61a5c7788f4774c807e334a44c1541bc75b972b11f70e42291468a86b2d3eadbdfe59e580a0579592393f41a52075f5455fa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b2fcae1f094bac2dcc39e652665dbb5a341f6f20fa85cca7f59211b9a05214c9631bf2a51cadeb8a3038ccfda5962e252b6bccc39c275f7b10f97d070ef0d63f0c320b1ba5a137e63c14be73ac3babf9189fff28b2f21f5a59ddd9a94862508b89c075be10195b5a29757c720372222;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha31bf044bfb0a93025c405fe4fedd44aa2a6e7c0390d47066d431810e581ba64d0e8eb14fafd4ad01e09b3f8a3c036de32768f8fc52ae6e66d7facdeb14c45a3a302cd33cdb3938b8112189cd858baa7a4e1e73b76a8e79dc6001dc20f1e419c62ee960cf731a3e737ae9d39d8023fb13;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44b205ece99163ea30088c9fc653f1d3d5d33ed81e2e56e6f44bfb18d736dcf46f530629538ca84ed327af9647baad3e5cd14f7df64a7e360d3d2cd9a091ea6b9aff3cbcd74b9eb7417e579ac7a0f3f25b9e58b1d820bf1b9805d94569fd29826b507427794b66f1d372fb26c57ad1e5e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e0228b69a5e2d1e793278a6a9855e28b0b74711685942ba4ebf05320da4f23e1ceca5e1580fc3c901700703e6bd3ee05489a779b8c3c0920ee283da53112b6065f471647b20e060ce3b1ec13913a94df50f0e64dbd1fa42158412f00c1278e8946845bbdd1fb45b8b94ac33fd8378aa3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7084c34f6666d73208ec44bf117d11fb9ac10f2f756e55340257f47925b5436ce15636752aa224ea8e46542d112f53a6ecd6a23879d63ff9177e11e84af222839efbc7d5d727e01ff9338be92231a2e67959fb7a481f3edef602c9182fae67502471eb3f4378acce7d5b880387ab18c6c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6395129dfd7d2e970cdec2dd57c6c28cbe8b410aa4cd6eecec79750c89c370558247b28ba690d727463fbfcb0eb7295a481b1034ac268baeec71c065897029689183bd34ce1085df68ff6b99e05886809add9b1ffbd4da6a760f273d0f6d097716d8a821fb461ad5bda85c7c8d60513fa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa7a722a2ac19aaf9da6d50ffea51948ebbae3df5526a5548b7f8ec27d3a5f20613014a6a8fcd72da67708241b09afe5c9ed569e5378eaac85df35f0c2abdb88310019df651e83e35bf166f172afbbdf633e1f9c6e6df3a24180f81c5af618cde2a25ff7f7aa6247fc0441a9ea2abddf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ad7ff65678707b12f00045aec0362bd265ce7e725997b5a43a8f08601cc00c7589c4118ba9560d0e24c9019bf5be0ab3735095b3c20144c36b471dd20d3b5672cc80c24271c3e6c89f6233ba8cb437eb36557f0196db3df13ec949f474074ae5418ae80c96633d64d21d4185fa2887f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7dcf6fb05dcfe331eec19fed5b6ff49b0854e34f93ed24e94217be7a850177c7cce71451dee2b252f0a6e10a1d14416b765eb4f45343893fa1e7deb483796e4c053b902e6e5c745e4a449adcd5285c48678884f54930c87958d18233318361443383de5b041d990b2af54fa5f71124623;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e5a388a77a82334dd2c16a17f5d692a0b23adcdf480c399a5ad1cde6044d78da476d5c62ea68d9f1c646154783af4308697b2dfea20824020852eb8af4c0ceb5feaa67e3a6c16430fc6ef3371a3f78040294839930cd9fcf6fac7b52e23c818a649a6b37ffbbb2e975440cfbb1e32578;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d072e361a8e94def95b600c99b68b8a77dffed9bba0bd4ec8866ef83e08df19d49e3451b1992bab2ed180d979d29f492c0d2e09204c4d6ac9a180611c3180dca3197e2346429b601aac2682a18b43d71fa5cee9df402e8c24fb21714e02e7f94cc649ea3058a5d386946e6f793f8ce6e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45b4762bcc5dcb387ba6459c0a664df1279473a4ec4d0ec2637ca0d966428a75aa30afdb1cb5ca9a24a9753f0b31617871e7a761931fe92105aa3298cf204119b5865d807a34228cb74af688614e9805587531b9965fd1b0cef81ea2a959720e363dd6ad4f97b210cc11dc723e4374471;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h454ac826bef2d44ee1f465a22d381769053033107be338fb21e34daa9dd18bc52deb93d409612ccfa9a5e8db342cd3a99306737cc9f11a3a87d6771560a54ee18d1bf941a8c8dd78cc9d2e8b296220bf440516c03e37c1824f7c3b99af263b976f53cc82bc093ee4189998b68f0491ada;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6dcf84cd89086f49efb69f5e03256532587a6549311d3d35c0bf9df7e9f3640170f74b61fcdcb4fc5ac36c2bd368836df5cae7079d7ae6f431b5c506e30cdb7142ad0f44e18481dba577463be55adbf8c1603e467a168d5ddff843870302650623af51cfc51295f83d04f374a53e25021;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4498e1f70cd18422ee3c2b2b5ba91e63f5b6d291d91e7dde379cfaba1e6cddc8fbb7597907b3fb4d9509863e0c08ab9f338029296265bfc022e54f6d3bdefd5a2befd085ea0b2902496c77f4cb933e0a391997b677a6f386153f7c02c1909884d5be71f4b913b5d579d90623bc2b87d4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d99cde79d777eef50fe204fbe5e0e59ecb8bd92291fbb721f69d433cd18e32b8ae17db9bb097374ff0a658bf215f57753f4864b4d50b3229be9fdcfd89d6379b3347f33ef9fd7719887742775e761985cfcdf5e0ad64c4460bfdbdcf7dbe3a7a2d8d087e7da99fe40a5a6b049b29dc2b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h99206e6bca0556c3e47bd2335c704e6041d9641827e15037369304ee4d2f1e534abe7fab8df6b196085746daa461d8cbed6c077b86e5e02902036cd03cb5605419ca09a4b70e46092c6556a2e4b92390d5ea0b6ccd7a4dd575d22fec67f7352332e9a21a55389c61ceb90bd182e4fa4c4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h909719685e247af24118725a1440fa6d7bb070404fbf54dbba3dc1059ef67fefc357b9ff58d29cf05bd9aaee3aeea88803816c46f52ad0ce86e2526515b152aacb52d57beffc9df2df9e537bf43bea5017c5df1b2fefcc37ce758caacdf3dbba9a3f867faed1ca5eea7426b48f7fc1c4e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd254f612d97742eaace1b23e6cbce5ff844507816d5e0e8673224e2717f077567765889d0b5a51200a0ad3bb4cb6eeace4de60b5e003283a17b3a9c76ef0c4cac0c15465768aa5f504a1f3eee629e5faba7677273c978ce2789470866a78672bb35933b83f819ae23135157e89a6721af;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb5f3e4d4b6e9e296c34c3c2b84133559732fa8505cd701b894cc11417a7909bbb614417fca5747dc2c0bebbe5bc614f7ab18779f6f0ee7f2e0f37c2803e759565d9f2dd1ad5771305150288f68e4c69c86f3dfd474efc328e1559e2d891814aa868b093408e05c326dfea0f696ac8d2c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55e1f20e1706e198a63194cb07b581f304ba7ddc01ebb0e90a5860318ffd1d11c00f55cdc6fed57318a06bed30150d71ef99879d91b1e106dc73780b6f88a36805b972f20800d4cfacec12959df0b933bbca29784353bce9288dd2e4cad65c80397ea99611c83ce6e9edb3244f9553eff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0e7b73f37ac371f1a7341dd0f86a4132bc2000b9524ac79bfcd94d6ee3b19575a9d90a5101fd5f776b46561f355f38862cb8c33a0943a0e11bfdf7c29de75ac0a381820fb62330db62326b86d60719c5698d4075efec72cbfe598cd99e6eeb940c7f8a4cd7f295ea85821deee50c2fff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74f394d379927df46269beb1ca4b141b044c56dfdc8003182d6410392c1866c52b66090f22b3422b751a7a5628f880b29cd50308e11ae33ee942e68960377a85dece488a7f6f8c1440dfa8a8cee6eb4f86ba53f12047e7321830ee892ee9bb230dd806ee1184e845128ae8b60a5d36ab1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfbd68424f7ca790dfdfa74b86acbab020639dfeee4590f70eaeffa9cdf0ec2765bd5b6ddd174fa03dd14585db35769a0e171263b2d5abed1e049fb740fb2c0b67e10c0b6247b7049140a36a78c133969831184253ec882fe888a7af15504dedb0273217210200e90f5b8ee1272784a80d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc77b0c269e7fb8b5847db2936739de94288a1892af300d5132139f5ca10ecac10d2c482b8321d0e6f7f35caf43c77f5b3834e1b86e472596a4e7af891ca782b33eed35d9345206fefe35a814388bd97752b0291a0fadce9f3efafa05e1e5ca8483a9bada85234996523fad6647965ae;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h572be9648e94e2af981c676887e93c068568a29c6f1f1ec2e1b3160d3aaa31953c8f561e872f6bed3deb598402cf51fa2aacac87bfac6b12eb5659a86f11f413373143114b58e99091060062eec0c2c4a01c054ed3e3d0292aa95bc2e675d3a2f029585bfefb7c3478dc854c822acafd5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e97cc1631421e386d5d9ea5a40b4efa5513c6c1f3186ebe7f4815fb0a251988d75f4ace381f4e05feb0c8e5067affe8574b54d6dacdf20481808c4bcee5ecbed8fc2a7f82720ba6c5e77507a5c6bac9fcf2c8fac4ce3f15affc2dfa9662000e22bd78e55110b305015a742f2a43d67d0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h16810b54444de0df285e3e58dd598d657e9a12ec6ee9fc86ca641d0a2a1dcf8c4a5382b601656c6a577019fbc320488f60504bec51a1102c1e3aa9159b2a7827b6809cac20739e7f866746e9a4093d773ac147471a1cc61ae396091065726c2b7379cc8fced61c7f81846d34b1a942b88;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab033d8a0f45ccc2240de374b3176b2ab4131c9bdb2c65fd01c41af982076fb06c1badcded1fdb94d1e06e50fafcb6d2425ed21e2d9c8262c1e1182864401b080b6c9e5b5787bb6ede17c5a7c9d7087cb205602ba06b0acdaa89f419575a2e7650a6050b35dafd278151f220ce6f5cdcd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4acd88192e4445956ca01f76f85796b7bea014095109cf1cf35de8b33b93a0bfeaee8a5f322d7118b5907c5ea34e98efe86a6d14024143cacad1268d44ca50668151c42f0b99600148a2ea8db63ba61fed80768918f2cb0589fcc88486f50f02cd8b0db8fb98bd918745b2d25bf5fab10;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e7c4609057a5cb1a7bae049534e538f351ae626f1ceea8e2b0c9c7b4b6e2264641e6041562120b278e742eb065656d6976e7f50464a2196c5be0e8e4a9968eedc4c4767da92efd2bd5cbc14ec2d2d600112b4454d316f98ae19407dd338a1a08b8f3fe9269844f7eec3bfe4793f31a8b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2fb4102652a5ba9baa8f99b8cabb41a0f0efee97d3a6b066d99a41ae41cd6754de49c6896ebd992ead69383e2f6c2ca31788f3fffd65cd11b86d399063ad639a1baaf937b78e88b10d9b0fb1c4cacf52d5f7b7dbd45cf6ec1ebff68e80840a0637175aa359659836ed7dcdbf8ff01954b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88ba3d2a586ca266b46bb2a960e5989a363622b94e646457dd3a60b576ea8759ea43035ca8a24c089d8e350ac80ae17f9362d725b7cd78f50cde361c0be7432b1eadd70eb5d38d73ed86dbe685772a3635a5e38ebd3defb8396480ae507a5c8e4a3a374992d1f7b2f516c6a3a73750c1e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b6dc6ff0d368d7033065d2c75aa17a8cf4346e31f96c6ee83fc70737975d98c9352dd6ab7a9aaa154201d973a90a42efe8ed6553c5eb3ee2004d1d99aef2401f654899dc7e0ee80649afe3de508dd1f77ad01e21429f83e98e21910364508a5f143ecb5461d67a334d84044f1bf950e2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22f57a6612449cb00ea3b78ee6f3438e37e5ee298b8b0e063ae6afe605593addd1df7b24f848d00042dfc3eda8a84ca51d25d25eb66419065550c3229ae5530d5f9c2a2de82ee14bedafe28d3f7fbe6b963432905191453db96629277742253ea6f169ed4848328646325b977427ee449;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha0303a15ac03349c2cdcceed1ee547a9729130069fcb09ee681e50bf120794b70972ddde7a7a622c4b4dd065b83f75f7394fa70de24eec1ef8617938ed42909a99b803df8c1707946a603f5fb8530b50c1876f927f9ef02076e679e9d009a48c8d0aeba2160d8d566e09611ab1ea5067d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf78c92c301853b594638b607a31c4b9f95f6e5c6898a39b18496065b2e28d45c797110755ad185b51055833cde787b396906d0ab908bfa9cac7a921ad82baefb0c261d7699f3678cb757f6468cd9942aeba93967a53997ad67a53d3c90d8b416e50d1b12c6259d768865902b5be257e2e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec678f831185a84e2a8704d8385bacbc41b796e276e5e7549325dd2793919d76ca1e9b0fff8b546613a35635ad62789c684ec6c843cb8ad88e5bf0771c646b25c48f56ce65792f80c4d13f843a7c37309739a3b5a7419345b89151d25a213460202698388074d1410367843b42515d9fd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h463b8dcc1cfe9978c7752ca2e907d5a1447c87713a9acac25dea5fbdfd60ccd016c37854ea492987cd3f023eb7ce8c4c6b258d529087af03d0e89af01e0d88b100c085189ac4dbd98ea606a23c475107a1be5760c0bc696af41df7c5ded3c51efdc8d471361b991fe3e536563cd3eaa1b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4cfcdf7ee8413cabb557b6aea64fc71c2ebbdccfe62c590478e2bfc8d57ccae7c4042e25d7c09141eaa9d9d0e2038d0250241488089a366d03da1779eeea4d762e047ca584f60057b59a9452da395b92ac1f893a8e3ec562f341cd7e632c77adc1f4c07303c361efcd821f889ced94b78;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd9f6ed472c06825ab6d2e9ab5447469c08e1dab5fc1a766b4f929d87f4d884db7f1b2c357f0b2b7dae2e448097f1a812afd9c4f06f30b038e08ed4de5588aa5c38e3ad55e41f5ecbd2c75e867a89562291d10e9cb4abe3e8acbf7717daced52377cbbfda4137ebcf5ef99451b5842cc3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d23fd43e126ca2a217a00104916396740ef1ed4ce4eb2650911600d672f614936f88239702202dd8c3d2aac8f7d27b5ac737b466eb330ed5eba1ecb4bfedfac02d3ecc1b4b6e991bfb0c053b7d60f552487bb1b15ce5db6f7a924fd84ea44325855ac96dd0f160456bbe6dbeff3e17db;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9fa83444d8ef2954028cd635da1f663039321843d1d95b1ad50d7d1ce2ccacded6795dddbda31b042fdf2cfe658d9641a0f40275bbc5b56dd50bb1e18cbeee7f0144748b4282ba4d1a193bff6b7c5a0c60c19f581ad93e159b99c543b6df46d70ab2f437ebb2bb31c9101e0d5d2fe9880;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32567f60bbc8b81e513f68553b75a2b4d492d6886f2e28a2610f3b73bf5e544ddd6ced185bbe1b51030c092bbc61301ff09de3a76591fe4c6af76ed698fe215e8bf23d11308ce8fd575a1b3b58cef61cfc15ddf30fdff8c3c4279ab0b1f4492e9a67cf9418f463a98a4dd24b2d6f81641;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4280893266dbc9dfcab04c8e9a71212e494df98000d310fad4d1a352f3d45d47564acee8de85e55700b03200d0574e0c48cd168152165dcb92af9de8b65716b47081bf4108989b0b7dfc457a5984acb0140cec009086dfdbdca6e55fcca84b963df94abc33ff391a281a63db96a127226;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc4142c40668c556564970f69ef47172a6f1af4b6f57faf4f039d915f64aa47338428a5f93d12c83896b29f409ecfa93b4388c1194de96f62bea3699cfe014068b1ce51781433e5ac27e4c8566889924182dd6e591164c79e50d6e8f6e653c6539b0838dba7186e5e160a231f37dba67a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc9169ee725ac1010c42582d5d573c3ac8e7ed5ecf9bfa0591f47856fb9160403f773b428dbca445d986548c02ae704a937a147e3d24e038db19160ad3cbaf7ab441d329689965fba3fca24159580ce5b4836a38139c48d2ab43160f9a876bd38d52e2859abad8d487a5f68b65de97a0d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f6e15a0e7640a945d99e6d5652c71e74031391d56c385560446c144bc9e55239ed452f3315c7e97ffd25d997c0aa8c45ee836d917cd7ea16a1dad0b7ee73e9df60a2919332b5ace0abe5e2bcf6379220168274616af3a712350cb25ee00d03d6fab1b4da360a2a2146c35a087caace27;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee5007c4560180d29411b63ebd8c9c1bb3fb9401539c9c403482c01be0f5897eac3136252142b3750b565d25c74bfabf28ff0176b86b1ff71caf0cdd8d98db414a779ebad162395ad544b0041d82ab5d004130e22ed45c031a4174863d9199136188e6a124b211f05496a5a74d75b78ba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h485de20c16dd746cacfb0fd60b0b7fb0368fa25d497061ea307ff8d0583bd7cc54a281a6b8a508de20dc00c6131e502230e50b85d8175bd0f7c8b37881a89be96705a83fa09e8ef6f04fe0278573b301bf8538c9cf390d6397b2368724c4e4421ac7836142699e3bc1f5c7f0c3978347;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a8b379599766c04ad84f539828a79c8847d7c4325177e06b82d41c00c706ad6bc272a2f251a6e64986250781425721e5ae7cdd3d328f44b39943502400656b600843dafc195c69b6897d17f3c13ed7c99e246c9a3cfc137429877bb11d7a16019480b7950da8f562afef3c78eb21fa11;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c6d99010551ef6fc99a715f73a15ec736e72e783ffd3eb04ca654abe9228d3b889151dd3a7d1be596bd6387abbe7788a4e525fde7f9bb7c14bd543d03525d5cf46f59c26d6536eaaeab53c8b91647b58a01182c23d99710b13024330e7272753b0c5208a021867dff50034e2d1b6845;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93ae201b08e7ba47f65e1c87c8dcb6e2c2b403443b0d97a18bafc94f3e52cb48e1f5e9e47629f908f311bdc47292193b0a5a538dc6af105d248eabc9db93e6485b16ccc5ac210ccbd27c2fbc3be5962656efb85e525cc412fb1f92a8954f7028946e75378836d14f875659ff85e0efed7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3865628272326cd944cd301a5a9336d48e8a5bf67e979a3ba1be14eac8fee57ccddf3bbbad6b58ab3facf1c9930b467124f7525e1d2557844087d2661e693998edfe4c0c767cb385686c2c5f783485e1e29631b34b3b6da8661873b88a3b147fa4c56c967db5823c10f012305ff2eeef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb65de76bcc0243d968caafbbccf54395f15ab9d409505315461e4299bda3d8136a10562819d9da3339b4c32e181cff0b19f9f0c3dca87382423126ffa0a6f23951555a79c40a299f99006b0f35a2652d08dabe7a1f2cc9aeb7e44f8fbba63a3f59bf6608696a115714fc13a3fcdcc4f2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb90e2a448b74f45a244b7c6c1e9702cdf58c8fd15847e391ba9dc5e2171a6e21d900d7856e0e154cf61096b24fd951c600eb2cad1ac5594b0ae665affab3c8ff045800c069f6239aa2ee642d4fd3c56b8ea5186c924957615022dbff01619761c4f742dda3b55b240fd89da4607ca15d9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ca4505a04bb111b3d1ce04a6b81c53799d1166d8a5b6e165947f132ae503ab5e8d352460f2583764a5e7ed8dbde24f9b9d49d07f21b58d2c6b7688f0fbe41b5e0c824f31df4e3432763ef70352373bef93ee659de6ab6eb186f3faa620ee3e0f1e4b8acdda2ca76033816eb1665dfe11;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h273da0ffc803b83484fded0e3a77f6c7ca5e61f100ac377769227b85326531dd0d7233b4b6b0840448c5939c88d2884de7a595a857efb094004b7e6a8074893044452647e26a27106f610608503ac96e352c6b38136388a15f05404aaac45155c5a9e48111728d49b7dc3b67aff18d82f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h815ee038dda4d0489c4b7159b32008e971c165c7557156ff60d1fb52e6592a10ab3980842de26b786a28cf2606aa6beb233f744358ffcd08f049c27a843e5a36b2394819471699340e09dbbf7c4ea40b0e201f542da23947b66ddd0c0f1b91d92392983d197d63a9598d96b5b787ef9ac;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec6e2e478c16905f20d02167e634065d9ab73b0e3f79a76a6f62eec29a7b255dd640a525a8c11428526a8b91ebaebbefdaad70dd1a6011dcab1d1b01408a8bf90030b4d40e688c8f7cbb032994537ee3e4ea0e49e56765964ccc84a1782da73e6a3abd1bf234e486dbffec0815f57b5be;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc771478a869f2b6b4c39b03e07426c85048239acac73d6881ec3a379a3db56f0d4e89a05565344a473ad9e853dee5eb74759b2d113fe63a9c7bc7bfe0e6fe12ef13ee93c8119714eb2bf1d1504eb8346b39f89a2665733724b23862a04a16694cb235b339d94378e22518c07751e45246;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hade089c6fc3008899aa51953c5362c745c5dc08207d12d1d23a87b8d10ee9ed444db8c2dd2e887042afde6553ebff023cc8b55f27d766a7b972700d1014dde21b1c65fbac923c5a239d143b8faf3c445474201bf7f90af32ed4ba65d4925a33288897fddff1b60c8c2449b27f0e717ca5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1cf0c6c6cdb62919adf1db877ba48e08c9947bfe184475c440ab8dc704470e0e2697ed98271ca12c9f4b257810a63f8b9215e13ad7d5fdf192016ed2e6d5f0f200dbf64668d6c13f1aeb400c2a057dc30678fdf501bdee781c6bf20adb9e3b9551789591ab16c2e652a95dd1994ecf807;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74cd24e90f61663096e65cfe1ef4da16695ae1c4579ee614958db50481b71be03eb0d432b2b6cff92a66d0f455b816369a31868746973f865f8d445e01521fc549d7087ab8262a2572a2955244402c19d0d332649905684c8a462fb4d32e135e061fee075fe2b62cdca14958ce3f8b9f1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6dea922f62adad1852fea97e1c1834812bcfa85bba9c3647e8376a691809767a9e6cf825b9000ca8db97ebf8058304a1facd37cdea14a08fe95b73d6cbf43e2acee531d35c3caaf725c3784cd50855338eb8252f0658b9fd2f1bac98254ca68afe8ba85afb817bba09fb13ad5914f40e3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf5d64f382f2680c4d9728ca77efc45370917327a0ef66e714a70d8f0fa507802f70fe684d64db60f28640ed62cadd00a3fd4ef8d59655c681dd5e342b972a84ab8fc7b1c51bcd4a4fd5dcf33d6709a35a035c5c595fbbccfbe39dea82f85f183a80ca1eaa0b4a8b830ff59d7913c78f45;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf90bc7d7de712a47b7dae8faeb2b4a21c6c6b2a33aedee5b7883389baaa32b7478da5785844af24660ec5f6b4a29752863708a107dc0a234075a622113621827900c890808d61c101b707e05acf6c024a2e9f905e77c316975a8cad3e20e363f28301c643e2f15063659264655871242d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50a3fe0a75c8cfe3f018648a371ecebf97b698157c05e6ada0bacea8f48a0c3ea5a70217063f66bef01c6299ef20953d30833ddbce303d7bf986c010d37f6d5dd196824587b28fde4509258520a5b1bdeda5e50e63f54a297c0f31bf77d7f541fb8c1eae4dcbc53441ca75bc68691309e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h16d835710bf5798843b002bb3738f8e55f8f834bfc063848f82dc7d49668571ef185b39aba10547bb3d27b75102bee66765229f2fe253dd7234d5d29faa7e4d0795262d3c7649fc8f05299b0de8990d1d61fac3ec4d450bd515413bb9608e3e573a898545bbd34da51951e8e4f7ebc5c2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc659c21c10279ba26a1572403e8e17ede934317f1cf5bb1fc4f48a6d41cc93ec5d0764eeffbe057b94f24b9d6c709acd373f7ca3d14477cb0ab430147547818628db3c76ccd678607ae016c84f5fe1abf48bb55c7551d85252cef08b9c3f38ba4b0d88e6dda773cc67d3585ade073bda;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5ee240eb5fa06dba6973b4b4d063c821e814799797484da17d22f655902bcd39d3fa684727956e0912c7e0c1a38fcdb8e09aaa82bcf27269f04ec1e9d8760d377ac70d83289315c1419345068a6c3160aad43a995c6d33752ca18b1b4fc8ea274bcc045b8c2aa0fe69253ca486186135;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f66b100391dbca917c47c4ab98d6f31037e076e87c350bb3da380003ce75826bbb17ebbbc924080652e98d8872a35e030cf584d3a4a418a3cb065790639e85fca308550135043270b32d9fb448f6d73b2f40f2053c517f8813e8968c5b93eedd93649fcd29007c834ff3274b7e216ba3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1170b7394954d3dd3e1c9d3e15d2313a5754a7d99914a3604c942653e53fe833705f19e5293cd6ef5c776fd06871443d22c3902c09339544b7d60ee4e2cb825b25e3678138f6b0070418a83fd408d7eaa9ff3b82ff459e26457df8b970c5569e36c730dfed9137c9d2eaf4ea092fcabe3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h766a680c9337dd2c7e4adef637f3964fb9bc3030591a29e0504ce7e4e785b9b6dd2728f2c4a1fb5bdd21b390ff8cd81e7d250efe9e30ce57f359e00f4b77c987c94f5ca4f70fe324cfbdbeed1da0f32e1007e135c89adfa848c178e4014761ba33ab41b26e89231f3bb426011b9938366;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e4c7942773e4eb925b7555caa46a3a12df9a701f39f6c174627299d689853d2e407f02326d96b905621925fb459e41465a8d54d22500df08d44c9f5efc2db9e80f4badde6413f5f107b155883ed774ee5bb2e0ad6f8e25abfefc4e5c3e4b7bcebde4accc427163e64c7da81feb8f4527;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f9a7b5977fe390c8530cbab83b7ad957d6df47a60226554737528cc014b4871767a0c012c5ec5c16337023832987b1015f4ce5f3caa64793031c8263e7e6c9e7a6841b5dba3387e3296c8264f777fb85951591fc8b7937d4c11cd3222de187330b9d999e836997df85381b6e9641b11a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h431a5239c356fc59f4b6be783d167b11417c7bfdd067f8a7ae7bd02b67e6bf3c31efaaa344f114dbf66ea691ea94cd6bc159d62c0c17115b4926003eebf46b0c3846d908915c1fd7894a5388faa1da74aa35dee6dcdd2b7f07d09f89e69770e8eeb993460d3358161cf5511bee5684d8f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c482bb1abd2affd295d00862e2f94408f1c8b3f9739ca0bc0ad24af143a8deb87fc6740be5778949c7ef7478285badcd89518517eb20b1abc3321aeda240ca438b82a6d12119f5b32c88a89ac1bace216c173b61a8c603527e66e4e3e9d31eadc453e900935f1af0d2d00035957587cb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h19e7e7c6098b07157e3c499566bd8f492bfda0690860511aae26ced249089de303370ac373943ca89a0d5634d8ac8bafcb52ef4e341c8d53af197cb40750181fbec49589004501ce3657e5865661067de8fceaccbd98c33b071cced62aa5851590a26dc7a71ec27724f854fa84872f33a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h291f8c726f84832f611c1045c1d10e8b3b840a912a8083f019bc9750c14817cc9fb03a9e0c515a162d21ca6ed546242f7f754ae15a686beef467143cb2296824dcd0465a3a5159cd5ad4986473a0337a18bbfefa8b0c0df6444ea508f8567384137cebf5ac302610188c386c36446b0ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd19629fbe745b07663eadc250cb1a67de5b05b37ebfb70328d9c476e6fb0da5f274bd46f9229f1b8505722aeb3a70b944c9255672f8ec9b1d350485183d5160f69fdb3abaa5cd2f4b78f3a8302b7c93dca5a1ebbde210823f2d8d1bddc0bc0759be64092e61ee566c34b8020d10d78f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc221e51f1b67ed36d6cf4810a7cd78926d74021436f95fb2a59118edbcb9e39d7c11e3a3c1402b8c324d133361d43c309a798453913bca43482957aeefd8f3ec121832f856318d2b351f19b87153d86d602a38eca478b45261d6b5cf5523848f5c29c44b3ee56d505f9052993badc611d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf3477237fac152242a8e77dd356d6d333fe9eb3776e6eb28b39cd03ec77dd24c31280a704e17fe0e638ffcf78fa969f575b360e6fe32f3357ec4f107d5d8bcba4af15de4202f7d795c73b72436d79ad2f74582954dddebaee1f2d2b782ef2581324dacf337ddc00034a6dfa19d7682f16;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25b5e37df513b6fc246aa0e3194d2ff108c71fecce56394edbe0f515260c924dbc0de5fa1c8b5cb17b79805477494e33b4302a800efbfdc980b77fb4627601dc9cad1561a7d92fcf1ddc8f52f186e613e437451d6a8775851b3aba944dc3d54296d647abcbd869b28c630677bed8f7f69;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcadaa04aa96c42c668a1d6d7a57d052d2bff236c859d6c11d079b0c1d532c8078f273952ba908eff15185f6c8d9e07d5a62e81b8179c0dce3c50e230f9c5ddad75b3125b20d73863183c84be10ef7f599b4cab3bfc17871bd3fc2d79279eb791b3b9edafd60c0fc5f5bb2e894d3424367;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14b4b45953c580628cc6b3c1e61232c63b125da1f75f8e53936c14c871f07cdcd5874c927e4b004698719f5049bbaaa72c3c706be53bba8fe8325047779fb674630c1265a31c67f2eb59dd8368cac950dcce661d1b88e0b674cc989871aad555bd41319ca25208a2cd320e9a8412498a3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c38df5298d7a9f76532649ae500f4c9eec5b37a4d21d8b6467049c92418d27dcdc340bc9205e1c62a249c9fe19461cf8cf533c2ad113038d751787e7d4423f04499f1a5bfb73667e1833ebc8c7b83c822e38b72f7f5724805f7af2434bbd20e3f047bdce1faa6ddb6dd4e26aac26dd3e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd385d8b29b622856739bf3b45ca8cf875f5ec2a9b9384361d12ef2412c6527a6b2c638307c3a4ddabb615f732c8f6047e6d604f36c6d48cf45754d9fbd60ce68b3291060ed8faac8839a1a4a8b785566970bd4e7db9def15483b02d0bc733cc5c29aab71b0131120c38914476f620a58;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdefe650ac7379886edf6c3bfa6863c1c9df81ab061313813ecc0c8f2d642756957f40b4a3ab149be061e751e44ece88ae9e09cc42bc6139cc08153716ffa66d1941823387201d777dc450c08e37629f189f2fb09377a2142dc01bb4a46547686b5f904a658dce03ffa642e6f1caad30c2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69f323af8557b021b78a1218fbd2fb2fd9a5d748c7fd8bc6103649e848ea9d54d8b74ae2506183f5cde004b9a7df026eba535f8b1f5571ed83361de6e35d1a98992392a2663fbe2ebe764ebfb290363cd48360ea90f3ddbf3dc6b688595fa4dd3750e8800b5928630e1814083b1dcb216;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88f5794b6bf023532857578f3c0ded188c4f17c3b542c6ccd82e7b239d1b6df3e6c1263b8815bc1d6e91ba516817d266b6571cbed55e453181c349da471160dcc92ced421ae257828005bc8ad63c85418de8182bc791ec2042b9e63b8c51a5f12ded40e43cd5ede43560089abcbc8ee8f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h912f89883e959b186484e32f7d429d8b607277d627cafaf7bfb7a06913b5eb98d9afb674492cffed33b3bc8dd5f805a911b8d748231ab2472baa7a8c816e498643280d5a2b70e451a06c2b0fae77195e6fc8f40153d4e41e42f6832dc7c0881c10faba3cf2bd4ec2ee96ddd5dd7f8d7c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1c9a0114c1bb305265e1f76f01c94988734e52b22d2e48989e90a3633d18bfa52173ab555376bf2e3eae58389b4886b0435183c2556f56d121634eccbe5d028c5d8c8f01984800738297764c41b72c6c2a8f385bb71aa11479486c722aba81ba38ec7d216c0ef691e8e61991d0a450b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b59a8d47fcbc0ea742ba4bb2593add2f9a994d21da6d98dbd23a0c9aad8b3ea2e093a3aa499fc8659f15bb9d35554711ba181211e03a085f4f5d2a5bac26fed059e1ebacfc44b7c507fabde3d42eb2098af3222bb5790d321051096e68cb1963482cbedb9a214a2cde983838651fff7f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9089c5a1f3df0773a06823f4a70dc86d7999ec3c68dd0ab6fea83d3e38d0367431dd26ca14507f80e5ecf0e57a63f031bdc656153600b44b469ee6c6f8a81a5049f95dca97e5a884490e50a532dc945980397e6de0ffed19e46addf37ed68fb2a677dcce46cee3e602dbf26d32d78dae;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd496b3f14f636b8911f88e4d6a5888389882fc2780e583211b283f85537597c98fef89a710cc667c4280733006ee018bbcd424a771b570f232bb9187dd2242837bd40d30ab0d145b8337ffe257b8f686c4880b52db7440cced8acb2d72fb837fb0c0edd4add31c72e842fbfd69144e77f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha3ef4a999f20e1547a4430b5f607f19ca1741d18a3b029ef825e45d8d672eed1dd2cda1bd9c8ca1d49f1f308cf5eee40cd446683781d1fb9a1c7c42e561c2c3326d6fc3e6e9b6153575ae7d0ced8508d3cf3952c46deba407d9460c73941a601e8e072e3397b57f08ef51edd371fe0e5b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2df1a492220dd26f36f5fe359e5017303beeb2a30ddba8872c895c1e66669f176096ae9a46e20074047921cb504d5894bb810cd846ad5ee92302553016dcd236f4fd5cc3411eec96543c10d4c7dc000b3fa280c8009412c113aaacfe749a872958af0af1491204a318769be7c0decefa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he98284846daa164305527115c1a8f251f2faa508241295449ff2a7970e80c9fa8dc5f4026d4e8ba4ea9714625f67c0d0aa2bda8ee5ce237c457409889656a912eb4f3d28a34efb66642263677503dd1e82470addb9e3de432e3cda4eae41cb6fdfc82e43531ba556a2f153090eda5dd4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e54a17a2a0857fbd5aef89afcdf1b55042a5cc24ff91419be70d09b1896133a70af61dad8c655030c46e249fcfe6b1b6d97485dd9e66146cd953043f0cc75cf9f21f25426da3b5a52092f9351feb0cb1e2bbc4d132a8f15632f5547731f55771639b3ac593698110c98fcfa3628323f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee257030de497c94d19f0c4f64380825666cbbe11ff1a998145f6670693544cc0768e766e5757e0a7fe6eb59ade5f3b2367f0892feb6a4935c1877a363d703c5063d3b376b6be7764f1397f89360456fc18dc4da7d6f4a37997d80707d7f91b29a77f43a537907e3802f82a2352571ba8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b3f2ea26b4cdff4a51efa61f64f71bc8b4e485dc86cccaeed03ebd244bc9eaddb0fde933f2415c0bcde3360eec84bff557cbff80fd9647eba554b8395bd9606247988b8d25b0d536e24c3d6699fe990d0a833527ba6bae0709b09b5bd6a7d9b736e2c705ced0a7cfebb93ec976fde14f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h577aef3a8ce5c52563500fc0ea657a5c3e8f544136f2ed2134f869caacc12c81369a0c96f356281057fde73c3cdac2eb66494c8793673568e22b52f1d3fd5edc9a79096edc92d6613507deb029ecf983532038456ce9a31df1a4361de7460c78a4df3eba325f5a301d8d71d2a520af3b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha0e7d7bf73ade9adabd81e444a9eb89c26691b789b46b7a8a05b6c95d660a067d07bbb85a204df5ca09f4c7cbaf5b2ae28b75f99b5d276464ef89eaf0fe8cce66605ee220b5e23cfdfe05d5200ddde5b5a08cec019778808178b1c6a1d642e5e8a6bb2a49b1c0abc3ab7bbd5c3dc8f254;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfac828581d6e25c131fd6823c1692079aa157c314ebf1e04681b8a52726b04e79b2d7a0703b17289e705e402f8efddcac948b1c96782d9d860a328f29b9c40cb43bb9f29017d6255587b2ce0c73056fff649cc3827ee3c4967c04b07869c048962065b5e2869d6aa5b8c7b483f0aee764;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb1e6c777bbd0db21b91b40a9bb5ea421cd85bd1095066531a15ed6818c1bb22512b42c3d2b0555a5693dd2d87882c16b424fe31a093dbf59e04ef100366fa70a593d59ecbfd2f17489eee5b1b09b286a536327967414a15202272fb4f6d6595a5ad8eb75d24b34b5b60569a872499350;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb1fad801ae03e10ca99bbc70522d9026bf2c8f4f99b35ef64ba1b0a4d7bcf562ecd4dd99be8952840e7140858ef7b8dfd50ab4b9281d0d0cb66287ae4929445425cb4ab8446d52a7b26cd4f15b101584e095567328d0369d9c4d71b374f1284fd52b956be97538e3ac6d7364f71d84e3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff9f9ee2e5f7a830e7fb76a515ca0543c1a54ee77531f40b4f80a91f62eba7cfef0bf98ca4464d98bb664be093b8efceebef8ffc7893bb421bc39d042139e56244da1c8591dcb6f3447d9e10cbb6488f00b5ce313b0cecc3842e61703361b81a3f5e3b9f5e22d3ccc7ad570016b0ca88b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fb97926901c577966be86577a68a30db2654633869fc4c219b02fe07d8b99ee0f43b8a151e2dca36222f4361c30ed8d27bf38b6ce3a7a9b38d302e547d101d96fe345d9e5188b630e8cd16271882125daae72bc2d307a175aaa27aea944c39bdad9ebc9d4bf77a925b5794f3000f3372;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e3d5088738f866e36211e89bea72e15c59a473df7f4bdd3d8d3850ac98769876653f10c0fa52abf3efc633053f562754450501d913f74017d3f169457cf0359f858b470ecdeb2f670ac220d1bd4940b32b6427ef05fe5df7af240166593eecd9c823df4e0be5cbacdfb1e6bd650fbfaa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h691c3cfc096e8f456710a7743a7ab47d2e04e1b37249ecee7ec0489f82ec56f9642713b1e1bd3c0b94951dce96ee282a6af7e30ddea68e2e2fecd0b11336f12f29c996ab7ad1c6ad001c0efc9e042cdfb4a2f4821da8a4ae7a62d23aea575d163e91297f946397367ddd74b8cb42cc68;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f62f402654cb51a83d1dbe1ec9357c48cb08b4749b9ada94831ac3a08b83270f95dde47f8cc7cb377d9de0845b7857bed1ea8cba56109d08b0815f586831c4d54a615a0d8dc33ae86a56dd639f1c0370f8672143a884614a1d574568e543689e07fba17fa41daa4f0bdbc69850cae5ec;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2bbeef09018ffee082fafdf2f7fbf2919c5f289155e9f6f4b4ea1919d1a07dfe1735994172864e1c857e42d4453c1389ceafb69c915a98635058b3ea3ec90d9fe6ba91b2a66fa4bf0762703df17b0a9dc3c989a329e4187379ab7b4d2388f6f5c48a80b843236def2461e316e6db1456d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4121407f355b1a342b77ae33f20349102ee45325f62fa458ef4a364eb6705028fdfc0e5467acb7118013475b7ae1f98a77dcb3252cccce94e3c260745d144fa8bc56a42252f21efcaf913377ebe4bf7fc6cf728398a35feef5206ff4ebfacf7247ff10974684d04882dbfab8f3426b59;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5cbf648a7834976f138e7fca15499dca84f01bbba16073542a10938b7fd77c9941a0bb05d23df9dd70e39b5dccc00e0ad1429e8b5f8c8dbf04921a40b6fea8087b25696fdc443beddff985fbe4851efd67ee469f10d4e66a48a99eca93333d503ef8050a28b0c6e4ad8201a327342cc1e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1a9bd6aeeb60b592102a777682761dc65cea077a43dcdc377671aa045fac24d3e5b71e674d03f882bfcd8a4d020af206cabf821fd16f1187e40d4dc546c31a8894b9383198e462a5371fd9ae9c6e3f6dea66eb90fda9f3f9b3e2b9030ac49d8f1bc1b3aabfc032d1aac455ab032dc31fa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf72bbed3ad6bd20a6c83dce6a554a38eb6558b9e6abec3feb901af1eb94d6030f8634d7e487f2f4c1d88de64fb58142ae6bfedd88153a89a93f7910945608f220444be391c6d3d48d0cec2e50f20100d13309ba412c35255d271d34b6047b71084d81ddd13b2794b21a4f776442b0a7a6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75c01da28bc62512c7b12563e03f6a8eb31b714b9b7ea3a76e2377f429cd3d4bc0fdbcaac15eec8c8abc02d133f032583f4e8bba9956ba36ab304dd439ee27a61dff56763f89280bf9cc9f6d4e12cd7c3423045a7ad27bf34fcc98fa9dec5355c6f762709d5647172c208d4acf3582154;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc31537666e2174bb560602787259d07e2b66dd455cbad12feed314e3da4aa0bb712126a1df4d9c8d167fe7cc57de6315cc6c6aa0cf5dc923ee2df88adc943c61d2760d47fd1b1f708d57a72ecfb94460bbef484e020b833f706802e5ceccb595024706cec6d872b3543d6943d390faabf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59b830bc32e2db24b3db8218b20a913effffe23394d9dec86fc20c315d57f9b22ee10523626a4a8b6fcc3ab3611d9ce1ed8fe4b6c66aa2ec0b64006ff4acd8b8b86481bb241be85c4b85cae1c6147af83c69532190037eb60c99e6502670725bd06316946764f544f8d2c5963627a8780;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h82aacae85e7bc427c7ed02bc65ab7a65591c96007c1818ff3d5340d4ea3869807110bd065d14a6323002e989f34725f1f900fa15e866438e9dda8fbcfb405ec2129460bdb6b9c2eaf6fcbdaae3d03853a8eca5dfb45e9ca77628c4a0e53241cb8bfe275f6f277763c9c1dc442065921ef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70814abc530af26fdead01c4b267f51ae46a0d1453d56504ff3fe93716daf31df2d4f52b0c7e0ac93ca2ffbc61b3c2ee84c494e6240d9edf14c4e9c728939eec6ba97bfb5c4eba6d61690be373620028924ca1940cac30bffa0a0a4bdb3589fd2004210ecba88049ba8b7d7576e457aa0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90f6fc1d5aed59fb60c194ea24a78ad3331f93cb1791c9360632de7175296e621c3ac77adf457619e3474c6cb05bacb1f778d001523a56ae37a7aa61839f4bb92669b3c473297a57e2c38c4d456148e139b094e3b46838396c06e48a9f82a0690cd0d559f344fdf028fd94bca70735635;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd828c1515d1739a8ad7bb22d736a1615376aec21c0804603f587243a56a267d1e100480d2739709dcb7fe2063ea8ab6844e6982e750fcc99662e4d65bc3031cffb19153192305df74fcc250a2d79e6042efd7e067142c7c620f219f97d0ec027665c9bed4cb3f7c8063a3e9e144afe98;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd91a4baccf301d6a67c125e215fa37b494ddea2fb313c53b6c18eaec0545dc63ddf71406f9a95a78cf76f69e586080c48efca622614a69a32922d41df25e9348627dd8c10246980cf66f9bfc0a47776a901e201fbd7431412e080105d2638ba370cea0f2f4060fcce86620394e46e73a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1c3529598b55ed5be4368143a0efdfacad75a6194359efd064419cee351583458d985559d81c1a1cbd84209a691fd109bd4f5061b763a0186aec81b9702250cf4beb2e47661af204c6f37b31d789e576ffacd8e6ceacd56fe93f97281e967be61fc7d9e8cbf43c1a7df8aa456e22c764;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c6384bebd0dfa21138c4c99d151a9643a2c19abe89ff85bea8802996b48a2c098a6a69f008fd39dd605fd045aeaae21fc790475e5dae7779645720aa77316dd119c952f8be395cbcf1529707b66393935bb9f14ef3587b6b6df7067324c9f0bbba1455f9e2d089e425583a43f80bea0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7cb5c8b784fc6dd8ad7b012d13a6f1273c7e5d282af42936ecb9a8c9bfa51c6790e3cb08fb6932478f0baecdc0ab61779757450cc1b3fea3d036d074abd15be2ecd1347ec26c11fc1094576d96298927f2b37d214e7d23ae90630231324946482e7e17f82716152f2da60f0ea870574a5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h964192efe3c1fa548322a83149f007243581bf1202b3f92eec9bd71c8dd2cb2efd8a99fb8ad89bee1292cbffe0a42964687277669f7e2f71af7990c47efc51bbe8b77b2cedbe61207051093b24b511c355f30148e1362ecbd1c3a885006d8a01222b9e188561d82202ae4d12db7eb5bb7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2507c0e4d24008823402f8c3b421309a39b60abd76a3e0e4336264b5b3dbed5961a8f8de9f26013714aacc06aa0e7d74a583c80ce3396250d52deef27d8985365cd9d172a2c1765387f701cfadb6bcb89aa83627d96ad2cbd84cee1e906df7784566c623bbfb6cacfaff890013631b703;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h40d0e84be9c6936d909b0377db4b9513130cf066a20238c34ce9127abceb5dd82937731b25b02f3465a10d7d3722c68887358a2a483a04dd2b9546f5356ebfe670288a760f24bd4ef24a196852fb894279b6fa597f955705238de52e5fe0be2d410faf43ef9708b80a980d4328e97fb7d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85e9443952a74e4556a45864e949a7ab43e0a049a61ef006fa488ba7207197d7e26401cab950e6d0bed24a9027cf26b590d1190f95e205ae121cec27f2837125df403e2205750d72e4f579099ba592248726767b8ff4ca793608652c96173f6e13163991363a5adf64c9dd16a0c45b4eb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha287e590ffec54dc19a2fb23bc0c34a123742d343a2d973ec1ec6b7717f88148eeead701382d64d5e1a0a15bfb49ecb8268ac75dc4b553d1c7d8ac4a9faa7339918f1cc4cdaac6633a000a49db55fe26833b8863416f56b6596999ebeedcf93523d4589ad3f25a1ab22c25b5241563a89;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf666a08039282d2c931713b2bbd5268c4467494a1e1b57be482179b71b07b17162c0db7087090b2f24aba4751eef7d40001ef2d7068f74e9d1eaf804f013d226697d22c95094907572b2e77bb1788285c8dc5c38abb7863fa16bb81e25e38d144f704ac54db079648b9bc3424617fc7c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h65a8b4e283f546c776e652f7b5e8d9a1faab6854f0f2931d31525f91fa58b71c9005ddca07983aba2b2026b6bebadb17130456ff65aa3c5ffdb891ad97ebce98eac47748912a6499edeb04b553e9f8d01a7e527b7612edf08047fd778932dd3dc3a7e10f07437c036d360001d4bf4209f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8878deec9963fec075305671aa7634d9e1ce1394aac9687c30e3b5d985866aa0929adb78100ccf848afc689bc34f711374db2c7f8a6dcb6fc3f9073c0686163449fcf6d5858eef1cc3ebb76b8dd8515971ce1314a630bca6329f3e8507122ed8a963701d90e4bf150e6393f238d7dff30;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdce6c678302c58853e2c14a0a1ad8fe0e0c2e561164b75253044ff9abc0771ce71641d68a86d3cbe093768f83dd273dac6c7853f172827728bdd858a33807dc4d1cf02a82934f131c150133d92709f6a75160468d42697c9260c82cc192f02cd82a76512f0d0df2b0ce09620a38b2f5ad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h808cde579ace07c8c6e9d36ea92e3089f5325626ed41f6b8b0aa9a61a74cb3f530577d9cc5c9b44b26b9e1fd3551bb1c371f1b6bdedcee731664c6ede1656cf0a9ccf529e71bfb585b36184c835716dc5eebc270b694e1a4362217a00a4bfa0d851c41c03bae74086c14aacb2f1181f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha134c2c8f4a0d525693df1f63920f5be9f193887e1f25993c4f4cdede20bf291fe6ce0eabf24307e85ae5f08e59eac12cfb5eaccd188c0d55c5ea84a9a5069bb617c0f20db256732bf658b34dfa84bb7aeb3e06ac3698e2b8be91bc1e893b54bb7c1bafd7f92e15be8e6b19a2d1de5ba4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2cb05a4cf21b0a2a337e5143c4015795bf38b43bb0ea3e2a2160b4519674c8c04b4ef4f33df90dde3ec39d07831794f6a0c303bc15e022c04e44a4df591d8a7d5547a9dadc11774d8362ee16c37e462c3439d25c54a1745fe3340b83922d0e5cb04ac9cfdd536a54eacc963535c61c2b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0931c255c2598bd0290435c1a9f22f0c1d5944954f469830d758e38d4b4f2398f2d92ce7e3479b8cf587bf7b53db634c20ea8a3c10fbacb2546e598337426722bd20a14f8d1c13ac84d5819d266b9338d719ef34b7b2e4f398f6085fe62954ca0a0af87159c75127b61063d7ab558415;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69bf366aa93b4ecb3ab8cc8c497d26bba4ba3dfd7ca25dd35071bf9f904f8f9ebe1ca7c73974587a0023d66af45ee980181713f9d03a5605ffdd7ffab4272f2a70b5cae55f73580b81fa13733546a896344de46a5ceb6a983c7f235c874fccd099f710ff984afd391ffea1bea5631fb5e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37479a9996d563ab9bd33bf068de6e796aae963dbc302308ab7047017afe4b2add180d4fc31eceff746fa65c52c6fb82f529a9ed41ee0ddda6b1e8420a6a2ba32827fc98c96a1a39e902af3756e510ea74aa5e9c7c3aff2604b89522f73c210504fe552bf3f3487eb3f4d510b8d10b332;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hedb0cc2a0a2120d89b5a72942b2945c2dd23300db9514b8af1e223c3f9352d610d19bbc37b9b5a569b4634a4fddd6a14ccacb61baf28898a4bb9009e33eb460d835d3b0bce1c0bfb61c2ecfc2f78c719fee7f2f44a93943cd8060f764d5f52aa0a65552910a550a35db03df9bc9105adc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h604189ac46631e7592ff639434c60f042fb7720e21f34f023375f3ed46ad274a98ffd24f83842cbb6d91294d4d636f91abb5a8fe27eb75261e9143dc3c8587154d75033b34e0124f3012748243a0eb2caebe25a17a7290d328820956c1c2b85957432bcb48a841f13ca2a44152f90def9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81374f3f5021c27f4e7d699558ec8bc6f91f656970083f39cb8979067b7784a4ae1036c996ab743856e869d4531a4330bccde2236956fd1afc55b4af572873a5c429a92217f63320508b7c17e5b7694e8dcb11b00673a7bcf70044558b87d9e63aa30f9569a0a0843ac57905a2752ba18;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d9944001e7fa13ec9806cddd457ee659bfb9eebd8b32989e63d125baa7b72a2d7ef35844a6eae576cc89d2b696cf743f376b40010792283fc3cde0bbf52f6141b079c05a3de74b797ef09471528ead3d946727070115c03c57f50f83b759936fe3acbc0ee0b5016e48efeeb464d3e003;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f8d519ff36b86fa04e6518396ea95f2cf083adff0efdc1ee5845aaecc64771a85cc2b635d9da8ee7c5198f9f0d4585779a21623d0e797c31ba6d7f006eb7834e3a91c670c95162e6cd5ee30349c26310c14c37060166b437b7e9bafbdde4e254cbeec87c456d9633b601c6555ba01650;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca9c487fcfca4afb8c48a67affcb7df99eb1e2b32251a336d2b72c5428529f4d821301d49e2c2154be9c26ae41d0270db87b50b6d40b5509ac872ef3dd41b2be78d85cb02f49a91170c86e53d9cf3470cb8850d481ba88517d7730a70d27ade11cc43d234631f6a0d93385e8f952cdb3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdb07b093e0831f09541ace3bdc164249bd521ba9032b4ec726cbf37eb4aae2221ee5f4fb0f0e7fc306735d54864ab97a18b2b05ee15cd80a48bb69cc8c1bb93d0ba05573ca69da5107efd600f9831ff07e75a7de7ad42ffb8f5dad69d7253de3c31a9719f0ff5bdc9dfbef87559fc39df;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb15cfc1b449210affb4cbd132739396914c72abb83589acb3d89d7574f085c1ef0521f3a6922b1d33417ec6ec377d8a2c48d2bef93e46199fe856bb8ac9657e3a0fa0ad64b907e2e2fca5ffbb0a18b2c90c2e95f3086b24101917e1fa26cfaead6dd5cd83e345698f230c53115aa0979e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7599433be01cc24dcb67f4f60d55e466db5e5659c05b55253e3f71141c1497a96680b6219eae2afc8758fe4e3e7db442446a7f63f26e23975c6974dc4f597bdac183d30154d56dc13f493b715f39b602455c4b8276da8a25dcdc89b1aace24e8ce06c6a4d85aee68cd1f1790d005dbf6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h182ad82cc334d22cec1a2c0badae3b7413a853b64b1c34ff346fb283e3e14e2d70b174fdf32eaa15e9a747efa520317a34fc1c8c47b30105cd5b31f00f0bcf7df1250ae4fd463e43c3ae878b5804f5171574885463b776200d2e0390090f6ca6ab9538feafec353b6fa7c6a173889f74e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1109a9ae5ce985df898b3cc845b382859ea80c41e249e3c378a8729ab1381181c96b4d7c6d88d657bd24f0a013e999c34db1b7341e7a57d9a6c35bfba90d50e1b33fea86b6e25679137c17763af93ca4c27f1e4cc79ee356f794eab706762d32623fc3b4c5e7f2751fb6eebb57a8e7f31;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55fd5612a444831685e5176431f3026a05350c20514b327b2a79f402e97cc3876196e3d0848be519281b5a5d67bfbc5770a92b14fcdcc9426599f4dd238c5b860df4f14c6fae21fef39742ef4b96024980178d6e394ca5a616864bf90cac8f060d4866816502839e2957a1b69b68515be;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4feb5fdfc49108d732d2ab85079d790d2480cc5af6fdfabdda350997a0a16e5e29cc723f59c8b9d02fd62a6e907b8066c437b001f0c2ebcc6203509cc4fb2c2be2a67d8b29113929894db94c41e806ddf2718716f3266b4933b006f9e2213bc20bdc69e7be7e565d1e3d7eeb540e8224c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d890b29dae94bf034e97fc38c54562f3112a58561a18ca852bdad8153b9d8500fed2bcff215df91d88d1a82279cf55aa10fcd7e21765924444df5b0a071cc6a77c7c03385df3d0878d61546aafbc48b1320198e939ae843ce2132633bc2d1015009e93a5a82929a8d0c882ba993c6c32;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8ccaf8d55244164c514239265838c9a90eaf2b38ec9cc9be105c20164b393c6f1e3461f6d80cd8ca225df5a3aabff3cc8cce46e1628cc22e42efc4bba91129b73601a171061570dd1876b20abcc6fc10c199cd76158158b5ef5480cac766a9090573eba72b7b47efaabdb77960d165c4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57f1fac2b4cc87e3eccf78f39f531b7a1d2478152354d320b839b5ce5a6238b66bcb1a9009f6ce6b9e367f0d116858acd82d66e040477a8a8e419477e0708f84d77db9c5d546febfbc45738c27ac786f9be9336752d015c6e25e46b4cf4afd148b5f3dc88501d368fd9f103bc07377ac9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c7cf41a981f276588e7dfa8a13794b88c39ccbcddb630c8e29f15739745eec78f3b88e9de5d9aa79d4b8ec090fb2525da02fb584eb9eb06471783c727ea59bbb2ecaaf4de6cfd0cd315c55a5c1b4d2b0660873769ce083ae81741e7d7f4b12c99e2c4d58858ab31de457332b1ce8bbd3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5fb737095cde99276cab18f6832087da6530dad734ba07cc10c9e3ec2095363ae1556d40f7d804aba9533732d385fee29751d897008c5c09bd00b7a10b866899051c8de72251eba42fc15771a44b80bbb862d0b3a5cecfb092e1e0e79bba9d1bf0e018b6f35ae9b552b04bc548f2f746f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3081b9eafcee4179e6617a0845f4774f38855399ce2e230445bbd8c1141bead860f7a7d493f839aa89d6cddabf20f3c7ab584a5cbc48918f0a6bbd31b6ab999d4c837f059156f197b2b401c88427d08a443f1bf84b4167457306ef50caee4982378cf6bc28a55d238ae5ac63d1a1b5a2c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h81d8a26d0047a682e4232530aa3f16820b2b94dea72207bc1f2589c7eb02847b0bc664ea19bb24d398533052eb73c21a8b4d15afc57017ea0853fd110bc77ddf0a3b30c83f5ca8182c94ed23fd6615274f2165ad992e52f2ac125ac9d24982ee2041512608c87ec7a8f896cfbc240511d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h60271aa2ca83d0d76c8a164af1e3aef54c41d9b849d0de000f0596930efc15db46d933a03e0616b7f9170dd9fe341356c554930174a73ebc24a9a00f788ceccd15be5cd47910994f3f4016ccf312cd22829c877559c46a69a0b6e735cb911322db1ebb1e7356fa65aa3643587c50e1450;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h973807591595c707cd34b4c604bf749171d810752533044e025462fa3068efc778deab968c4c38ae6f527f7be261957d86af9351e42f345248994be03bd65aff89024d58094e641e5afdc952bc79488bfaf70653c0deebe4e52a0c7a097b9a53ee9fd18957e6a09fb478a717acf9f68f1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91ffc793e9d8270090316cb507702df79113a6df0a75b058be4d53d65d378e0092969ab2cf4f705d2a42d4f999dfa45cd01496740f32e5b8f3eb80daf20f9009a69e6f900b090859a3093c51cd49cb2a6f0fac32d6c67d243fd0ba91dce1d904da830bb6fcc756b7b1d120bb8295582a1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96ca26f47d0eaf93400223ac061db162a16e4b285dcdb9a89c9be80a3dda6befe761e3bf010c95224c95660ea0244feaa43530b7d6341fc7b6c2836e6d901ae9e6d277514d10e4cb34ddf1e2c3c132ee3c18ec1b10e9d9307c3fed1ca2468bfc9949dec5da3a10a26f4f7bc058ab92975;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11c1a084b4f02d25b95c7433cbd2edbb4a395a98d0f41b656f8dd91dea4eac25af05659de12045fad335536d272122ba4872985f01e033b0eb64bc04915ad16e37c2b5af81a03fb8f0d93587c62d780d510d9b26c89a98846f0214bfbd580bc2cecbbb0a75d22b65002e8d5ac49eb517c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf862f01732101852d6722277df67f62af52e3b962a2dde0c0de5387d0aecbde47e37e86832cee69f02497d41331e801abc850d8e608eb424a7f720df752003dd37ba60f184e1b967f2123ce83e17e57ef63e35e6daca0f3224f089ba0c3829658f9460fe3ed7b618dcf8f4fd015c9157a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6943e88017b5815019276b2ac472a73fac690e7947721e1b93291206d7b3103a35b56169e7b62ceb64997373a7e38144fd694ed9e5a9377a15e36866088356a2fa1fb9f837946f99e4020910fec6e4898abaab79b22c54e0203c6d9ab7a224704ac821834cf73fa817d4addd7ffa8f24b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47e80c01eb9c58cd49698e97ae9cac3da6d06292979b0a78ce71dd1ad93aa77ec48a03caae32e606fe34f067c545f705e28943c6958619cf5498d5197f0a435950c5650d5aee446cc73ef349dba661cbebb30649b9f2c365177888e24cb9d756508bce1aad9c62f1d2367019b09559084;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcf4c8417dfb7ffccf8d051df9ece1466761ca20faa13fc985908c3938baa6a17023e2c2c6b2b7502a200d93727210e654398085fa0017b6a087a8a6414c0f7e7441e72493e527f03537fb6eec9c09abc20bad0b7b9a8f505f329700f6ea8833691e466551c3efc4fe8f2cc66f3ce92c69;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2044c6af5f25a21150ffaa915e9b25a15e3bf1f0ac055b6bcd55f2bb96a955089d4a6ce6efc7cce007a7546d93343b74afcff79970d9213fea81f878f26021be2684fdea6d708da292ad3a24d34b5cdc019e74cb89d09c61d3b9e8fec400f1454f5896b2969673b55d7bdf0daf7fd805;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1bdd555730cea43be06879740f48dae06c9e9ff5c0007c079b9bbf0bd66f1c8eaa54d688871ac9f793b4ddfb66836dbbd62033c391cc8accf2334e4b33e67c3d8a7da3c07a75260febf813f116408322367b4572e2bfd3442a537dba89808fcf8eb385efda556fe20d8373cfde88c7eb1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30e9b8fd56919fac5867baab2e57cabf62d6ee1d73beb14e27e1d97e47815c53551eca09729d0e740ef6a264d3acf9426a8c65945b1923e87d71f1e8e6c833014ddd84ad6c2f13c59d4753856b74a17a3eebf25959cbf7f3d82dea93080a7b3a498bc68e6141032c087bd0435f7c3b91a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha53db4994e9e45c4d3d9e1fd71b5ac9695e56466465f58d9a5eac3746c6a44d453d6be4cd151321b83716ba99daabfe2570ccd18ad929360b26873da1512d38078117af8d27d6ad29fb84d22e9b12ee7f34d560cb89368deb9607db4d18102bf791a9ff1be35695e64076675b56301839;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1cd2b95e3544ec04ef4a4b3b76eab9273fc317cf4046e2cf26acb8f837b08a98bc98db8167088b5f7260890b79cfbac141af0d6bc299a7d546c8ad16f253c2ee1ba1795d3d057e24bb88395e1a8e8bfa724d1103d1586aae1755c928e703c168531afa4a0836af5a41a7d38c161e8482;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47a8ce2d10f96b6369c73ff599be1d4ffeb9fa01ffe5f07763afb2d486c0c7578e9d5be436a83d4a7e0cc56fc157e5148052ded68b4e381f23fe9113445ae7e419a5c9c4a04b2ae97e51d1c0521c9a61f50962051af06cdf02fd6c66aef92ff1cb990f1a0965f315a8fc36bf01775972e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6527e0f6bb8e5e5f0295a799de82c14c0723fa17d2c062127346d44e4af14017a011ce1560e9603d00e8c5c6d9390654863db827afae3db8a8b7b5156d034c9d2d04ffd89f205d90fb98948d73b4c751dae50abbec5417cde8c6bc23cafb15e750513db30ec43c07ebf1e4edeb79b6fe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb5c9ec6a91a9d65d64b39d720ecc64abb17d5aef47a807a1f27e1bcbcc276d2ff292bcd82a8c74759b911efff0834e8704a89d7067d69a616782e7cad8866a9eb194d374bb2295fed03a0cc6b0b1465f339ce3169bdbdb61f936456011ec4b494e29e37e98a76e50173815bca6c6e3456;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h964dce11f337da19956dac71e79b015725b3b4cf8f86c2221e085d145a1cf707e4c2a1358d1f8b1d8a6a6b4189a5c808bc0e4f13d63af56cc5a35963c54f6efd01bceefcbf1422264a69d380cedc2d0937db59095842f2ca1b22a18e771f5c2a6e21afc21e41a1a3f1cba829a8e795977;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1ee7ef9daa16c7f3978f8689d3da3e913f436a8a7e022e9bc7e37661a1f696ca77daec59e211efb773830d5072e332217c9f37a69f440660277d1a20df67d571d9ccd9d66c3b179038c22a03cc6e33f730e21c6e401c98070d3ff920642357212cb35dfd8de2542a0f1ac247404991d25;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hecf04e7100697de13abc8c007a2ced6b75ad757399b744dc83f6ddcb5dd589af4344b43d28f46475c21e3184e663d144f47f50eb282716ff28a7bee7129d788e2bbd5f7e86638b306eed64b282e3ab913c5297a9645d0a81f12a44302e71de4aa39ebf0b3dd392e51fa284cc095912f52;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ea80b3baf99081cc0fafc65d3c42e78adaf5817ce3ccd9e66db80ea28cedca4310a2ea5d812a57a6f567462c6db1fde6111051e5de9f355730cc389607cac7e93ea40ac989979591843b4fc7921e98b0d66395f714cccc358f87f60701b51db8cfee79868ae9fa71308ab9b0140ec82;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb834e019a2c8fb214d7dfa582c4041c9462723184cf3f95f31c3e40354c052d22c4dfcd769cac8b2a5e1a7dcbf457276f5536cc5c4598d4708fb124a575d535773b5c2555bb93c6c39186420900a5abf5549aeda8995fbb212b6c4b1e4c5ed2685da8aca7ae8dcae542773ed4a63a5b19;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb5aa203672abc7e4eb882c2e4cddde76251cd78b0d21145cc48ab9446090d7afde2c965d5e0765ed3db9b70c9a2627d817cea5758eb3e3ad3ff30f5cd6f173f345bef20d2a3224d2fb9df4830784baa6b80b1b78096d8df8304280bd273740b76e200e992bca63eb782450a68ae22a65;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he9dfbf1868cbf84b677ee7189054f5d0178b31176efd148ed30e3215e0be841ffc07cf66886a7b6babc1c487cd4e64707f27a8eef8edee71d15104ad45b0324f8d6fb9130524315036ee702629b44a4ab5086487f445a4c7ef311bcae2a95c9089f8d93896a53ca36899d8f8424161425;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h98a583dc4949d44b91af1fe5e9c8f65120be0c76fedbe7745a4e90946f8051beb31d35416f7274afe8369d7d5c1bad7aa75e8c35b4bf5bb8cb7bbe2d9bbd810b6f12acf164047405d06527947bba891a38d0d139bd0c0be017044e84b1007c9af5dae6d9e17a268f6478ae19c8b2f34f1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h594cac82a31b913869ce9777f8723af3a7a025c98c0cb5650a449d1a240fb6f91cd4c59fab0976eb4ecb60003b69a62836f94292450e5df1375070b019cd3fc33643bd7c599c9aaa275d724cba452e255af6d7dc9f9bc96d39f93b1c35b60ece0ac41b09cbd48764926647b171206d125;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec9c309969a498dd73ab49e562df9d2b6e6624ce87b9941b44ba6f0d31bb0d3685992369d50290dc02b242f9b6f885a164295c593ffe4701739c4ad57fdc1316bdfa2ed85bc596899d5cf675a96605fb70cdd28e495206f45f104a0baa13d4c264305f3972bebed8afa873f5adf60d2c9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd63eec86102209271e7571ae21cc02b416b915b6dd566379677728e1fdb7f22381dfd5f513a14dbd353275fc0834360051e76823ee61bf0e33bfa47e7fc019cfa65e62207cc0ab7026e7528e9bab53d594d11b113d86897354764802339b5ea125871f70518e6c7096187f3048499350;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he826b174c71988c4cab53ba14952a1014b71040c6354d71f2aa0521634ebaf611bff87db0cf8b6de6d9a2a94427d9b0b62819f3b321373ddc5d7c625f215c2d82e90bb968c79e992940899cd9094a84523b06d3b8f7c5d0593c0ad571ec793c449daee6083327284933751cda1f2b6491;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he07103363f34a147dd9777817cb3f70f842c4f0545098a055cced4e267153a8fe50ac373565cdfa03848fd3d3dcb8e1dd95b7236b1caac8e829c49bfaadffa258a4364c927713abdf1621d2fb6e79156f62faa37d7e7a89bc792ea51fbd4a15a85a254f8f71a67c639de45ba8567acaea;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hef45b84adc5ba0f8327382553652621989c211ee943a444d9a6dc5119826b7c1b11ddac292dde0f7f81a1ba98c7b7fb28b7fe62d5c5ef724abfdb217a0ccf278c862209adf092d562c3f9b7feca1fa57b48aec2a02c835f6e62b6744074abc7a9675d1e18cdef026a12489ce7b0ea35e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e9c6ad61442567fedb5343344006d95ff487a1b4c7c4909c51cf849323707a7e899a3d5e6bc0cce831fd0b360dcb6698129beebf4bd7a17e136b10eb679f3d0fef3cbb43d7561b6f2cef911d27016479983074722365f0b1707965b7ed7d0d134247f347c030287ff44a747f0c8d8054;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2062ad35bee7e7c0fac6f2a94bd244f0729ec9147f055ae5c95c450192d37d63c1b2fe0170e06fe1b70d071a8e8d2e60a7b6dd85cc94c2dc62dab73e559ba2f89dd007eebc8c685bbef3d6530af4295a530205b7149d12e305d5cd265e347f4f6d28b04bfb18a288174048728d2a3c174;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h377ee4b9122abfdea35390994b20f0aa69a6a1e137ae1e831f1181566134ae6367d921e0c25289a15e2d23fc9fc66d7205b92d37a82c60ccdaa6221848b256782b6c3c047792d2fc3feec594ba442e174c9fe362af0a941b57159b113f06db74228cdbd0c0d04c62fe7259d307c164903;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h972e4f3c019acd228246ce237a0683c6ae2576801d4a15f8cad54c4bc3f335b92c9ba05bd44dedafc033da365f93512035f9b60091a1533a923c3600ad23b5515d8f861d8da7261b03de35568a91929a3a48edb4874d919a9ad3789fcd909d8181cef6d36673344218148dfa5b6c4b530;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4565f87e6ec73f2cbc2d0866619a5dbee511709c5fd696b26cf47a58a2c164856836c98f8a1f95d5dd721b9400719302f5d21f5779d416350be56b3585d5f21107cee86a9d88ca70012af617a855099b9732877e18be4b2932863e51b03816a2cb4241908fb287cb617dff0dba7662387;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc2910a6bd7e13d562aa4187863b54eee10a80a00c5eb07e7b7a69b35e2e35e20673d5f9a945147cf950820adefd85d20c7a57471215b6da425a6687438ea955bd9284a7662cea2d46d18b50fdd702d56ee937cc8461030443d6a6742a203005e932779cb93f993180d47a9e2310e977a5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c1552d6e099d0dd8ee9095f5d62458495b5a6f657ca5284ef74960b41bf8e25145c96758f5105140e4aca47306aafbe5caeb32ab7ea485d8d27c19920f545fcc2915c7f00a28fa7b34d56d0ff86f45352afc3203780a777d2f25c8fd5d9828865d061dad663142c961fadb8eebbfdcc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3a085b5d934f1ba413226e1aaa76af9e1c6675aa8ac273b214e52af86a9137d91fb0671deb69edfa517a8ecb95736de88a5bad1935973fb81bd793868c8b9f503fff0fb90fafbfa6e1191253dbebb3b99712a17a0f57bdaacaffbb9dc4cedc0d92561e991273dbe2867e8e5e29b80649;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47f39c4c6341789365c6eab2034f58b0f491a63886cafa7223a29be146ce3a24b46493f84c59147b90a61f7fa66dd8b7c73431f022ce04928d46e7e52830774256c390c20e469495a8c8b34c669406eb6f905ad07b316bcc7d41b5ab29a4787b38b814d453b1a24cd9c6973b7fc652567;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h46b4d30dc3e7e24a49fcc33857fdada417f34520b7da8afa5df1f1d3fffe17d948ddf3794afa5ad197fd9e7af2a3132b4d9cacfe9858639fbb4aa6c1b0da1da486c2d231dcf24e5932c045bb40bd6785dd73cdef6c86e481bddf4a42ca7a46cc58ad4ce20d79650b2b59b2d4fd99274a9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h496731688ea1b93652f3c8beaac9bb2bf02d1347f47b30e3d28e47237b9b2fdecd078c31fb8d6204153bd0a440f908059d8d47174693c92df801181ab043fe50895a85fa9e7e42d5f420dc307208165c7540e39d77a8f2a69ca46bc5c4ab8ad7a1ec6b7f4aee4efb9e14465f832b86d3e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf6645837de0c400f6261e44c97bf6db3fff86c1ed25aac92e5346a8835dc64c61e7daea96f060aeebb2a83a03c4184d488d228bb4458b5f3464b2c5a14d0dc6fa6bd09ef277fdba6c8639f1aa523fed4d4f467eb6111221f50bc627f21c23ad2d009a71a1fa14130cae1166ccef7b70f9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h60f779f894b93b2a7596e0d95717afeed41f8327cb9344c4b77dcc1b31e69c94b5b64b091099dde93c12cf356803abd21e98e2c9643f8eaaeaeaaa34828a972a8a7f694be319ce98bbbc678ce4fc1caf58fe986d2e1de996e60f619ce5d60a7bb45f4f668ae3c942bbdecca6d1893bc3b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e6001e8d27399c1be171031fdb33bcb7bcc655f1dafd4dd153efd37dd996359c99505f9ddd534b477f8e1a598ba1d149eff6d7f9809480eaccc74d49a2886d3f32d603ecbb2dc222610a4b96a1db1b213ae6a852f957081f26bcfc9ca954cdc4ae6bbd7a616f783f110c861fc578fce1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h160a8ac4f40a1dc209a5101cb0518b155b83732c63edee411942b1855eeaae94963845c6000bc0200fcd861e8895978a7c841c3ab0918b9472918ef74d657163faaf039a8c5215b1b00ed2327c22928538587a6a5ad09596701e6d97e54119d094f3c5ac42f94d95d08bce6bc3514ac44;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h438dda8100515c4f0257edb70bd85b42df86f05cf8d795a6113a7abf962ab0089598cf1c2d6afb61ecf8540b75ff8903778bf38cd4ce65bcecaea6130d1df385c64f73198acaa15f5082cea592f6b4056bb63d07c989c2d6e87556d44459e35a1f6fe6dd456c51f40df3f5826fdee752;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8329d963e800399aeeb5d762ac2426144bf3b64feb344e8da4032b9965808478c0035d74ca3070be333b80863a7a9e82ce801e7fd66e92c7cbe7de40ac6648c9cbdb05fe7fd46ef3ef9829004de951b8a1ff6e77c630e5e42a94c1e1e6b295611ce10cb26e1418e2cd6f2817b042918d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ee6665445c62eef74903868d7c13100afa724dd61669357b79e6befefa58737e4e9ea11679d897ccc00747a151bd292ee7b07ba4a0d539ba6da783479490bafcb68a1cb0cc2339795b44a17595f81f9634b132e339f5221064b9586e36cca150ce678ff5eda3b25801369ea3b1a921c7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h369230a4ebffdf0179ca25dfc6cffd78c19d1daa7bf0147a5d56507857941b5a87c8dd94e633573c5afbfe4c61430be59fafe248e3528ac9055cc3b6a25d9b4c43ad9b4c6bd7002733cde4b05eb03db1367b684ee0c4c1361d377aaa23d54c468a39b1e1cdddf394f56e98b9b1ee982b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a02e501a220d4ea6b8ca2024995df92163ebd5a9736fef6764a1f0c5201208f41871689db78fcd00b7f6da4cef628421093e3dd5ac0bf37197de35279d5c0fea758a3e11432f269bbe2e31efda94cd5eae51395e1bba50074b6a24241366f259a6c935bdc583dc6879eb1479a4f88142;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4ffbcbc5b633556fd0cdf497f5d419e657cebc35e13c5a1a32119adec6bf34a9d2f230d7ec95f5c3ecce6541509e82dd428623fc6e25d65ca21907d5a1db4e80cfa7feeddfbb659b8e922eee5431d7d86dfde55c5d6e6856ca046de5d096f56056129f06ab9d5fd1ff4cc3f92917356c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8526e63e0732a836c96f1c5d8361a6ea4dd6021e8f55fc0a585e482097105fdcfa2e7700eb41089477672b66a202359d7ad556b8adf86b2ad98ef9d12ea64309ee1aef54df419a454481abf578b2f720b39de32694b6771cf17d9cb7d68cd62f86c486f6c98ab95b816ec1ddf6656d724;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22a9bbe6c503dc99a56f98111a20e9ea9082d8bc5d976273870765635ba6f5569bcf634491190bb26fa4404ec1535d5912d25d452264f3b507fc8f0c8018694898791dc03d7adf0c82f00f3de17f1ad4d9bc29164c6e11b06091c8de84bd4ab775f4c612593c51b4f8e2222e711c55fb5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9fc47220eaac2d7cb8ca082aeabbdcd127b1aa045ec24fad5b8ba6c069d0539ff6ad2a9e8d85f9cef91d116d6f0bd0416d0de5446ff16280921b257fd8b314a6af9a11a97038322f914475d36239afed62bf4537864e7210a2d1f7bd4024c280572f3b2ef10122213e5849883ec37d270;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47edfee97740a981de419b273d4db12a017ba4a715a8ef724accd5bf6a7d11d1f53fa18277a8c9076bad1c24d8be2cdadbb19d3134c3cc32915599be96434f1445a63b32ff8fbeb0cd84252455b777262f8e091d463653eb2a63e0a4bba6801d06aa125e2b3691d5f04f4cf086fef25cb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e3ef553cdf7a239f63f9e7854d3bda48508fcae62a3b6312bdba9f2b7748b21d0b6abb140aadcae06097e65ef18b5ed5591f45dd51cfc835e4256fa047f59b0ee5dbb251da850cf20bd0ac991e22a69f1ec309eafc069a12da59ed63f11e8df587513329634d57451761820f9790250c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha7c2cb501a20b9658a3dc239e0d48ef9a7e9a9ff39c80502e589f56587ddb8cf23fb4200cb70ee2c2bf9436eaaaae85ed3efb7541181684e8ab31339a783abec51390693c3f07e1134e284fd61bd1b0819a1b5087ff57f45ad14b9d5519be95bd3d40ae2efdcf2fa3ec968387494f1fcf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44b4e280273496740f8d3700e1d6134b649e0e864ea9298f19ffbab3df513dbc081d36226269c13d5e683a9ce260c38f3f48f8d13de17b0fec271a37a6301ea812dd50e29ebc792968875ac5c9e42ed65b88e1953df9623792022b7bdc839ffeea2ffe9d0def158e8ddc809a9c2ff20e0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23b34e62c86d22bca319b857c7db4b3cfb4e620f9424b705398f2d56ede39cecf433dd6b2cef7ee4dca1be30d4a01cf7fbcedc776a3543f82a57e967da077bf51dc31f20632d51e08cf858fad53158b2e2a5ea40978ee3c03f949ea27443fde12fa272a6cf10bca32cf2ff4a24998613c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80ed524c37436220d6dc77a3780d5e343ec38e2a58be812ec6d0d733c17c01644e5a1aaefd09fe0bc4690e8135708594092fdc4f20974b259ec81927a758682c74c60c1ab5581741420c2b7b8f78f609a6177b88e60761636b2fcc92920d998a8eb66b657376300ef8c091e56b1e161eb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b0e79d994f9138d8dd1fd3ece6c08d544b6b2f396c3e4d20301675a888dd318280628bfee612e0add8f79fd126caa4e1cc166c171f94e633cab1ec7c3d4fbbb71265fd7ddcc21275b234b2cea0568602d6e1963e80b7406ad3d2d02b1199d8c757d7dc70e53472671333d7010c8641d5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ef901c8edfd43fb15182eb835c8bad63b3f31bee2b7104ff33229c534629db13c19bfb187b804322e6263c3325fec21cff0a9e5f87b9ad4826aaca7091100765b044a660c1fb91a77c438eb30b47a7eb0bb1f75e983dcf1dc496544a30e3057cfbf4759c29277ad1739b39893b8396c3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4b73b8601df9167cb59ce2932a3efc30ca8f92a27bc5d054ef11f9b37eb662a379210b599bdb87aad33aec153b17e1cbe4a3af2441881b0eea07e32090d33dd9b8675dd4fb718686bebe424d17cf6cbc6f8264d3875a88e40deed7a95485945fe855d02d5efbaf1a30b93058b75c6673;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8b37558a52ef50c47b59c1054a26d16a1ec7e706c6eb255c864908df96d6478782b643564a1c66f8114074de224e61499681aee5138820c96790c93b82941068ae38bba6be51cdce62ad8bcea9e36bb9183f8bc3e65eda11e322cf1bea556fe74e8dd2d1151897e83b9ce2704ea3949e1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd1cfd96901ca4f92ff3fe3e71795f58b5e1683cc9165f104755d3172a60d568f3c531003012e8cbff8d54b2014445bd0de6b3d4b2293dff0d2841391b47e0870e004ffbbf0b33d6fac0895e6409f29a065489d55e557808a5188150934c090ed577f235bf0a2f51270502de57cb018653;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h403428a25471a0db54fe46e46c3306ad2ef45db995f3c16bf23c7d63305ec54f11215a6a2a8b5a78042750faed12c8526b26d0abbdab4a68064a0204ee259de4b760f25b9e0354a0bf24b9940b4df7e5eb65bf4dc71aa46b3e2842224c0e5843c02e955c02b12c426f21a25e8e605e12b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5c067a62401d9e757f7225b49f8630073f548a8f43483b80eeec98e9f63fdef5af489427f82f2e1a689278ed24423cfc512a20f176bb09cf787f432e7a740102cdcfb85a58ee328d1306d16a496b60cbaa5e23991317b154789581ffc2e8b27a2d96c5a1b09abcff450e113f865bbcb3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5effa38dba3d9dd7444f617e4725cb4feae673ff73f87b6b7a9ea8729937e3fce6745b72d4435a259f35291d388bb29388a59d226da4f632d330354e237ecda88a1c6029c5b3598cb1574e015251f80d3888e2dcabf3fc385ce29c7034a8d37d78fe5607808801674ee16c2b3b9d6d67;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d2db4ee082572aaf3397d455596d3c4e2ca206ddc728461f37b6bde2798eb8ea949603cdacfcc78c4305dd67a0809616ca443686babe2954d88947f6c110a3d037e48044368434facb6a6ef2d8ddffb97daedf39b78d5bc74737884917c6a33a40e6569aee3840e87c5a768800288272;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d475a25880fb7d1970219d7f60882e37afaeaca6deec959c948f7f82ec09de41e372b811c9053345438543b32526675047fd19006295cb8d27f25a5b11ab75ceb2ff8d4418c1f2a4d16c86d08fba1a34ab960d86566b10abd22b7a4df0d9ee955063bb5fd2c520105fce87bbb86fcb76;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50f32b54e5aadc1e4939e964ed9a7ccbaaa74302318920b9a0d02c669a0dc8670df4b43f2fa6fe125a39265e98e6428d4e2b57bb5c0206a3693bcdc1a1ac0e3703127af4fadd4a507f6714dddd8c312de3bd77928aa986692e1f9bd2adf1ce173ccb4978061b34ca15eb80379c534ee2b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ebacdd565ed91fe61a50257ed474715052559bfb808a411e156110213fbf18054fa796b789abc30fb10699876941335c089d81132e16280a1ce1610e7de3986a4e262bb5f86f9e13b235eaf4a283b7fb0f856d31e94d4cbcb230738877dca7e575a18bafbb30abf238f519c6e42b85b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haaabb37332a4d73fd9d269367d8053e8ac526f346dcb651e3b3d58e4d9d31adbde716f40839dfaafeb90ffb58ae67a35e42abcbf809fa829836583380fe2a8823e32d9cc5ce19d9c9c92ca1c11f66a5f2ea7c8a81dc068dcf1b85e2e1f473547f353ba666785d5aecda3b863c7b2085af;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42b583c5ac628f4073601f50d5f194b0b25d16adfd10b054017544cfffd6882aa7378a8f50d50db03ea47c5fd1116fd4f9f05bf76c8adf01250f6da40b2e651cf15d0b695a813d48649cf76fa5ad6a1509b5162defcc31252295822de1217a197df76fa878cd19bd9ab81abe4ab750d19;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9542e287e8b3b3c59cc29a57f2204b0c42a6cd823c7efa21d640fb6d6061bcf1cc8306791863043562a0cc04b27eef6ef4fc5ee54b0fc69abb74b0fc2503c6a4aa50d5a12373c1fca3b57ab62b3925a4abe52b022238da0aae2d6666fb777a4d7cd6d5a66364a87158c8c455c63db9c37;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30928eca2153f668673b402c872cdb61f91fed4d326c0ac5f4b6f0921ed3f04b78b3d2e6d5fc46c530c647110b270dc77fd8c25b95775ab6f5a245166f96c67dd5dc0fc427f20f95760dbd2a7e096f303ca63b703a54f2a4f6da17d87a12867f7891f74ddbd862651cef4eb81bc30d890;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h424d6dd6cc817f8c41b4a5d10388584f729daf38a1f8f7e19eca89853400a03d375454ac6655e95e9793a682882004d80e318831ef365acb963456981338e3f2e59d5f1c54089d947da98c943299982023114b00da78e88c6c8b18119b382a6633f1ec9c3eb54f89b9168a2e18d0410c8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h21e4b55ffd1f0067c5b00e7ed284c76ef11dfd7a18abc2d3b21f49be957539a7f547980508b0eeef762edc60cbb5312bfd470cd6a96c33ba5dc1cd20ec2cbfba7b9db9561250fd6ddf0a87d6f97d549d963cc34ee8f2e8f69e18119b3d1fd129ccc65e473094a593689c148105b832106;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66bf0952d55bed22b995634b34d99ad9d255b078554a17d484a5d88591930d14005f09afcd01c85630a66d24d3d7c58214d2241972505cd72df13534dafa7aaac00d12339fdadc4fe68b5013a781ff3d15ab95fef689effcf2d1a68ea0cb9551a07ae606baf6c5326a50b4082acb4a96b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a0e9d17d28ecb3db04d2229fcc900f661f78faeb4b8a1d88c1d84d448327610bcc47c79a2f5e1a29380ef9550d30457c7bddec1786d2eca0c154d96bb209e900f68c0c2533d808108d46e82c94d32648608254fc0f3ce3a76bff9e03f41e46c4d706540bb6677da1343938cbedd34b96;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61c697416950ef8766a9841836877a5e4ff671b673a1e12630b3c2af93ccccb74e41e860fd4c59f769921abbb17a5aab8f739f93f874429fab5ac169510a53851e687c7ba96bf3a41dbd02f7c8575a5d6698602ce254d320132c347129678edb5e58a8b457f92bb5b12d7645f58d86644;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d2ce0dc95c4d8177c37832572d7814f9ff54b0b5d49f85ebc5b494e8cbf7834564538a5c30181f03998a1d560346bedc424b1589400d4517e32f0e16e4dc41482d99d5851667971e2f3baafe8a72c8e66a06f56e2f64845a9be28e69cad1d79eb03fbb40dd78f14c8d2e4171df6573be;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h592e6631ae123c3ae01b698cc047f14d19b2211e81d56457f2d0031c8d89a62739c04a088bef88b026f13ce0d7d2d6d668fae605d9802d45d525b3ee41bd85f28229801b82892a9d0d448c4e6298616c90ab7ac707d32f157cb528598d6e4999d26bc5dc505c00a6a8f8a6225e8b15b5c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d0c3a94ce02d24bfa7255c3a56f6dd2a986752fb092a089344ca44c157402212788553d8d80b0b8476b6499457f1563ef39ad931f0f5b7463cdcad27a5f2635bd6810524bcbe609571904dad53bb8ef24949092caa9e680fa102b6b990412d9f963ec7ce4fd54f6af0e86894935c3d1f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'habb65f8fdf441957d1f382b01731fbfa1f1f4a7ee06a3ae2597172a407762ee87bf059eca666f0c34c19fc771c7239da0d80eaba84844f4bdd02abb13f0cab67a73674d0003e7ff409ffe3f7cd87bcea66113ba5ce8c427c12eb73d72763ba3c2121d07b99c2cec01e8e7460089ba29f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab7432a5e6dc9c9e5d59a195c4aeaa8d2fca65b6852d8f933309fa701255a8fab6a9268c545d6648ffb40fa3f4b0beb3aa3ee8324dc720ad88ab916d13253ee9fe9f810a767cb6a9ef69e7e5f18897e6341c60f1e02039cb3905a1ab5edc3c18b3ac240ea123d11c73d36ecd6f58b19b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ef61a64a0a0a034f6c05ccc66469db0ab2452eb45259c189e09e91160612d749029307738a282211b92fb6eab02df3c5d53e9afc017b00ab545d6da4011701378343bd5ba9cf072719253932742007896099b858856993ac375268e20df7d098bf2249103e9646fc62827e6f78b8a26d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f3915ee1108e4a6656157fc2198f57b60d8d2b1938af258e3021a6cda2176783c00d93e82bc3e61cb7e051b288766e22249ab084528f020260789e29b90ea73f5e7afa9395e4585a45e82d459ee0c50c3dbdca1c68aea8d6506ce0796bf66a32c81a8b10326040a21d66b1f4f5321bd3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e1d71628738a8ff2c81c4ad91c7c10e0193d69529c7f0bfcf36d3d4799f6927c12fe85538a4b255be90e1748b16cdd450b49ba5dec3bd4accf6916eeaca48f6cc73e47dbab32990c91d45a40d3aee896831c2fa63ad07c1e1bfd0e22ab53cd90bb8ffcdb1159e10197314ceff05affcb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55a8c6484280d9e728df610daffae76c318912df5f59e72bf801c408c415f646d308d787e6db6bc8511682472aa44b5f7e9fdf4fea4a6f72475bd1334ef8da15ed102a7c97267797d16e0defa00257b2d556e92fbd046193b2bb34ae481ac7f4e00919c94468da63a4fc54816aee2a519;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hebc8f0aef7588147e2d6532f566148a0289de339b201bf039694de2d8e026bef4dfa71f730bca73f0fcab7894d3ddea7dd50a5d2669c0e2afd1b01a8c82a0cf2627d288b696a6599fb46517791f034522e8450176fa5ba5f21ae8e1c3d5423a72436a01bd73b6d132fa9ca67f0b6283b2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b0249d33dcd998975196989ae3e45ea7d965a5fa4c030d177673d5c84d7db911d74d70dbce26e1719bcaa9a2424b645fe267cbbba7be34b5adb9a7c9f21af8c99f9ea86c59ac37234f6b4e960ff63d86509b3ccb6366049771d5dcdadc5a28b1fa141acaa860d3fd9d7a164a484ded51;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h683d4c03d4a947386f8d0553d20afacf8865436355d5e01d96137a422927a6ddea87b13ee50e009e88ea85b1c05a0b1775f1b0cbc0adea70b150fc291df61d36612459a5b99548b0d4059e04ecf692f6a3317fff4a18d50143846db2e4083f02a575cecddb9add11920b0b6aa01d30a04;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h141c79078b7b336dee1ce22d424a71445b31e394c62128ce1f4e42f9afbab81195b0b2bac96279fc4e7a579da47a6c98d6c270666a49aae0099d9761b6ca0f1b59f1dced4fca6f3fb79699c4cd7be160dcbaaf58ccf118e7e5b207d794b5629b1f19c8343ad22a0871f4ada4d0bc3ab9e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd19c8f3ce4077ce646671245633f658673475739f2272872687c5864246556ab1c5fbfabeeeffe978304f45526aa1e3c61a2c4959749dbf1901d3321bc600b78448daca53384391f0d12ce0d78745eb9ca9631a5d3c8abe6470869c98784321265ba8ea5964fcecbbe2ab26ffa8a0bb0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d61ac6d7a575158551b0181d54680ecfb2ce7175ca2dbf6019708dac9afb1816fd43c632863040485877082a9d5d0270300ef89b2d01798af76f1c20cda0ed1146499a5afbaa1bdb713707502fbb13aec3196c3604c474827603fdff7da2c7940a35aa61a2fce5bf9aab0a85a33a8bc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h330170b7ded93ba1ca9f6ad238c1c0c377913e781d63136d9f48d80d9e7ef7b9ebb98454aebd6227d74feff695e02988ebd3b412aa5afa2056b9746784b5838536fefcf7a6656553176b8355e3b990bc741c00a36c474703a6a583bc411c3635357e7dd9d4a5fe2779790083ea9dac7d1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h234667a3db41306c003b19c9273be0b55767b24daf1e3e4ff349e59f8226e8365e1930e3229eaf685027a71a72224721dd536a29e73b6c21699359071d7b33ba4a08a9499d5da37b2508454aee61d920b73b66153a9dcdba1f48ad0350f27aed3a6802c8f60721957e016d9f50b6e5bab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23aec954fdbce737c8ab91dd56ff546521be91517bb1c2741dff403443a3f642c3cc285ae930df742b7e66089d73d863291d64a10f836f1fd61e243f68b0e0236e00b9d74564b1d0e11e1b07b6be54b89f7a280d0a7432c1a22ec096a5497ef8c6dd1d31650440a6ddff156bd96386407;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h41f5119a61b5b61a831b605ce20c1c491950173ff40b6b6705bf81aab85b96804c838f08d06474b086f1cbd17c44262be569fdb771b4fd705c6603cd6f8028de6d21ea4c68e5f9d9b5c70a41e4705982321374d9e9ca23cd5d7a104fbb93bc243a7b8a95d7ce9f643a198a1feffaa00e2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f976f492b1823d2a3644ef58238afd8fb833f011fad5df3defa50b3a0a105eb36adee414d499c3183b9aa35e1ea8efebc7e183d8d66b93d0859c39cc4921d0e5bc4fdf56157bccbc7b9141285c56cee3328a54c4449bf57b5e8815de47a91519a943d4bf3f0e6c6dfd7e6d9f2c40de61;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd1f44ec79a8988fe22c080f3d13bf5ad44e1cc543474dabf3c57aab9f35d0be0292f01fae3a05cc3237e10d39866cd9680cc5c7cea1319a1dc66aaf3b1749c78f8df47a7573e615894f74497ab6ad75452e7ec21df06a03d6e26ad9a89cf8557a930d6a04ff794104b7dca3cd7a780fb2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17cbb672b1b7d47cd7a4dfc3c0e3f42e413ccf57bf7c00e4a91f2ee7fe186ef1e63cc98b63f1eaa156d53d07a6f3cdad6d582e2592098d2a525a07fc312ead1b74886a5109a539a1e39c90d2f7723485cce155acfea50fddeb8026ecb3dd54a8994d0364b9af282f1dfd86dac8f0ad1cc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1f958bf28ad98e4556c1c63f133f2e24c0b587d85dcf28da107448b362574f2360807485e7dc299a93e060fd02b293759a209bd118cb8ba17017bec636f7dc4adb2b68ecf1fefb40c7836340f7f9e27eb6df10e0cf95466a9d14e309f99eb493131f8bc87e6a2c0c90fed7849e46cb05;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h20904531e680f6191633f68397486ed83b26728898759bd6f3028e95fe881bfe4a979733af3ad1aaac191b641d345d8603ed3c2010b97a0cf7c3dfa52419f04bb050a662143565adcec097ab5710fd6bab49745b37972b67ec23bfd59b855437f65a5c1b2de35eda77a695f39043e8465;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha8245a60c8ddf122a5e5b7ae895396baa44fed30a652e69ec1e12c157b0c59f2a8e283eeac74fe6d91a58267250a1f28c71bcac177aee82e68f5f6256c8ac13d5f8f7366e4ffbd8bd382b1e34f68b155d2eb5f2f2d1b86ca20729a6f55805d91db125850f9c2e1b41604fa87b956cf7a5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9fcac9ceeac0a825495ae1874b110eb6f6bee486aa0b4385757e573e73c9728d195e735c029b390b660df824e717616710c29e45c66d8c3f2dc538de291660ffc8e1e44819824cdb78e3604d1e2d3139b1ab320f64d7d35ee1757cd7c3ec284d1660d8da9255f1ad3ca68941419a3f1b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h59764134f95c848fa64f94c3f7c2bb0e0cfdcad3d8cc53532a6c4db2d6e76ff76a53549b12ce37b7c5e48493190b7c403090228b8bf279887ab143266ba943182a8672209acc42230dfcf83c43222ba4d5902ab87e26f21cee08fec87d2c29a81ae7e99658633372f8cc92c4c9f7bff86;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe3dae9ae01d11b9c5e3bc26cc638334ca1b4557602c234021b233e4cb21d7c82b98d6bca202b239f05185ec54acd54ed9dfdc32b3e09832d59eba018fe99178ab96a7fc48a2c9fa7960ed3d01b288e97a63c9c7cd7eb8fed46c52d292a4e96864e83df0d71219dc6ec7b994c165062be;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed6a9f32765ba60cd42b2281a871d0617607c64e212cbd8816d6f97efeba940365b0a018c6481d8737235831311b4af6b4706b7d008b5987c813f5ceed2873899d9f52237efc61e7c0c141a7fcb7a0f369a3e1ef2c005e871d50b530623c549eae20925732317a4f97f62ee6780610175;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h587553b762a965c6a9e17aebbb765335bc692282fae322b7d111aa275d4b411d1c81899b8f6bdcd4851fd811645d39a2bbf1e9b9cbf6ac5b584e5db3b66870bfeab97f98042c4a7556fc4442da873c3ab96cccc0a18b0b3892eea86af7599cf88228255a6c2dd29f678c1c29979a17d5b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h831fdc79d5f0124ed2a2937172db977636e43ec2da2f4fa3892d429abc5b86fb6dd8007e49a9f70571383ea5c2161cf95bb46c6f5d884f986425fc5a02fb3401498d04a217a7f86a7ce0265f1d8587d513413f403ab37467075ff018c00b4cffd5d10ab2d4978e35c3ecedaf45424aa5f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a3e09a049508c1b108bb796865a1a9a1881a221477995085b58617a2850bb871acccfe14f9368e507525e4961e49bf59e64bcfed907258459a17c06fe9fd4ce2f708ca9d42418b07047ece08900647bc413d05de0fe431dcdcd05e3db334c7a5b164347eeceaac4545faf1b7600b3f3e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf03220d5429eb5e7ca1c29df467355ecc0a6755fcbec516fb2d8a8e9d08277151acc374a590ae793fce1a207a2bf4aa09cd1de9a4835e7e27b2d4da89e3af30f3c850693e4b8154acda547b4b9305ed7aab3b177ecf6d97b54f5891f6db03726487a6dccd0540152a993f7a8a864da837;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6742a628c41addf77f107fd505199a2bb9770e9c2bf05a80fd6501a2bb9b88b9f8c47d9cd01160d9fa645603d0d079f8eb26b1c2e7e003c29b4636f260aa0bdc8b88138507dde16f148b9c8343db184f799b40c9a4f4c9cf0aac9973bb10993641ae2f54dc33ea2a001f6ecfb62784cc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6aefaf1e211ddb56685b4792d0bdf2d01ff3a1f4f4f7347830c4a40b4cccc51cc5ce790861b61d31c3bb10cba8fc30a6d847a4e897929e5b4fea8509cab7b6493f7805028e9ef20840e652def3e22c7a5b6cf6ae1e7cd3a3e340be788edd6c1c2b12611847550a522d5b4b9e2353c5c3e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5143d8ea89ca895592ae67cf6732d0e9d187d854668a534389a30eb3402ef0765af5703b0bfce49de6a7fb189dc3f135c78e7cf0e957ba91174cdb5cabfe2027e8ca25bc3a99d065a47f40f521bdf1c6ddfc307d1965624f6e89f2319a4cbab714804b4cbf38bde5b5ee7066301cc97da;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1bae7adf9ed68a8d3af5f680cd4a15561684767453a5ab04b53ecd8f5e5b9f9b8a76ad895609c1ce0035d3effb75b00c691b3579395c261249f15a2c7ba7b68241b38d445fba9d01d65bd01b8e597b062b80c5fce62b93e00ef13f5943c4150ff9879cb99640e3d47f98d5e742be02dbe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87dc2d226bdc09cbd9399f11b8be312eb11d6830bb219d5e0a5bbbbe4c981c7fcb277550b25521903ab4571f9f34a1623d9f78f8bfa274ebc36076455a15731be9430c3ecb677aa41ff0771d230f804e523cdb4b8f628da79806af307cc5c94880ecccef8430e73a1d2de4c6a1b508f4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c6f351be61fa8e86a3c23e7b5a1b17a5e286586c83880e5d76d9a6a94013bbcaf20a7e59d9362f20c668a2345794ce367ca148f9f8a26c3cdaad02a1bfdb9fe6312e8b86d7c315c65e90d6adad5a2365788e6a23e14b0b6c8ade28c42cccd74a7b9d1736e87a8fa172392b0931586cd9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc93e4af2c885ec42e44369cbbe46787ac90a17b1a6d036656a808a9e9c2b7b68eeeab36e9d3e00e9f2121d0c5993b7be63e0b441862aa15800e0c1867fad79a87c971ced339a2f19071c073b9b4fa12d2ba29b37ba0b98394d0c6a78d39c986ce44ebb8c747dc2123add8fd4165292472;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h53fe63e1714aeaf4ac6d5b92ac43d273217e5cbfdf1e7ff802515fa9fed81f1598d71314973034aacae3c0f2404789dda9fef8d34320547ccf5081e6392dd8debd8751dc90bcb1ce0adf950799283240173a1088bf69e17e6df719949163937c5f02afd9ad358097e7d6c4e883073aff4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6775ca47d3555a90501beaefdb211c73f46841504f413e8429d6beed44920240cad4e653ceba23f8d62781d99f16dd61c51d08472f0fc8a993015dfa2eb94bd1316dfdeffd4e0810c534dff2704350c4ce60072de78432fe063d86ec636b21dd75fee7b478517c24caace902e9047df7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91735e2b3d6b975cf11d4ffc5f5ad3473b58284aad06a2498c1b426b23541517a9783f2ce27a0b08c83209aefb85d15ab79e002adeabe59d69ac882dea6d17b90096c02d361546ef395a03ab68c0be3659129a3440e7b67e4f39b086fcc3d761ab04006b9570b0f5af2e4c2cf3ed0f9f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb1f1c7f0db288c14f0268b2b6ad1853027a9afaf369d68ed8ec99f8e19467c218969515f935b6355e82885458949bd5deb295a61ed257b1ea5118f1d3115cc4923116f312a5b0daa5447cfa152f841f65da3366b15bab1c11adf86d31692ae9b036e5c6ad031213f0f5ec71a0f2c75e20;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5fef57af2dcd587765921f5a5d6601cf1c3b46205eb268f52123abb76bdbc22304a2f217670cde78d37b2bfdb9539ef192968cc69f7050043f57acc02c20005b9f9b8029478fcdaa224119dad33d21902702986f0642d071b6001775c6716177a2c5dcdf67b8c0f3c00bad1b633918c73;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe3da92d71fc6c2795ea58afa944bec3d261de90a86d42372e7956e4f4073fe6384630dd7c1c35bcda2555cce59ceef033d5b166bf903558d5a54eef5845fba2163109c4eb8662342a930009183b769a84eced287c3a0f99a059583d53cc404895e1b8b3dea94c20f3fb729a1cbdc835;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d9bc62d396b14c9a10747953175f68a80fbdaf876bc63f4aa6c7ef35cca877f77e85e8ffe2d05590f227772689887a88b01d5822572bcbaf333252905616ca6a813c6c8f1576c74419fc581e2f3a8e8483e5bd0bb2e04136758ecfa2a1590225c90b87d391448308737094c625ffc25e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h984e88c3b6e134e9b1719ee7224e633d3d97502f3dff9795197afd71cfb66b536928c59a3bd069f4dde091779dfc65d040b21e35b9ee45e6974ef4d958f3a0e813256641395e35b8036223b2b6b1225bd11fd4a2e5a5674d4b424a470c7eadafb67145b2b710604f0e3617523c2e5e3c9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb043f9fc0e4b739c5db97518ddb32abb291d624e1c1d0f2286e2e9b2b1c23e5052f03cd61843a6806b523c8d622b517c433f8134c58bb02f3a5b740ecc4fe9503f242a7bfd520823a18acd087bf670e34f97bc7a144db8f3003b60ee6de38cdd621255c90b421e62096f0059eb062e74;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd955a5a5899f659c51ec3589e328bcf8a579e97bbf47d63e54b6c162bfc01a1812ef16c6c4389ed214f754e2af0a5ceb730e63242c0d19d1545f44004caac392de7472419c8e215b5e7983099177d89b6854feef3870737b71328913d732d23fa3395b8084bdca0a7d5d224969cac043;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1e1847b0dfa44595a6b09e8e91edda60cecb12ff6867b3d1c5514e18089bebdf52aae0483d9544dc8c68437be31cbdef13e2e704b0b8b74e04875da39559d8e5c2bf22edf4eb0a8ceb1682b6b293921c166c6e23819cc9fed7f9ea748a15385174465834de2b0519e0017cd997d0114b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h747f501bbe98e2779aae06cadb1281abbd2d9081a88f9ec39aea19d90676f838afbc56685b43e3831c430973467cac0e83640beac3c1242f0bcfa4280415987de95596f9d31311f202ebbdc3ea948f43fb3b05bd326bae2920e5d47e16764844f104dd75dfc37edfdde9fd9ce2db7ea19;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd3609840418e1848845bec4e18fb86048f128487d125946ea9081a3d01fce9140a762426f030b2c39fc02d64d5ed018cb727f052af8d40cc24b5d0ffe5955c1f672c7972b752f11bb258a31c0163b6d644440bc2acaec988cd88356665ae39971adc43951329dd0e17cf7d0c99cca9955;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf51ff80f91390b47bee5361949042667d4e3f6665392e9101e662fc646f9a41e047450fe708fdd099a94dcea8698d676040cd4760b16880cf770134a1b614ff6199f7da6f9c92585903379a68d1d7238b54fa87f5e8d02a7548c355c2db91a9c5c8366988aa7c7b17d0548fad902a5403;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ddd9c9282b46e195e0215b402fcb88e3d5bc4af318e25dc2bee5d6fa32cf6249db7295536d12ef66d899881e19ef55014fbf79f791bb02b7663d8d48318c1bf19abb9570c3295fdc62a09a5526ca58389d95d25a3a58e6ccb552bddb1690ecdde1edce1afba57348abadbacf22367f9e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6dba6ac278e650bf36113ededefa62a0e73547eaa74252cb7e2934450597a31426cba23cad5f7536679955a2b6341a68e2a9eb7fbea6dee4351dfbb9a2231ff93fa92981def69c7d0fc1a8a02bd468595ecae315f3000495bb6c9ab8d716e3bb1f2e88bed0c3dcf47f8489f14991401e1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30e5be951c61e4e54905dc91e0e360fadbcd1533274e17a058dcccf94e06f204f09a8037c0a22e1f2bd50cf2aed0ad0557a215d5cf048a1ed9fc4879bcb236457a1b25c2c87eff38d16c24a044feec5945f1ecdb7f581407be38475a1e9d8876d8ce0463a175c865228b483e4b086185a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5a7c0f9907e2af2765199f02ae2119d70183f436a98aacc186abf605f5d7e57b271d328af75a348c232f09091cfce52fc04c2a980b87444e2a51dc3427d469518b505732a1a1e81a9fd0a5609a45f782cb90acba2163e2710da77cec50105c8ed301cb0d2226d7c8fcad5b1544cd0fc3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc91d1e5c8994092ab4c50bef5ddf6ee10ded045cf0ece9e111121a92d888a400a1ce7bcd4677ca6cadf96a1a1aa5f06853f099b05aba3e996ba7392ad4ef57f92d17f4b7760d61d0a034c383cda5eb92d121c9841dc514688a8407228a99706b7fcb11134b9eae21b74f6e1924cc2c5a4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5726473b1463ec665a5ffeda46af6eaef2f46fbca908d7845339159b5c6b56b579e9bfd9ea1c8086c0dd982544ef94c2504b9b52f23b5671029f7e6d7290af03a756313fc6c354cf7a1342051c159213d7c9a3e11a56653c98458eb04d13288c3d475871d6f601a7da41cf570f0d3bc2f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h82067e8ae32b59110cc081e300a90320748f579772eb4fbc0227039b217b97add65c5ff77779c4ed8102c8b1137b17dd9e58efa384274859abb51293cefba959b5bc32160b93a90b821422ca8ff73b8786a715bf1309758bf9ff0dcf78f1c5b3c8c63d3603bc8f9fbf7a44251e391de27;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb92a133a2b48749d299d3f2065b8b98f968529ff3e6792f562b971bb4a2703dce561dfa5d000fcc9992836d0683665933ee1aa0200acf29b8a6f451dc24ce605af3f8139aa74a27616113d280c83f98602c372a06a9f4818620399039b4791593770f73d75bba5928d670de4b32cad56e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc33418aa06cd80df54d89fa00a849f0238fe0240cf4e2dcfdb211766634c5975d3034699a75d71b0cf52d66c4622b0bd992ef694464896d0e0623a7476cd9c61efb51b751a6be93b9002165c0ae365d1dde2b3e6c4a87190eba2595d62e227434e1af0a9cf3bc3c53bc8f09a08ca0cb2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h68a1ec7ed577571d0e2e2fb519acf157a0374f8851fee7aa546cf6b1911f3e1bc62cd8d96f7b6c9a25dcc48ab4a8a58fb91f22448a92d9e223ffe05934da0786dd9eceb0c5ca6ed74f33ae657c3f22c9a94ced2192f450ef2d6510338f14bc4f4e98681a400ff7cfb443c04c8ac2b176f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hca055c4afb1ef91c050a2e02a00a0f00f52cd1cc77ee784fae7bfd2fafd57e33a4d7cb68f0430802ed77d58f8c42e3fbac6739b5146da985d82bf5b8daf83e6c5d8909e1dd5b44040bb8dc6b5bce52c3ce337a682d4381cf89b0c9bf71577933a35f7a1873c7878d5ad0500a647652449;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58c58ed8e8975fcf3e9d14b548cced823f597aafb1c04e3876cbde4d205f5039a4901a3c8a48e3f2b1119d91b1b1647222b58e8b2955ab9e7f562adeb32bf64c933593e17180cd86cbb87691c0c4e048269ef68b1c01ebf6d87bef75abff299163df58797b988f0de4949c061286fb20d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5a4cb2661715ca0894a57dd5223016f1f8d4c18315a9e8e6d2e609db0f6bad603d599578934d9e29917ca13ddc855ef33449ca8551bcc8015c807f3859cfcc80edba9de4a3513a2ce114478667188676e4ab10df1247271fdb762bced43e111a48bbc19f2e3af327899a2f58753d83fb0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcdf1677f434951b9bc569db55216156c6f14f6a909abc6d373d4d7d7b0c7b988b6c951b5f48b89a0277faaee6324535f8285eaa039cd4a5c93db979b4a97b8aefe5156d44103701c5499c731eb5402328fbf5d69bdde23fc557f30630945fb2c5df0090a8cea17c82a271e0081f1fa844;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b3020260b77172c2de64f43726a942fa9375bea74382fa5c5ea8526d5d94794a9d86a51d0c8fe838d8824fb7b685dc46779dc12e6f964bf4caf26eec7256d530c355af3fb57b3be49f6853efb5192c5698faf0b4b24a3a7a88b5c2b315ebd744c4c8414f80109f1f81ab36914c62a786;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee38dca6f5e584aae1b7e86721dafe7cdd0f318946a7750acd696edef93f6b3a7c23ac95efce07cc800613ca943c3aa3ad5021edb36479a05d4df14c3911c1e2b260f4b47692404f1af83cc31707e11a503120207b06b14fae4603ea9a0967c2973f61119f7043e39df2e90a01db5c952;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb091da2c4c9d2c7ff6c1700591fc7b63c2991290885c107ae33aaecf6927a47a746e299be9657976f8e5d325457e744475c868ba823f82cc3fa7d2fc2522123ae2e6e8a25867cec120647884b723ec1e4d0b1f842dc80020f31c408757a4d39067f1732415aee24d285cce966eaea37ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e6d9f92d6536aedc8c5fe579e9124beb47c7257255f3f0285e5d2f4645c30b4abbcd193940e2c97f23f92f5cde4a7fd9464a188964c669441153045423aa66015d8da66185fb2ac2e8530a267243527fb4c6d1587455ac614c678c58d1a583d1c9747e97c7735baa6d172bbd6af13cb9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8892d8d2e240ddcf14aeb39decb6f580ee15c156810fd22e26ffdb72bfbb02613e3308f3990b7048cdfeaa48480019830cd64422f7e3a5f139a6723ec23a819a8c213c6b180aebe32f9d07ab8ede8f438a134182f8a714c4629eb5d912d11b4b0970c68c39d3f3b50c150e027a62a5394;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45ef5da4409078271cf21f7b88fb8dc5852bc3355aaed39ee46260ff7f4412757e0751028356215ec9c9879bed1151ec359d9f31d70948b496d3bf031e04c2fec018098d87669753070cd427814f9d4e85db5972d33a00f5c1ad8448d38c89a975acd56637e7f1f03502737b890b4c754;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h698663a33f196a23cd16c6ec8e40824b0bbc4ecf2294e3eeb9bd7898a02e0280f9d0182232d865ba2d2c2d4b12fa08436112fe8e17f82372acac334e7e0f8eb91773981243ae312fd4648a8a11a7bfcc5fba243d16efa10ef1e13a9f568ece5129bd7d488cd684e20fc2e91aae5ed7a46;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heba0d235f7a8ca318e5ba892706a68a61413af9f3b46a9191b4336b38c593539d299831a4c948c7265b4885a0611a9598eaa3c0e0be846e2c5080bd7807fa52144349e3c92995cec255ae50b4c532a8357ca437e8e85ca6e03413eb66e363a1a805366b76b3257b304c11ce267c581ab9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc95eef9abee2c5f6ee24bb488b54f01ba323b60543fcd5da9c5210f3c3f2503dbeb502d61dde6600ffaccf25b02967a2a6503c6a3f11dd206cc14daa049055a7cf210798c69983fca2e16cb967217edcc4c02109d68510cc2975c6679ec047e1e5bec839fdf376c0aba184df92ed26305;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h73182f48bd6a5506d82f4ad3194c6c1e99f8f03f21ac801a48a17516fbf327c412048ed469e375ae761e6277574428833ba401224d2dbd39d6aee6f518bfe325db8c657602ca48b7d8556a0269fb7d7d848f9f409b43c64d26357f44921d8deaec82336ace65b9387adbaf8685bc126fb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7a9d97a653c9d754cba7691836311bab61f5da4cb7d12afb940e32fd15c2d65328193cfec92b4adf7e1fec99903fbd1911fde4576534628580120da87f74a0c3c32e82ef1d994b0555ce8bc15c435b3510a8031945111a0c9ba25fbffa874181a0bfdae0d277f81a5e2fdbd2ac68b616b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66b3b4e177ff908fce67c4f0fdd26edfdcdbc4af07f9ba11e533a4929f2208b3f84284722cb45f147c31c6291b94fcc67384cb85247d37833c362161df8f65030fea1b2534c6d99ef20ca8c7cda258b5d368c4fe5a8f8407161a7340547cdb9bc8f48f64d2629c49c3cba26f6a55b6221;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4eaf05e86b4f02257346c880cc2a392c456450c25d194ad6ea9ca5ad2c09d46a432be2393da7e8bc4aee7860479f9e47bd2ff15722f50c135511e64daf4b78936ae448544f96d555aed45cb941e4516d596834f716cd816744bd6b076423725f71c5965ebca67038aa296ada8b997e51;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb8329ed512db11b4ea56882391008001d9d74fb16d2042346713a801dd9a22ee37a73b4708a8467fb80a391bfaceade0ee32edc116acc9c11ab03c0680caaf080e982538ae2e4e9d79a58cd1fc91f1e1d32f0ab9e905641850a66aff2792546c9331756b3ac57679045a58697b37d90ba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc0cd65229e62e63e2531fbc0d76a66ae63de184c23a55cbe2fb96d94a25dad9231c90331dcaccd685e013f6dca09e1a776ed89cff0927e1471684e0fea6fca881fb431225af47f48f3fa780b4340f7088399844197c0591a28df3bd8080c67e9b65d79c02179b38fa77511bc3fa7bf0f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1c255a74a83d5470d5e190bd668de93b2bc10b51ce0bdd26ddc3de26cdeedc96c50ff9983704cc483e5d7cc6e28daff1028d03af2cf256f696379bdefa301febe65507b6bec560d740bb7048b6e93fc3f6d7aab4f2806be5fb2de527ee7ad53289c245d11a5938cac80f43d17d7b5165;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h671b71e3d1e72dbfbfcff1f33965830bd3ba0fb769b02ef725c0bd020750ed240170ed2aa694ef597cbd91866ecb0c385239762ca46c9af2fe7270b90e3b1c448bc928e20e8b240dff6d3f459720494520e323ee6b7d7962d954d6b51e357ba214dd636b15e0394b05d49784c1ad79aab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he697553918a512623762b9000f0d4810af36cbd58a2270466dff556da2819f776a299d4b0857131ff451d37449951ea8841e93d59a8c4a3d0e3147c6a002a3d3c1a09f386272233ac77eecb11e219310ef00be3b975cf9f9c4c3a616c5e19f5bace09bcfa12c78ebef05781d9148fa3b2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h705df596326b57016150426510212c16f985eab0ced193b96fd990597adb430435942ae9fd111a7e3a24b00cda234e8b1593860958fd8d335408694604dacae0a3c18cf5cdec01643267160580a404998e20ffcb407d08ebad0e709ea2112a3012e918e96f6d4dbb51da2de5e58341b3d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb023ce11dd704a117dba196e4aa72d208300a102f2c4c064f89790f6233f9265d3bb25e4defc1488c274cc9f3b4fadafd6fb1efbc0adf128f6be04ab72b6928d1c822bc70bad55ef027d72749e0b62af2e37449d1d0da1392369ec214247034829ef86a3755348a843d216c3a23b3974;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87d8d080cbb59de38886327d9df7b26d8ae73a88b52e4ea521904dd75de05648ec7b4106705d9a642e9fbf111eb76add0d75acee656ac229d027bdfcd6873420b316439f2b47bc7df82877a7ad2944382a26cebfe4b2707e37727b9dc4a780dde363e7bea61199adc3d661380ccd0eccd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2364b4de7d0757bf115e7ae9c13161b5e8ea86265b6556e0bd4bf0ec388d04db2c903bbd0930fb6170d2cf7f245527ee9961779a4710609bdd964b1804a6b8d6663e0077c01014d7bfe7e1a60802cf5c73ca6a21a83b6ffddbf930acd9e7f51ecb13e79711a5111479da812e9d862c2a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ffe0e3ab7de54cfa8025facdaf98edf8679fe5d7d8ed5c2be2bb33cc59c311524a729be42d2e2ae680ed96d9f77a1bfe76aa28ebe45165d12de20703d66ca7313c88c8ec66fc6c9259e40ea01ce78f79bf1c6b2ff639cb251d0c32ba233c9f9d674dfa541abe6812ca503b3e10dedf8b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4aa41077765afb247a58e18406e86d83a82ac1b94f51f0729a873fc6de96c64a05bbd5befff627331f8fb1b64810ce87b1878f828ae3d90eef2ae85b7dc3878f30bf92189001db0e06d6c176a460a3012af614ebbdce96b4b51d131a9de40f9c5ff565bc7c1d1ae64f6a14a459895d7f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7693db17e721b5a00ab457a7d2f44305641486c773894d914bbc2b474fe6d854bc06b5cba3dc053e06ca18cde427afe7e671e7f269d3dcad5bb9033e450e82230a4b1a1cad9a9ff3af296d758b418cd3393a7c0577f510effdd5d5165f58c86dc452dacfcb8dcc390cfe8a1f1cb837802;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1d29ec8557ef64fe7fe54d4cafa7fea9ee098cfae61f30487cddf043e662b085c193419f1d90fa8624d71dd21666dd88724b3451ee0ec88265741823e467d5bc881b315be64bb01dff4035823fa10e5317750dc068e4e9243f74f973b83d20f7f86a512d85add648cb268dac826d2ef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had13f8329600f37cd98b591b210c9a67172f2ef6ceccdec8aa0f79e4e64c1f3d7827ea71df8fa8e2577229c0c81e399f41870a837a19f04a84771c3589dbe08fdb33549ba10cbc942e372206cb743380998d5a6af8d8736ec412cbf3a23888f3dbd9c537c742fa9999ee2d69b96effcaa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92b556982d489df25b0bfbd10ff167d6b84415a6d2d8182eb0c33454c56328dc08c30bbeacffc685f96e0762c3a07239c11a73891aae79328f69a14664b48beb42b09f941beddc4fe1b12aa8c14631ae9742583230de2761d7d477183a8745c394f03e86cb4ba17320034c370d3959fda;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2020fa4184a3116bec9152579624f644e5983c9ef83dcba68acee93b60648641263516ff6826308d29d8784215b1706e1f1374ff3321ac925e03032fcbd5e903773bb9d121ede2e6e3e585600993566bb047a0f07a4491600b9568a490ad7bf436f551396a5770d8bf6760d248916042d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8c0423d321630ee4198900ee6c1421cecfcc19dd99ddaa7864352a1c074bbd677b9eb8fc53eb98c32a208f0d41c15e70c18d0497beaad43ae3bedb3767f9e1c331493b69b04a8ac57d9659ae037484aa8748fd65a1ceca36ffe8c2237791bb2dbb08b52eb3ac68e313c4011bb7af11c2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e8e227e25cbedaadcfc20cabb9b557fb72e2f5175271487b636f47af7ed5bb4f42d1735e396306a79628a2e879195b31ef313e8ba52f739514f3d6b8a8adc46419ba092ccc3e869217f68de63101d2c954dc24454c7bf1c2fc91fdf284b9e19da5e07cc9a3a868e69d14028dbb617c79;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff911ba9f9f97aa87019e05ad82b4289d198cd858a1093d82f5bec55987305a5fa855283a38645d31643e1669803b50a5298b756c6829e4720ac17f890e00824133c72fd2642db42085f9077c003637a134c3498823277b5e56863d04ef67eb6ce760505af395c2fed81a7a7c6355860f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h39b2a5f8eb13ec2ae9f4b48c9f824ad9ae79d7e7d289b29a7362611490c4ed63aa8fe74e105bd814031dd41d337a985e3115d7bfbfb2f7a558dee67a1d830152ff61cb2cdfb703f6efe8e81877d8049f861c10a5b30bf04eb85bc5f9dd4461e5ec20d4a4ec9b93b0965093985ffb47e01;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbf6c9c7c85ad7496bac022e5ca3effd7c51d5fc37bc6d070292d5b6303d3d5c4d99d8695d5174609a00cccbb5289dd954d7ca674642c2018a4123f34d8eb86ce974867e58d1ccea95702da35d0208183f807b638b9b87e3e02a7bcd5839c725ca530bfb9d0b7f05f01f79c2b927e035a9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64658f092c612f62fe802e73450c9303fef67469c3e1b8e03560c88fadc87509f6960010e32860eebf3b6ca3fcb67a93df33f609f085086cfc54caede52b6f37d0fc1c60e993f807cb78499c29a04a96d0296cdaeff49b622dce968d2a28c97e6241a25e1872349367aa818d4fc20c042;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6fc5dfb164e3b029af8810bdf8f44e07335e3f8ef1a94f30a28ee2807b39211c551d55e694953daffda0af84b1743f583c217cc0eb5fb805c6b2d4aceaef5ea15638f619bb1d13bc003bc74b1400e65e62aa59e91963a4a50544992cf9b722cb6811a82321008576717bbb9473dd9c3e6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd08bde9ae2992f00a7edb11b9fadd132fc2a08e8de6760d777fdc30aeea4121b063542563e3df5371f7e7d92011f41c35b02a0d52e87ec1173972fdad0f3d227429346bc1d1181dbfbc6c5ad98b7063b540ae47591cad3982fcac04caf22ee5a96b595941601ca31642a43e4cdaf2d4fb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h22b22fb13d5e7b310d39dc1b043b87e74f3dc2b61d3acfbc8225ece0daf3da371f6de9663502425795b1f1807ca5e9ed39363ec1df3e38eda43af58c3d599d171d65f876f61916d54d8623f7a231f80851d836aeb652cc361a678eb81ce47ae0f5d35766084578bf9b08015ca111d965;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4726468bdfe09701425ac5ef1d1dd0e754a0e6bd2cb8c5aaf6c7547abae27ee582bb6fe572d6a07c57615480493e5452069b18bf9a8158bb329ae8d5b54e3051433cfe8ad0e45fa5f6074328c489ce80fecbc42d4ad0cb938ec880332097e2c81e2fa2ebbb7b96b204948405e6177f09;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc6783d47edf98365d64e8df882aeb85ce257ae12e1ffc5edffe5be0a5810cdad4dde5ada81028af56ef259cecfaf8488641d65d7f8910378344dedf4890386e2313c4a8ee63582ead12066d4eff2ad7aaae96e3ec2cd21ad19e9ed60b49ffacd04adccc7a8503902979c5b438687aa87b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e71d60fb121f7189df67527951fcd25f05ad8bcc9e9fb95810e1a008ff44a287192b08eb81af9e0a1d8cb21019c2b90dff1d220cf925934b020b94b8528628aa7f0e3d1561d078eb10bf4755c85c9db0c164ebd49640bb6a18e43dfa35b3a3af4feb8756618fcdeed3ddb5da2c66dd0d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d912281a4930dc681e3b426de1b69564d281620188aa65d2730b075af4ada5774fa8dfdc43d8fe065f81bfb812513fba7e68a4f7446c1a5ce3377fd65c7f953b620d9caa411b4095994fa2b0071c763ece7ff56d1743f2d21ef42a5dc94a884b590aaf9628d8f80633039d8177ab524a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h962a60203246282942b4c4d2ee4f9ea9d7ca59eb5b5437d982b5df4c58587c1858d957d9e982a316765de34d0f50a2fc85a5f602952ae80be285de59b51ff5f8219611851d982a91c1ccb2571bed8e150bf7eb9d734149e33ae26ec8d6a6ca62cdb26ee1f23d244b7a4fb1da5ddf22ab7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4103622a7862370b68404067fdaed8d6348ca6518fb6bdb44d6b8c2d0af278276641c4d7ba32f9ecf5c63dc3ea0c51a68c6a3e4025c18b232c8a50aff246301eb0b70681e40692793cce9f631efa106b8f5fb211f4322ce5c38fe547abaf8e65caf3bc4ba06dd8bf7551b196a823ab722;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14b59c8f105439312d712ea29f21a2d2b7ae33028fee63c210c6b69e96eef7b40c7e892c57904c64ab54a43047d5946885b4a9aeb3c149e78aec1b8910e65d1b11db47be7ecc7fdad483320dab2ef66ba4076f3a818127a1e649ec0683b5ddae2b54a434d9ba603c45f26bfc453d0a629;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5847cd4b0f1c3575cac93c54b3a1239de89550adcc7ac993d5001a9ab54df448847e971892ec5eccdcc1830e9be3de7afeedca16443f5da29fdda87e7e690e31c65c80c7919cc0f1ee7de1353575ae7040b0a7ff0994088b4b10b0785ad67bc1cf3740175d434d45278b7420e051a6268;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6efa946c826f1d01785dcf2c611ff83a6349d1fb19d1ca5452418d06c3a3136082b7bb0cf3797ce371fda2043b914cbea4ce93ddd2c157e01e831189132d248825c7b1ad3aacbda399caa1d1136685515cd7e541ffb33982d2602a79d973a3de2d820a99bb35d7cc5c9c05cf85c72b203;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1a3a2830c1514867dc44cdf71c5b912c160f7453a421557b68213fd4191310279992c13e8b73282a32d3aeaa60a84996ec0c759b7a5727cfe0c78a54de842abbe29aeb2946ebc562bf09f483d674d74b50ccb746fdd8c6b1793c37fb1c664fd585c08c07db3f3bba36d99e595236e931f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd837de5f0fa7ce9b76f5d595dd0f22891e6405334c211edb8c69a72aab99c407b59830f0075e1b5de1b9d803f6ff825bfbd5ac3b6d24165d4d23bcdf15ad99f897577d13b43bbf03d69b7ad2d53ae0ceefa4590c2138e043b41a032cbcd5561430c414b3be445c1d4d52c2cdb98ed4d21;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc66bc5b13b944a45528b92813400538d7035332ecc04374ad68783d809c5e2587aadcab107f88b1d2ecdba03280394f2c7f988f61d7aa6e9df65ab0756f21879360f4788256c431882358dbe3e51dc804360553fffe63390f2f1cc7ce61027d2e0421d76ff4214c99c3925a959a895007;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h42c74455bc123c68776c1a09c86fb15e525e8b1a394ac71d285401608dc21692264893de313f91a9abc141b3807910f989bb4349f405768bfd931a63752051a94a4aa20d8e2f2db7cedbebf1d38548bec226fa98f76e7b2b20b67b7dbcb2fa1489b85e4c85ef5c9b1e9b436596c3c45b4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf926eefcc190924489b8347fce609626a76587069298b786b6f46fbffa77ce024ac3e7412d1c9879a48e031f3108029151076e14edd685067ecaa52f72ccbcc2a3e5a9baa2d53146c004e55811066811c9fd40d8447610286fda3068c1bd12ea490b8b7bf1a6e53c1f5a250a3b0013871;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h91f7d73c991a6797daae21ef256366bc860cfab9b5bd519a0ff8812b6dd95ae63d5fc0cc3ee51b34e2a54edb50e98f41ef4c7b970d180cdd00e6174373f8f58e219281589e2ddc0db9aa739ff9796c3c5de732ab2867f13b0566f15f1ea000131b561f004db9e29cdd599ddc944ddc472;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d43365d06916892d7a0a0dee406a6f44d79507eb3fd2c7c90948b26a52d0effab1e6746f7eda1e24ef39a63bc6b541677a143f2c9328327af2f5ace6726386e00ac5251958f6cac6a616ca327e631e42edd951090e672bea0cba4d8ca117ec7b0209d193b73dd014297156cbbd4ec90a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hccb19f463ab5518b1949b26911cec5cdbb82cfacda8e5788b48b35305cca4d89299643cb789f0e5e07435463d8134bc2c25b8c1ebdb49a19908934008cf318ef76beedd61128df6f9c131425e4abf32b95393bb615b0756e6f33976e3077bb4124360d1e33109f1487cba0fd5dc938315;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4fc6964c1c31fb9cdcf219bb86acb0f016ed74b38ef28a16a5e0ac99ef2aca4f9422562565fcde70ea59c0aa3bdf97701a239de3f4f71d99981d7088a9d15d6c5ec26ffa1ab0553959e8beed9be43b7ec937f3ad2470c5e424ae56605e7b20e90dbc3748b4484c26c5f1bd1d7e49db2e3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h815c1f1cb876935d7833473e7a895320ebb02b0f96394885078a5dc08b97c27f2aaa866c0a5aa0566d490ecbadf701784e608c097a83fc77db5b16a8ce61c886a5d71252365c11d1c8286d35628acf7c769ecee9214b264faeeec1784d444f9891c87d1e0e932957ec2621c9030aca3b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3dffb679012b1856199318568d84734e1e8ca8329e0b6145d32ee42eddefb43e54ef088045a099da46e0eed0d20af5964875d934d0e65594cf58e6ef7256304dda925dd0d7d03813edf70507222d9b3f90716e248a1697bfa88f6d0a38f17027350772cbac1be080a95a3db4370f96711;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8995d0687fcbb76ead3594b0d359de1b1ce47d409d1f3fbde625a55d091e79304a372e502e41c5bb507c10af14a5556848c929eb5219fba4c083ec40a0ae6141b67249fdedfda979a7ff20e5a6069415a5fc3fb5f9a1961a8e7b80252d9c2d43e355f2417429c58fd921ef6ddb90afbd9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f971a4415a377c905df69fae2d5f5d57fe74f24e2f88ba9a29dcab13839503c6104b2eb78b30719e4ebe87dbe2c167bda55f19622b8e47f0439723a9bfd9add149bdca0c0466a08b29343ceda8212871c432f66032a7bd7c991ef1550f89adaac0ca9e75545d36105cde7d4898bc2581;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf2c8f881a3194134a05163e973d24b60e9b6f86786b49773dd3c9ab9d98dd9f31d2d897e110945fd2b41f93c2ad3e5115c8e34cfe89299c10eecb320db9f50e7da98ac33838f7a26b3c0ddacbae70aea4520df088ab37e0882495ef025589896c262e771bc1c5ca31cfa819c6f62a543;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed14c72c7c71d2d61c627634bd2bcf8d70109e49ab8bd54512b20f7614e0afe7ad1f4137f39986b9f82408d324073775602d631878d5c4c27b70edbff40f664beacd8dba7bdfbd78499e844bb1a69561c816ba4220e9e26549804178f2638beafd9520d8040a49c7b5422368366d27e62;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b8bee85ea6b7159bb4e3448378088a028b912879782b8cdd8bb9e164b9d7da99d91931b56f246a872b93109c733530824c91555789fe335442fc5bb2a514966d132e6b6577cbf6319be4bd1e20b16c432825dcb768acc159248e7365b3c9616f6a065f1ccf715b74c01a2656cc4d7a9e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0e79e314e79d87bf6615efb2aaf9281beec54ec28c7b573d29f171d444a98bb15bf729cc24d7f1669e0390679e3073a914f9f4a4f98060f8f24cdd391cdeb142db13ddb90b203007013ead12d85b72a743adc1db66fb0ea2fa9b2ff06c832d75551da09f2e1c0aad83201c2d70164756;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbbe5d79ea871dbd467f091a2a3dac06ae7444831664d71a279dd0928133337a717aff179b10a16398afa3e9c27b2ef8e971531845cff99d11021c18b7cc0aca5b659dc3d5ca17b6ecb97a1c5d3bd583912fec2e2040c9db57f72948fe61b8202c4f3b4944882db955ba95ccc5f5bbd21e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c01cb91e448d2cad2c223856aee9cd220a6ae84f41fcb4651515c5b5f3cc74092685ce30f9058f58a5dd1c43a1b28360695cfceedf246d626316d6fb54c000d986e4dfab5cd6924aae625920c7091adff80dddaacbe0ccf70a4bdb9298069075bd62d2bd266552f7e8d5f1b420b04fca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hacf008ab0acee92afef48d656fbe805cacb9464c7c1818299cd2172586b5d35a5950be6eb85772a1af50a1ebded77b9900fcd4580cfff5391db2cc6afccea07c8178ae353b2b48aa084442735e2b70ee3756dfad10d2494ae1c7f064cb7cb3b96f279a00334d38efdf4092c785e3a85ed;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h658ebe4a681cb09713baeebc62e81097d55161a70a2eb5dbb4d40eec326c8a31fc36ebe28c8e9ecaf0ca77b5773900c00a710a7e2c19d2c47358929385145f3a664b99e91c1ea933b4156ec0b88e164b0474a305f2c7319679974e816566f67e929b8515c3fb5fd4855aefb861a0058b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b8665a43b97838b926d15d28ffb244e928a3f50a7fdb98b521a6efe7802a972b82fbbe252010d0bd00fa9ed1fb244693328d681fb2a2916e6f2865fb0e3e2bb7851a921f4dfbdb7405322f1aadd4bdef8b145e4548d3d51b3f8c67dec62ce2360c2888a09d773657cc618e0d9871e363;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h46d1e97f5285cf2b9d86d2e2abf424446fc0a84fd6a81c5b57a726cb3898a4d03d28815c160f1a530214477adbe1afedd562554a7cf7e91893c33d58ee597f57c5940ec10717de797b43a64f5385bbc67b4465da805c1402551711cc38f0dfdd4466d0af1a76d7fd9a3c4924853433ac8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb34bdba49d854d47a86c3d763b6871c72c71754daaef6c3e10cfca8b693ec3bcfed9be0df309bae37e42a8370db3c046bb0b3b318745ead425640bf37a7c2593be480c40cc88e7ab61d00708321be2a6e895d221093bf8d304b4cce1581a4a5c042d2aa4c386536acd542f21e056d84f2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc11d72cd12f683a2aac53147e8f5d262d3eed57b0ab24a5ec3a76f431cd15cd1b4da9fcb88065b26ee06625698deaa4ce251a382add3f1b9fad8415bafdc24f91db798f79ef73695dbaaa6974a446b13887ae938e37ef68931125253fa1a0455e3edd2cc317a2aa5bb87bd2e00f3d736e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8f2de9a5dee5ea2a91c8054e50a6b1435d4ce6a279a3aa44b7e9a96a12281235ecd6ef43177c98ffaec5d57cc5f9483e50cd46250d4972d1d12730556e644687ae4d87bf48b443633784cdf6ffa43e04257141d82b1e066a0605ba82d9efd9a9de482223acca8209c921f4c34bd882747;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48f6a60d6d2e2cd61f2d555513596fc53065164aafb70a475586b05afd7785d5955f238a8ea6727c1abeaec51dc373addb1ff5b6481de139a049bb5e1ad0d2971e795267b6aa2c1d873c329ef7df8848904a95059d7bc2fb14bb03a17c0c75c8b44307db42c55d23dfb0f8bfaec85d152;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3df5f68c654c4f003d2fbe343cfe8ede322588a39d82b726148f1d0dc3f2917754e6d4fe2e0098bce5ed4438e9a12976715b2c89dd1ab6175f21c83a316eaa6520db0eb7896b011b95f02d44f2a444689b8de02b3da4a59305dfef36d04b4b3691410eeb7a1ee03c1212fd4eb74b6c04a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h879e74b1392b664d64e94461a7f917af1bbe04b3e69e824df3ddae66c3268b470ba63b34544a492af597f43a0585f3a7e441d5f36e817a7d7934a4dff9b2ad26929d6f0a85cac70a17d12e1dbb663e6ba8a52e9f9f849e8450c46d84c11a999f3ca47fd8fe9f4baccbd45381cab2d4bb2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d129430b6bee1485020313b7c77cc5e649ee9fdb91825a2f572bf5196dcdbb6c834b686c6595945aaadadd87fbedad7c5c9517b6c1cf6575f1db9dcaed187ff72ecac39b42dfd0ff7867f415a3f78495c843140833715b09bdca01b2e8d8a5b2b3c3ad2b69b049d63b5f686541d3f825;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9f1de98c1c0b1c58a497804facac0c33630db7f2f5c835ed51af34930aa97e4d60fe510844f7160af551f541883a296b9d67c9fa07ff34e025639ecaf5d09be805d9bbe72e5e5ada0198b099e68dc0fee74cec034b6b012c67f1dbd9039afb61c33a300e3d6066e867ac1bea2f35bf60;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha311019dddddda79e3c77638c66fc3242ea138725d0e39174398db5895f451dbaafe545cf986f42e10d4c0221b9819daf78df9e0019171e25a96996f0f5a8a30698aa19fc22644529732875f2115eb5c211e5df6dbf39532f790ea42d1f36feb54945287bf5d9b2748b2716d9b1671c6f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66c4279de751621dedac39e5b0fbb3da5305ba89c4c6a55979c917c76be7b7cc26fa284ca1caa56a49defee27530812ef185044b46e01e66ce11d09402dcde23214e8d56f21bcf3a8e9f9913259b3024ff238b0f2f37ea54e5382e33aff7a7ae3803619744a9406bdfa7367e58a652750;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e56ed98ff73aa7d261a1e9aed1f0460f4d2e738a708a1cc5e261ae88567f04e8c019915e8b4fbf68f788426bfa1a30cf42aae8166b671669ac417b1ac2ab0df0ff0c60f195a4069418465dddf84743e2ea21e48e6c93dfcbf4968bd8fad51484526c184f873c68e798c17925265ace12;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h318b28041da00244226bd85b1f970ab11a60fbbd14479e51b5d759dec8bee8431fc334999dd9aca364e9fd9b805e811bb781e056762c2a65badd070efe3a20adfc6dba1fbfeeae2843925ebdd6c527241b7b82ab05e95ee1daaca85c7d622ee2e49e5ae2e9cebee6a0e4257d5acc1fe9e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90a0a3d31b0b8bdc27ec3a901e8b6e02e9ecc16a1524222866b82a56058e60d6390cc70b0d8074c0b25318a5d52314aeed768bc8dd9db1f552203ea8897607b4bacb191e6e4b4381d8d9a37f401ab631cbe63665cf402754764c5b1704d4e400d2c3c041a13ca13ee20f165e9f094d4ce;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h629266cf00f5f71393fc3d93f6f08dfb75096c057ecadee1a23201503eaff6657cb66c6b83de31ca95da6851cadac2523b453f1971e0e74cd04a97b57b1734fcb8ffabc065a70b7e3fb928d42881cc4282abd660277faffbeb364581df8256790de6a7cf132121ac584f2feb72bfef52c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdfe2d30843c7750bca21dd3aecef283087875887ee31c2c99475f8e1bfd217dd963d1b3ad3a662254aac907f54ede20c2794c1132c9f778cec39754ffbc5c9db37a002192386f4b20556276fe1f10c9e0907fd1be29b8ca8d22c48721f7244af5ee7cc23bf7951206d12b55e7792cc76b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6036ad82e59953ada56b0082ebdf592731bfd516ecb09a4945e8f0451bcbb6ed6f651752d211dd581ae47c5c82a6524bce04afd4d9a1799e9ac31949bb3288d2083283114dc6f54d9de81de9525203859743e7f1a1e6db2959fdd12b689fd29977c096a1a14e0a0cb327fbf274ba9f46d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54186dcaf3d2731a14381d9768d4621b9156a06d0980ec3148d78edd220714be873f54dcb87f0cda9d06279ce163dac813502e82d2add2382f61ed69b9d3db74a4aac07b31ae70c66609dfb74bbd22bc63f1b5e893b95355b7249092d7843098227ca2e167697df258a8250d00302d2d6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb91dde45ce684571dd7ab2241552fd30870ac084c433e41febec99dc4982706fd52829c81855e698b89f999025553ff4cab4ca055e35d8025f8cf0c7128799316fb0aede3d17e5e50696b6838cf15cea1c2a162592c1470a11d051921d3554ea3e211151974d6acacdc37b06f91579f5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha60890129dac40bc0767dec4b02ce6b027e65244d55e5ded15a42adc10d8a0b46ba13275610db8f81ae715ca2a841ae8ace4c959dd263d94cb5b8c9bbe30fab61e1a5ebf2eb13ea01e5870cceac6f4f4d62f1dac6603d3b545ec501bff767c1acd72522e0fb5cb68ed392c07efdd830a3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h668c44d58a73936179253ef65d101188793291e44c6bf3d4de821bc229de8daadb01f91b00aafabda2a58d018fc951e40a9d2919a48c82d67f665d9e4acabb0e9da0d8a8da81f51c51c11dba1ebe69c770fac96b8a1d9e3437004176a460e5e64232c436d0fb1ded836f45cd26b9d9e95;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23b3189d9e5914b09a9a88dbe1f9ed453bd698a4fba4ca87270dd5d7e6f551487bb2b562c6afc659666a6e8de9e5e35caf7788b46ac4a535ded54b6268cc210de64ee30f1600f2670e6652576796d81d86656a5d65149cfe996f495493cb7301d08ad675069bef816cb98af4f1fea0ce3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1e503ad15d2ddb2d72693e87669ec18611d4e0f8983b220391eab218e1b8828148bd813997d0d38be5ee49f944f658b0a866f7e58a1c336315aa171f1643499351f463677fde0a14533ac717dc9d21d930414a7cc6896ada7595864545f3b5ef59bfcaef87d6f0d45349ac164e4820d3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f065073a350fd4b313c3ad00f3caca4de779b55f2b8b8d78c3ccc86f8643ac6267c03bb09f32895463b6ad028aaa8f81e0a25f9246ad0ac4a4d841d15133ed77bf241c158e31692c0e6c84aa6d90bf9971c0d70f442c014c73709ec09d3b2af3962ad4a19b5fbe883d48e4cf3a4ab6af;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc366a8898cc9e80891384ae92659cba010aa9c2eae38768d5ebc9ebb8834c316c6e248a02b8a1d114e1c60ee0af806157c67f2680ae3919539a576f55a5db9aaed14b8847e03badb681b355c01f9e62468aed0df73c92e24f87aa2da6c1e9655f52009cc55201aa358d389b2696a92539;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83669e37c6fc79c0f8046d87f2b159211ddba5c2ca1dbf299d5fe1ecf90e3a0a4860d9d6c9140c0cabef5ec4bd185129f91a357b65426757f1b3e2ebd572d16aae12b9d91fd01f306096910bc9aa74e37323253bc055581a9ca6f888d95a3b5f3e9f94bbad79bf84f6c510847e558752d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56d519749b4bdaf72998ebd6483831334c7c1c3b6cca209a46e527d61a883cfab0c63283467f3fc43caaaa37b52ba15d2df2633cae076057d7da24212785f3f9dc5ed790ba44278067b0eee7c8b11af3544b84a667f45857c97f7be2b87c63e5917bfc84da7e2bd71922a05d12f075038;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d7f4efd966590152b6fd5be795e73353ca9183896c9652c287a6dc14d10537fb2bac670bea8445ed5bc811162ab166833dae397dc26d910e5f23736056c0ddd8ab3facbe4344e8d3857c43a52cf9dce955a626431ebcd3bc9993f8e1de9a75e092f0df32e221cc7da391f2c183215b1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha2e27660b63399a708a6ad47e503d843339a8e3da5c7dd34a37dbc0843bcbf2da103f1022beb151809c64645aee5b23951b61b531382c435924dbee55cbcf4c4a5abe556a596cddeeef90f8735b8d67adb030acef3b9dd02294b88cc504ddea82c972fde5cccdcdba7fe494307ae85443;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28e9e5a921770969bf1440849c376bc5e700f03a0a29106b8199edef0a860444d55b9549e1e5f517e1b1f75cc5de65070be961eb3ac5ba51b6dcc0fcc9ef57cc20b0ade9a74fae65a693a867083b3e62f3610767252101a4a4fe83c552c061d26f8accc189abdf0519cc29fefe0283b74;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h712eeba018293a56572a3053511bd85755aedcfce2231f59fabe7e86657479243e3a3350b28ab3ca3d2e233f8a399bd72cb7f401caa2f364fda1be2363f3b1f05b5e3d35b0855856df6cc6ca328748f481aae11a873b02937ab18008ffbd5554b49b7feba695c269357ed0f406c44ca01;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha08a4fa479a032113395fb4bdb8ce174018ca909403d4832a3db7e9c50b031d38d394e693a71fb1444507da7c17e87788aa35930ee9a727b97067d2b15015c597fd7a56037556d7cbae05222d2f42f148213810d546139209255a8222f2d9bda983bc6006520494eb2bfd8180e73cc5e2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3bb3d16c48c2549309f203046012962ad7fa824a2fad347569f2dbb295cd94330f9c94f54bb47f9a3188535e370a26d4413357ec6a104e86b5f564885882b2daf784d0d4cc5b2f5c2cf0c4766ab7b3727dd5080c482379339cf82094a111afe6bb9f409d45b9787528ab40b61d0d88b6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6d733c67f34bd0fad163e719caf99b765e62cf1d79899a8764a2dac2a67e0a898e13db760d3304a3286dedeb8cd040af1d23a070664f8478ab83e4a95164d19e6f1e9ab166381c89a3e001a63ef030548f64349189f7923efaa0a704a2b570b7cb3bab1a1e6e0eb62ee3b45d170b87915;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e37250a30b1356bcfeee890d75a69a38aece7910fd0f710c5cd2e746874dddd59bc270550cef7802eb78cca2583aac1ddbb17ac509e95adc727bcdfe2792e432470c63ca1b948c052884c3e8505f4fdb79cf7bc0611d75115b4876422600cffd27d6c03ea700e17e41453b2384a2d202;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50bac2b5ab49795c7f3dc6c7b93fab91168a3caf75f05157e2a61711df3d1c73fbafe2b10407868d19b3a8beb09a125546ccd687bd1a77d474a0313cecbed6f717ac261fb32832d29050963f717839e60afde8c5391315f2ce392930d1826392c8a96a6d7e64c8c93095429bcf739b0bc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6bed622da7cf5680d18418ae943228c25903f990a3e4186e92cc241aeea4aeb0f2b46501804569725cefe392a587bd35aa3a3deea8b9a761e576a5ed65373e5816a86b9c3d055ff36aea107eb35ad7ff228a268f2035fa35519883f42cdd39baa8aeb51d473e65893965b40fe484a712;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf7a1bb4254564a83690af3e43f6479e58979ec478d628b34ae8d94aa39b47c7e61c253c37912bd88705eb83cac4bdb10c723ad54d7952dc6730a8da69101770388e6da9f0f9a859e328a7c477d1fdadccc73f51bed7cf9e3b2b690a2b1efd002f847771ce26f7f897a03491bdd7d94e43;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h570c8c6e8a17d7844ecc112dac6338853de48bdb50a2fefa9c5b9f17b8826cbccb11cae16d0f0150daa2258f49cfb4cbab9719e5230346be1a266cf121e2427e1e5783fda4a53f743ee231a35c061076a73f69719c762550039138e1c0dba20c4308ea27f7c00a749af0da5a27fbe9379;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb20f1fb36b6e35039a25e33b3e35b1c5e8d977ac79a805c8c82454e21951835575ac14e5e586b96aa76c6ff04cbfe8c52757e0eba7939257f694abaf7d54e65bbe1f310cfe8d86ad86153c4ff89b5b7be4bec65647ebd5c60d3e319515c28d5bb5da2d7a012a1e7f2385b19c3d590291c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49bfc134fd9da51ddce74ea1052c36664ffaedd0bb9553f0a06ff773a9f888facd341b643a030153240cc5d54e94264300e74d49ada9e2a10f4eb689c3a55aa78fec2dc788278da3950f2851844cd54f4ffe0dc63a6fa863200f94901d97d3e4c3b4e0a7126be0e17bbe093a07b2352b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h255515f9a95268d6340913d33442aff39d553864c007372b4b029392eabe8fe66165d2bf47967b86584d71904bb3edb6864339ab1c75400283029236beb0f7a95f47b2e16cc26aa46d440a2c248e9a9e962ea103dc3f37dcf5cad46c40c6c17a1906752779ec50087c7f33009a54bf022;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9aa9e4de2c2c05c574a88faafc76667e433b0d752141e7e3b5b88d9cc1f24c7e45b930d1b285b748680117f6c3be040d8d8195236d8a53693ef48e2ec6e5d29d93b5849fc57d8ec896b746ddefa1c8a17c127851220a98c5c029f94d21e18bd63282f8a709413cdaba6f072843aae4712;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haebb3d937d4ccc167c721c94dfb77afb24a2e704354f1ea949933bb187979ca3439768b50138bef162291f75b50cb70ddb1f1da43b2624dbb6f57e3c860957b0df872d5f53236b99c014510f02ef401683e897a3d8e82cec5111116db55eed5e5c154377cfc044ccb470f1ea668b66578;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5bc3d6ca72cb4fe2d9ff5cb6ddd729459ec2d0f03b7d9b37ed7823a457bc4b0ea6f885d0d560df9b48f2d38deec72808ca47af767c534388d69d0c09ab96faf5bfdaf7ca42aac7b913611454af98b237016671089d3ecf319f80f8617f89b8cb8df9c1c9f8c5ecda5f3eac10c13beb81b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26c4b7d32e0c5ea9e8b1a4176fdf1f40ff0e643a2cbfe4a95227e003a0d8c7434a061e9da77918b45902d4a4283eecd7de9b78af203f9593990b352f46760c9ca04935b149de6ddd97aadcc41e85c797c25b2e5be3ef63c088ca33ec93c4419c804d28a8a3b602a24ac3ab705bbfcd471;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75f4cccf1a2c8b69897ca43f8c72572f25a55da3dfa2922e2e8cce067ee8f5b6e310c17c41400f972643afd12eb121b8156a7e16f306431ddbca71077581687e9e7fa13264cbd0b3f472ff81f0dd54d4c20adff7020596198e54ba52d1c50be5efd8324b953bbaf789b0af38ce2d6626d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5eba38524055361c9093624e6c9f9e71beb191703a17ded50d399e2ff6a93ade3d8c629fd1d7da3f8c6371fa4e88013066c1e49a384ea877303c76ef44b7e86a68379dc1916b44b2b96225ca011dd110235bb4ead9e36b889c18937a1ffb0b9ca1a8cc22c50d9619cd615c6d4a43ed06b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47739b1067022841df19606f901af0b23543303ace1d39ec9f913d2bdc53ca7e3ddf6060ed43e07dbc1d19f4c1430260ac1518fa8505db60ca2abf89c9542c6c80d7f0a28c47088c560cf56c3e93fb138588f4aae6e90bd16125c5312fda473dd5c1379c80594d265572bf8e16042391c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc0fd9781513ec7a81fbce6deca275edfeb8089557daf852072bc88ac1140f4f95dc6e542d9000c0f2353790b82ef17e064fd493f5565d0b3fff683e44e21bb2f1f693898a317905a046b3344be35753f32e8dc8e3b5470adb198435dde764fdd7c1e67256bf94edd6943c71a0d359a38;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff6b7bb6f93278dba5ef15c59dc00f50f2e142831e59c3f102d3fd021ce86be3c7c341f36b452f4adfed42a065871aecbbd3aa86e853ba57c2eecd6c8b96892bbf5463d853a3a3ba6a659efcd42613ac3cd7e0ec2d31411b9c2233bf3ff44d3d1beae5d187106a0f76308af3c24ab34a1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda1a1631b6b48b57bb62fc2d9dc3f3be8fca0d9148ab35afecf42073b4b4fcaeaed60b95743ab3d64696849487580a537ef4165ea7a0019f3c93f0ad2bae182c5c3d00e18bbe089c53bf8b5256ed72d6c2f082d3e95f466c024d75896e550928b3d71cd32004abea681d9845f0af809fc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32fcd52cef601344daf2848dcfc21724be12aa3b1c86a2c371ac795c63091849be6e4b0a5bf75dea7876737b8719a0d144ab225362c802ae102ba3d56c879df5f696320c14f806734b7e699762a222d449dd86e1d542e7686a99ccc49269d8f33ba2136a3510691224377cd0078fffeeb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3872d314ee47619a0805520d943f730c0744ce765725de00f4d3d1039dc801ce381d0f068da22bdcf7e0e1b54f46ed0597a8df11d167e76c32d5596dd9443751c9c87d85e4ce74a6f9af30091380cf5d8058438a499247300c0cbc4ec7e649e6c9339608a661673f28d1269caebe0e49;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc2adb1f8199986b3ce1920a4572d3411b587fc28d52e7d5c438d3e0307d63ecf12197ff3e8d8c47e4553f36669032cd3653e3cb7ee9ebc9b18345ec8b3ece2d3941e42652b291ab318db3ee9c0e1387939c3cba38bef497c6982f56ab74c9f51b6471fcdd306d38ea08b9d70b293ac77a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90d6acc161286868e4c11332b266e5218cc1d42ae7ebce5553eae4d291ff561f526a6f837640802db08c8638e80f9772e9500f05fbb10b2475735ca30e7b15b9ebd8284cd3184cb0ac9dfbec508b535cffc0d49152b69b15738644596a628ef61e8f96f8a082800eface097a4556b62b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdf1f94038a335b7abd610cc5f091f7b22f62960833df8ac00dd215674308a84730a353eefebf07d1942ba889ef7ea25388e9f42a23e8330b6c883d4f78cf1a47491104ce21f8457078ec6dd986525650dc5f3f28be05be27cfe911ced9cda159b894c5b49f2d52a701a32fbaad27506ab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hebea381ee2a5c0c3083006cf267b15f9dcd2111ca535f41b8b70a6692e7604141253fab4cf039d38c336644ce94e62121fbea0ae9c42b7358763dbe8f2a1546321777f0fba21645314ce67b0ddbf922983292d27f82e123ded4e6a8b52f38aaa374af8fabcfef5c52552f8afe9fdd2c2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7fa3aded4eb133cb0ec6f612caa2732cef6e78cb397d797c403d0135e027066a4665fd83d1eb4fd21e9fb5e937d53a736aa089f0b21ee0e670d2851b7ba5e89e6eaf09175379f1e088956b1ae87f5558db835a32bf9107f091e33da9a3d230d05f74ca48706901c52d73e1d55b47f980;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45462754fed6c81a7439901015de78ca2fc1ae8b5a2ba702f9883257d4868af0e3f7726e24c35350ace63c330b85d0db1b3a2d935ec6d901a3cb562fa98804d4f868d062b5fd55a2458d00d43c32419b88ebede79873ba55af3ce63c68fcd5fb1fdfb22f2328397e8a40dc5282954ad46;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96769ee3e4e77c7fdd00f68df31db20faf48e2ca6a1942dcfd6809cfb0a6087bd861d1a94d7aa45f9e03febf9b9d9d074fc03bacd2f9f2297c09e3d87e85f8d663a1f97533dadf19dcba35f14cba62cfb428b27a3b4e58986eb3324959232166a1d8947524deba306c30f4b6142e430f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h983a95cfccc378e3068c69bd9db77400fd23cb64e530ae53f17cc2af647b2db4397b7e95c78acf1a3c25322e3cafff3db576d7472f96aedb0160408d9c4db0504b6db418c4cf92ab90a60925833ece0d5514382b9a45db4bf803689df6f8555f3a1ee05153e5c818ee5267bc4f487ef7a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd776f32a6f1b8676e7cb0b913fb8cf67fb31f1c98c7fc34ea6e95670820a4489fe722aa160d5f78d9416092abaf884a3d026a63565871dc06bab4877ecf705b3cceba6cdf5ec048ee6060906c22181ea71396a7de7f328085e80e879ef49a453821fba8cf28cd08e536d51e6a83530e4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h780925d914656a07856db319e86441391e8b2e54ed1c5175ada087ee143f06ca067faf35884d830f362cebfc8fabc3a274f1d96b962ef6ef56591bd1c7d335208119b74474df7cc9107ed1d172ff368fc126a26e367411ed21c4bec25359cd8b5055f9fa6d6010b9c4780a0a5cb4d3351;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a4524152580f04ac3397529a84a8f597b3d9ea21d434ef0454f82deb2ab5f0d0451ce0435a49ec489edf78af4b9e99f5b1da57a1465d2156ceb10e21f95487e4636e79607cde7cba8ec9f20e2e770053314a9a4518802eeaeb33815f8ef11359d171248fbbfcd59aee9ec905977be161;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc707e5b2a14a3872aa62e2e76ae0e58d7b5884bc19bf00126c8ccf6cd21140d9ffb87d912d6f4cc57cf296cc1b1066aa89c70a845b5f9bb4c0ff1202f4dcf00874fb026f70f64d2791a344db8e330506dd5f116070bcf37c36c293408cae6eab7d2a19a184a928672e586ab932bb9f65;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3b6ea9b0e5540ebdcce86948b8264faf0d13ffee674ebf3b3f500469475c794f210ba5b47717263331c93757d97ff0890de6896fdd0c1c786a3428da7295a1e0ba047b3f00856828897fe43e4a0d5b4f53c855fcdb7c92256077d7fae6295df32713e4651931278f7e541e18d4c701a6c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he20fef9012dc49c95f4a108d034335f9e141eb53a59fbc1f7763aa3e440529ec57dbe537a65fce9f5a63f69e778a7f2803a719f4c81d6406d0483ade1d10a4dea3de50a919e41ce4a68c90a751eba40f7f8632a3dc5b6327e42a36ee68cc1cdf8d14d1376b70c778b71464d63dfcf77b2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9df8be1915f00903afb5e0d16edccdab8ccad865fd09bf687123b3b2f6645cb7d60579c6ba028104719705b88d8272f061791341b7552c9bf17e2a42346f7aa99ec9bfea85cd512753fc7e64bd93ad0a832acdde7904a40713459fc6cf0579cc7101e70a42349035469ee6507b394f11;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfb4ac74dcba8f3343313a3126dfc57235c107eeaca7a95c3d311021a70ec200c837cad45bcbaf7bceeea468121d41d74b4957c15b975d63f68e8471db2bb6420e357670095619e0ea8dcc605a5b090296bd94e55c1032dbcbd9c5439bd591669cc4145951241a0798aa35765042b497c4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ac156ef006844b0ad553879168b3d5ee606fa8f11c0ebaad4f5132d716cad8c6b589b66cc7df0180b3207fda6cbbfb934d028ec514dba9301ed393a01dd480a49aca9a22711d6a34ea8b065b7799eadd9db152789d9fa48143062fba5060bfec7eefa501b38ad6780db014158c2746b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43d88fa4c71fbd3df0a25b37bc171ee0c801a68248bd1c64eb9e8e8274939b5ebae386375b79e20519bc50ece953474ee12a212facba45837c5c773339e1b55500d5c749f6caad9510a48ad42875ef568f77ec476f8c337f4e132cb0fb0d1dfa96e6f83ddcbe9a8e66fb41eb41553164a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ce63c3d7f6918c21131479b8bc2f5d96b9b43ecfe6fe2b49f54c31a22e0ed12c5bc7e616463f086675a742804b8856eae1bb1140526770399abcbdd4aede853eb154874f577ee7f953c8a15ff2d479b0fa0f83084f85a5ae144693ffae95543c1b5e261a1bf484027bcad426c57a1a2c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb8b00176646013e48cc2390144f4f91d7a95a852aa4a4a50554998dde35f8228441a7bdf906c1df4f52fa00c5367f7df86d4ad0780ccc92ef1aa8f15010595292e34a67556560bdae99cf31bdd6a93ca09e3ac08f51365eb47632c5c054dadf9731f52bfcfda2e4eae9347f08c192c41;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5406e7faf2a1a3a5694dcc8ba8d398d2ffe883afb4b9411c7fb632542a7cb24e6d96b34ccbe19467ba5903cf9ea06c76cbdb76681bd287032bf0dd396d071160af081436567669227397f0d82e83d4e88e049c310778023b518db2f16555fa747ae53ae9637a9115b5a2a8667f42e1e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90f520fbe3476eb955a2ff0af7254968bedae9da572ae866efa3c97a305de4e356061b264d169711900388596b85f73e7b0ffaaddb34dcda6600d5b621274cff54488078fcc4dd8aa32a61817103bb00bfebd169abdf6b44122950e1460f923c29f416434fc123c37dfd719b953adb373;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2f7265adf48cc845e1e6ce7122a9aa12bf403738558afd5c24b4e677b1e0db7110fa7d565609567bff22275a84a67a63c64121fd9bb464a52e895a703de724a39f1d4239f7197a000ecf957d21feb39116afd173ea21da023781907f8aceb3b693d188a1bc0c3b2c7ad94e2239c6deccd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1783792f4c70b6f83366ad3981f45c1e40d4207582781dee3c7fbbb097fecc96da2a45dfa55de7177fdc29e2ede11be717e59fac40531385a9d9777af5a9cf47da81388c3ac481664f41fbd00af3b6f084d6bbd2365ffa3e4ed1969284270aeeaec7bfc8bb165d36d8f98c74210479bc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h77684ea5b1c47a9c1c59ae707f53bf2bab94e60b41b765200dbd6abf32678bcd6e015bea4d207296d446ec497c5b0701ec3d59f9a35739db64e3f7123f1bdac6b819cb3d1a86ab21c939605352c6c6f18718eac1ecfb2f2b0ef3ffd2b6c1ff5c80a2b521f25250987fa550c778df11b2e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc97ce8cd7bf156a8041cb2da7fde41b83b33cdae1f468a2822d9fdc5412e2543f79c7745d197f01dc4b2ec064c86ad9d40435fcbbb43882a308583e704bef62594567b0c6b44c3f3bea6d3b6867bded236b76174a6967af3a59a2cfc59cebc0b64c97b2d3f65564033851a7ae8b985d87;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47a89cad36e63a1f205994e0f0017e2d8ff38dfe315c5452cb81a06efc9243cd1dbebb4e7d7451afebf17a009f0d2606107771a925f4ddf64babd9377ba1d508fc8c874cec5fc9b9d7b51d86edb83ca2f416317252aedb02ff8c2d4ec60d2da9ef0752076dece0f3e263d514cb97efda7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h27b5cb1a8a652a7fe3fa8d2b0c8bd23c2dbb48b901567ea24a100afa7fde28719bc694dda24be06cd9c09aef21b222098f5690bb398ae04b1fa3d3cdbb8be70965073452a60f3696bcdf521ee11d56a919061e16a8f941d07e4f31ff32542fd3dd0edbfd57f35d165f98ca774fbe265a7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbcc96c282aad211618f394f4d32bc8db96881f7b836ef236344e41be0c9560e21789d65a894bd28e38b88775489003f98e827dcd1faf04c9074d69690062fb0c77a8d29a4194fcdf7ec453c6d7d1acf5948da4a5e3adbd5cf958ad9271859add65b52656b2b6c8aa6e6f234cb4095aeab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h318c3f57337f8e06c23828e8475e5c96de8d04b6edec021e39df2e6b6fff1eac0fb1e0cc7aa0ab62b30052b1629abfa1da48aa961d1f918c7fe46fc36e3395eed9c56658ed1b75ae6697e5b74700e3ec8641a856ad0d51164e479e41c33fe79a102a5196de60f5494f6ef42262c6400d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf939c733a7c204e59d22545146469d7c18a0a3041f17d7c6a16b551de8508be97297f2fdc1e81d06faf008d6c97fa5b3571978fd2f054ced126bb6ced6015f2ec84922f5c54a3d3f1eee791b2ec37fc471514f854b78b634f8b9bd484a4fbebc5175341f4f102f66e388cddf09e5ddfcf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b5ec0c9e79eee99489f58d36f8ed67c75fd5cbb6d1c0f563f8878940cb5adcba616afffef5b2c643a6d720221be3b5c5dc6c879e77571f703cad35fae5359cf43c27d2b33517056547a331dc7eb3872bdaa4bebca232d14a09a87ea121f95c30a59ead2d4c842bc99b154e60fcb0fb36;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d4bd35ecf9b896a3e69f51797c284600aa6d829ccc710551ce8a825757ca1eea824aa0dd9e78842404756349b169f99dd7e0c3df6f94fa76e4e71f52eadac6aa77fcb4a2b19fd2a563aef66f9df35013067b9d269edc23d97ce136acd18454cfb26a1a6961f037e9af163cceee70764a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h74434529e8f15793a8e65b00c6cec373efb62162415f8978fe77f924dc6d67a6502943f201b26abce6873c81f61746b6406062fe746d7df068b1667430d96212b4f6be73c2d5018cfe651cb2cc9a296f911fc8fee688b375dc1e68974e441b3e56faee6bcffddf8a23629abe0c7983c29;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88616087c43b6e748e2babf9fd7827f92241cd1783d0f5e7e2844518702a3fe8f254517e5608e9bd61898697cd01f1a051165e6a76fe0e95c0d64ea4f931f89860daa47b254fb659f43575fcacd95ed8b16c2dd026dc7451076794f060c810292c115322a78de635c33ea487117a910ae;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6575d7b2c5af94308ac52366d663f3a6d502be79bf0d013315f9b7ab06933829b540d16811575fba20b9927d8e4dfb1f87c6d584b18e4c4595401644a4e7c7bd212a48375c4a6019285a46bae29e049a75085b45e9dcb24b9d712d8b70144e6559f86b47c99dc8d985e62088be764fbb7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff1dc9397dc39eacfd54611bc3f2e1780d3c13cb9f150bca05c262e39ff4cae76059aded6528ec06a3f2e83bf06be73cfb1e24fcebd19e5f6ab8b3fc12af206e18502c26cd3d3e0dddf27c8ef8a5ca830467fe7059d31238691e017976b85b8b07af7881f464554b3ee1f6e20cfc4a99a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h23e36e52787646b5d8d1f426170915f649c13422585e916eafd57064ff20ee5a19ff0bedda7a8703144dbfc7c5e41247b259e64969f125eb95a18fb784691f0da648aaf605d39e7d6a4b6bb907c5fceb3f8e437fe5c3d922c62bfa298dd2bb5d113f7176328637b1db3fc534edbeadf18;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h290bf5666dfb096fb768082e799437b4a101bb095f8af67c49752b25b223b07d5e4a014fb80b1b3f06828d1b027fff20869171e97391ec4e48adc858517025b8920d16e9ce314b9f317dbf259932a5f10f741e6b420f65dc9a2d75b2e28f56c6cfcf816364dfc59dfd17110d1ba796e23;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe40e47796ddb2ebd18eb1ae1de36dc9f4bad80560f33431b766ffa976a2b13fdeade7db3cb280d765b5c6a8cb323025011096e4259710b46d1a9e448ba5a5f324b739a76aca5ac836f5e5a1eaac57278340ed5f5ec59fc8d4a8dd471784ced449d779bae1e0ba4857ce0fbf96b15b8b4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed90361e3658698bbbdbb1e0508b7fb2a9efd93ca2010a626724ee7bbe8ceb28ef8ad0514b2d88adb353fa6c45659383d2091ffa73484ce2b9378a27e046ae99eab3a4d360ea373e492f0c03d0c9d5814805ac1187f9e2d3c687448a9432779deb06e5ebd2a9ab397fdade28afae7eb54;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ab2d2ab70ffa0a8f5bc849e9478321a3b8397c51f2f7909eb9841de0e54ee7dce5350c3c60322f92dd751e4acd836d05e1382f5e572da14b1864b2e1103025d14a99e5a6cc5cecca4389ee26fc6c34c215357db064e82324b01c81067a9eb8ab5b09e3f7b678fef55638d4f913b75538;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fe1b570728342e85e8a1d09adbb173e7e4448f808ec5f3919cfe54c5e2279175b996cd957debd57135641730470969c2d74976496062f972a6bde9f067200bff542029d15b9165e504106b2cab77d3282bf30618b7332557dfccf3237d6a031a519d2d4c8fdabdc0dc19ad0232f086c6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf4348eab110553642615cc170f9aca724a37f3e4942c78dfe545f028085f8d8ccb28e04dd400c4f692d26af3ba897f7fa96b914d6688b527dce5bc6916c28c6c79508669753631566b8deaa56f8068b2735e5792f52236e71d03759446055ae42f5f0098dcdcecb4d38ff595e0cd07d33;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4170632c581b355877d95acf4e50ec1a7492fc28b323399585cbaa1e1d003cb956767c45d86c1595b035e7c056d91b2c6a3021e71ce6d8e8616f33d868d8f60d8c623acb945babcc2538bad53a66d388b22aa48b77eb99815d5a52588190b27af6fdfeea3bbd7e1e4a559d1ad95e128a0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4881d25c39bd7d8cb3640465aa428b1c537ff9b650f778dbcbf128354da7ee569ad7273c23f3746c3f7343171c2d4cd01699feb9cfc05a39d124a909d645297c278c60c6e5a4cae7f8217eb7665054588882fc413eed8b8b9ed95e4d03e3d2159fb1a88506a1c4950eb74265ee6c5c627;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf831c333d4339d3ba1551e013f74930008eb8019458b96e63c70efbefc415c28ed5b10303f3bc36c4554d3194b7a587afa4c53c495ac3e89dc09bb061b729000adfd0d2c61dbcbaa7c11aa340a9c8ab118cb73df9d7af4745b78fad6a2eba4a358dbfb67291d8a0d80fa5bb2a955e2645;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h34743e70ff52d691c130a6b0950c0fd28c8aab2df80a4f6a2e9c2a691df3e2aedeb9387eb749a7669a2bbe93358beb692d5d41c3602e8ee69a0f76ece60a70eebb61d239cc6d5b8f9319c67151e8c1171753a6d4836361095b30efc078c17b8f0e12fe825a951920e4db4534a0b2e4806;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45c1f19343aab76bbe5299bd8deb97f80458937310041e82aa7da354c20d940092909bb0b0b86571cd3fbc96c765c3b377ba5f052726588e822e366b1ced6c9d6261baad7df3e96e797da56bd63afabc083e54669cb6321187e642bc5dc41e19867e3c92d629ceb6cc346ebc5d53404c6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf8d3ffbb06a692fb475b6a025b7fe2c9e23f2803c1599da5a7802fb795dd3e24b50caf6e5b6c1a6ff384b2c54e07e2eb28ac9a76d43ff90f256b91130530ff4137e900c4d85d4bc91322fd104e9d89b04939d4baa6a2aa382fda198b2635b71264aa09179c05cb280e7fc1054ffd8a77d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce0dd04380aa9feb74236b9664aed66910c65a383712bf723dd1609ab98019dadf0d7a21fbacb9f15708fd4eedce2c1e1b36549d9b7711cf69b36560b3d319c29434e0c6d0c928cdf155fa65c7d8c22e3d8cd7f19baf8dd8151b833449803967ae62fd9774c55a286c6751cfc3c49d47d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbba3f5ce0483edec9f017cb845ec1ddfd9010de372830b5bea7b6c908bcd41704c7c0f0ac5bd4116880daa23925894d9a04305a615b05d39999a77359a362737b588008f244d74df638090637599eac8beec62a2c1fee1bcd8b38cf8db240e7211d8c038fae235a37a31ce9b1e1b1e961;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8594726158118825f1ebae526cfa97c7d1198b7fb0908c321dd647520eb3e2b35601c3e92789b90c64722ac658279eb54ad833cafb9c48aeafde3f939e87bdca10f0d1b4cc8bc89297d6c3b089833741e8d6b8c32fff2305de67fec6eab1b09a2b64a874b444ac57cb4b2c85d5ce0b859;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14304f84027750b41ef5288ca6b102b69cf1f41966a1fd5edafe8b7a5cc029c3f7da6531d9ed5d0ad4397e80cdf291ba80a822966967cf229b60cb08b4ab519cbdbc60f3d793e6a599d1f57765330bedb03ba4f26cd0af7dc01f4582e7fb3db6cbe0cee761392bdd0484cb29fd76561cc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1411cebab1b9683ce81dc2a2a1e88723b309ccc4eea44f74b6111c479cf85af9d3ff0fc360d5dca84aedaf3fba815514e6374d6b01c4dca4f0f286b447432dc5b96fed236c95382b77d4f021dccfad0da36f267b42c052d7cb23cf875a72e041b6185d365c8571d1429646d4443b90c35;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he33675b073b5eaefdd43b041e1bb2f6a13d991e5d3885e1ec242db452019e2072d1ece4d2d6e031b308c740e753b08894b405e3626dc62729eb2239b029f22f08fdb0e3b5ab6cbcf581d3f83305bcddce0bf863f3e1842394952ed52aec404ae491b7682acaf8238923a387e3b550038a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78162fe6c99dc04cc3917b5620a18625428824b079d1a1afc1e9c58d098a5845b79e9bb65462a991d7643e4c8970c33bbea26b02131eb774db4b4d57a55d72e01f1d69c1746c61654fb74505e937824f88135b86f9edcb89d98e1987861d462aef3e5b249fc8bb2f0eafe05feb4ed901e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b5c077c6f70a6e19eafdee991b21bf82016066ad88ad017c6420c1f3cf82a51dd638bcfd74c740474b4b00c0b2741f7b9cc9e538d7a0d8f7df222f94c90aeea6b4c401f6949deb311fc3b467b85a621690b6f7cbb19671970c3011f43abcf24d9ab36432745c5242fbfb58168630c439;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hecc00565aa758e91fc5676f6e39c1a2e51e25e171c589bdc61fe29bfdbf826af30e54cf4cae1da57dbfa8ac5b6772c5c2e98be2ea053df5ce713c6f7aeb1c59248ce2d826faef059234a7616931e7a8dc606d433d7741b33e35c5c4d25031d9e9926495a82dce91990adb879a9bd70e97;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9545ad92bb9cca1aa5029dafcbf9d71c51d41fd522675c917d77a09c65cf6345d5cc8b3f4ef4ff6b2e65592d677b2a0aa51c00a91fe9367080a05c8e639d98b825261e36a42c3e4cbdd0045fba4d26d08cbe3dfd2e26e0e7ea999d4270e8a326b31dc148902334bd8153d24e520deb436;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e281553b65f8e62fd41446bf5fcff1e565e5aba6ab0061ea264c0b3158830838ccf59db4baa2f3f810fe73a754434610202d473c582d677c41a36be742e93e5be4610d2cea92c5db14e425d0bb32786f1c2290edefc86130959548772e14c591d52629c706f74778386c1f38848cbfb8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb4a9becc0627836dba4033343584714b1ac29d2cfb35c2dfb8e097b8cda5f6b3b0f37a939b213e3e429e968e1a30641db95715d7477328d9ac51dc1e32c02e23ffc01385041cd1187d084a77c395a89ae632bf6dd339ad10ff47347ea592ebd9e78d4fecaad2e5002f63b2905fbf8d094;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha6e064e0b8885681cbfb1c047d5222cf9e0d343e0cc9f5293cfdb339b8c7aa2788ba91f39a84d18a339d68fd38439bbe8c89ccaf63f1d51b88a3bbe66d71ccb3ad96edcfe465bb4f7634f4150596b8de496979308822bbe4afc202e626b42888cd182e39bd87fbbf2c1194d961782af57;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2bbf0bf85da40700a14b76aee26e95fa3b597b9fe0b83aa78d90602dc88b56f6b2a41d6f2fd28d9c98201783f28931f860f10b400111ae56a0a61f2deeef3b3a1f13a60ae109f4390cc542c75d027bfe1a799dfc0b0057eb48f3de7191050053751f0e7d7cbc59947418d7d396f2321e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ce4e58699c8981d077d8e3976f73b9181cba7b626a0c5979b825c0dd3eb17cdbd8e354ce6f4c7ebbab0d45c15a369a601ce45a0d17c0cd72e1317fd0a1a39669db63460c7d6bdca6f7e75317940bba8fc9a0fdfc4fdded0bfd54e3cb044340e160250e84e6617c173dadcb141d48aeff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2054a2d1999b364b0f6a17a5db834e218c7582273d2b3ac84f58448bcbd4fa3da675b06f113529bba7666c941e34ffed72e3e803ea9e09363ec3d8a01253460a5913eb6c7089a4137fd3290fb42ac3b50148daba076d19f673dab7edece960070ae1abd70c43e67e3b9fe585b63e1061f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2e00b23960849cc656485cdaaabcd311209793a05a6447b4fd89c7849a8088c9d12c53e10e6fc0221739368c277699f8d6009464f82203081e2fde1f0a2c51aec39ea65efe4ce32c0236d16de033bd0764e7a819c8e084bb08101c32f576413877b28a2a21cf759e235b71f0fa1cc4b61;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64a10625cc33f9610e89bb87cd2d3ccd98786d6b3ee1c451470defb39f8d65d475e5241eaab9630548cf2b37f367913e2f4c754c25eb6de7bf4915f89de69e234ccd4e70564287f8c59771c72c008acb8466a4077a488ff10486843897815dab4cb3054026a69e5c5bde33653967723ea;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h466d4d9d12971a1de2733df68e218999f4b907db15cc5d9e111fa22f2ae2ed4b0e7ff3fbcce63d2a663105270fc096cf7f340ea8d7c01428b93e67c557a6ef5b7d43f966800aa7e60e52c8781888e92725e7dd3d852e272d45cb71d015c0e1ac9f9a61ab0adcb68bcc64c7ee2d376d2b7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5270fbc5c515615e484a455c3a3b7eb98e80c681c5612bebb32beb4eccdbd4192ea6975adb92685aa9e9d0b3aaf58b39e7e43bb1d47a430ebc012bfba59baba50b91a9bb2dd63f3e4a3d5bdf229bb947923f0ecab021240916d88035c980dc86efac8358b988eba0a5bccc437d916986e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e03d7f42f8250623f9e30a4bdf5ca3ed1a3693cc3f25a000640380a9289872ec620d4f0f1dae40e667cbcd0d6d2ce8716450119baee8fd90fd5ca67b233952a75023edfd3f23064d2d5c66e15bafdabee35fad3f1622b3c3ab0892373c03def1e2762ec1365187bd3725717f7efc969c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6cb9da7c13ca1dec7a31578f4a26a49f7e33ac16cd82b39d06b234aa6e6b0b6f1b23fc7dabcf28bda6bd3ad1b51d906c09629c95208cc83d055dca4f05c2170ecf2245599e3bb0f213e259ffa84bbf1fc5103730a4bbbbcd40bf8b5528b0551811de2ecef70002cd466dc27f41633a504;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ad640f4ba5e124ef47b960ce0467ae120a5f6da4341364b09f3bcbe9d05b783468bac55fa1de0d3586b02b0029d9452adad1c398ae560ed73d0895d10c6cd6a32d4cd0f8385db2165fa1dfb228bf4f208913c1fb6e43018184e193082d01aaea9194216c614ff547cba5a07680789753;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4709a557d62a42f531a2734fca38bd8c2e84b9cc1d2c3a8dea8071de8bd4183fc4a7a6726f1bbe4b2966480ac865a54010dd6593c326c7e4299b8e4ca36e566df8602efbd9b2b97894fe37d3bd08723c8053c4d28dc9be88e6fcfe04cbf860f2394dd79f7ec14c9d933a08ec607cb24aa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17c0fead276e40f9b15029924c1e173e065cd205d4b8b1c6f05e9882b4a6e71cbe9bcc79b39f267ef049d2eff0a206e45b53967789b5f9d5bfe8fcd24243874eef2d68e6abf3bf43a9356abadc689df9d8327fd4b8e8eaaa6ab2c7082165fab048276a51ca419a87aa7ac18be8ca0d914;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa6d6b2ce737fb600b918757b160c1f5f5064bb692bd14d8be0d209f52a9543afc6529dcdd9737cc313c8e8ea21ace7de1fbd965c421cd7165bbc94274168cbc85b747a7c9c6cc3651bc82b2f7c54d3f33c8896ceb748d15436fb9512774b8f2f0bc86cb1996d57cccd2c1af6064f71;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc3179c51ac773bf4916f2a0d418500068632c29d8b8c23e06c93cf2d91b68d3a29cd9e1d16dd5a516c879326e6db379c799d67c2872ffc3899105663a2b6e1bf8bbad7f5e934210fa5ac3aedbc3f7f0abe34fe16783f7dd15aecdbddb6bea4f62f7545a41bc09d824f3ac949dc8a3d4d8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66f5c8dd1bf7251e01ab0ba93c99854a4f5ff9af170830eb465732c6c525931d476f97318ac41a432f0f02a54d4d13493076da7c1acdd4319644f1a74d217397e6e9eed94497d4aa37e1c99e8f4d575521843f81d26e40c679ffaa752a964739b1b64e9d554544da15b2368e661d3893f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d14cb5dc70f57cf7707d3e8d1feda3f04aa7838d623c19565d1a7ee318af0b9ffbe045f003caffafe371112f704da8a1b7ae5d267898ed9a38b935ee8acddfd0c892147ef73a8d6f6f680eb11cbe290ee61293c97bebf606b5d683992489b771a012c198d8fcdb494440b231fd88db23;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc8e1a805fe70355aaae8f5a371b46f112065ade735e4321ac74bee20c4ae419c126e05cf2e3e6388b7e8a2ea9f4d2a5b39a090ede1b08e4232bc950c5a133b7335a23edf2e573b4bd241e9f8289d1b989ec98125ae20805d675a98d7e7627baf0d3312ce2cfb1ac1f4871b3d066f2899b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he6256ddd9df24dc2b3985b6fd3ec1de3e43c88061a2c43e7604dd4db28c608a2338cfe52056a126ca7aaf01912f6099083ac9672036297664a1e7af12dc4e60bdd19a1dc832685a564475c19cba18259dfb785e649fdef17f6517f4aee0833e45f19f729ac2835101dde4f034341f33c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h167069cb0a22ddd053ba5e71f8f04dbafea97b903837a73d7d978d8befbf9930e56bdc508c45c6925618e41cd4ed5fb7cc31256e8a5104f429a43cfc30a4ca8039c0728b341ba22bc947add8dd695bcc53ec4eeb010b3038c634ecc3943cf549276b077c2d562e27aa6216c20defaf8ff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf2b9ef37cf8696422ad4ffb65e7a9d56ae451fe5bfbce1d0a6915909c859896c35673eb9b901e526e3d8ed93ebbb59c7d6389233be7560df62c2ca05be236c51cd9b4fc95b92b151349287f39249e0b95bfab70adcc780570b7c54a00f0e87e1b3e7e51503b4cfa2195d17a8ec3a041a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h72bcfc312eac7592aa5fae59c88d2e7b504bc9ac74aead340c6d6324ee8688619c0e77b5f68c3321b2dc31418058093ad0243942d9f3e147504b64b1365fb8f9a0652f82d881e16c9b428953506823854bc1bbbd2091a8ebce0b913b1b859f16966983276892f739e795ddc0c8fe3c219;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h521a7e8c47a87c7a20f403bfa94e825e751750a78daa9a1be43fde74e04d77e32fb0b0a08caae0fe6622274144857bf5c97ecaee599958ba9aff0a946050918d047dbf08d63475bc3de36e3daa45a2a07ded52f940110439bb453e3f5a9648d47da1deaf3b68d8fed01dc0048de4bfefb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed1e3107f98ff8b0511e086d7dd4dba0d36dcf7c72579880596d24d2018f5bdb002beac7890f336fcae63dce4c44ce6fb27b5d6300ff6f0fe844f5c3cda449c5b21b658aa440d5a43348cf5ee20ebeb04d1c872441d1e6e7c5201c3bb5c8a80e71e8d0cef38b4d388b43318631f4ae16a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10aba4a7eaf1041a2edf5b771a7b95ca69fc3e838b9e127e82d605db1df036fb96fffcfc1dcefbd56db8a2cde811e0ddaacdf890d3dc9f391d3daa7bf7a7aedc81971990b54cbedf3c5ae4a0f7fd62f08d7625549b579cff486b475d786b6be6041109c44c132ee10738e4366511ed862;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c5fed6077bdfbb1374b0a49cac4f5eb20d2141f1c43a59fbf92a7edf03234d1f77bcad600b4a6c4c071e97d99736527a09b34219b193068641dc3eb86721a47a95192639838f3ab50fc6319c403d5e7ca7eb488aa0528e145e53f6acc20ac42333ef7cfe18fe8af217031284b8230ffc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h112f85f28a5ea5445ae6df2bacdd8d6a5a03845b6c16488a73178394f1d4c286d0482e3dd95b786195757cecc35c08987fddd121e77603dea389e28bd40a99aa86a3f400466251991a60cfa6167d34dc0d2819c692e192cf0af3e3a6f47ddfb5105e94e6c73bab429eeb6520cc7e15ea4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha68ebdb8df375229d8bf2f0d7e3f85485f1cc09d3a2687883d455510ad525f95ca253eb6e3fbe10fedb4f3be148d287adfc427e9d60b646dc30127b606bbe7f2addcf25237182d199571979e6cf71b638e99f211560463bec21dc9c7702381ad628922ae9d788b1d4fa1941554dea6582;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2540f57ef2506c9828c6ea285f3d0bbb8d637dcc9e54774af9fca3ef4b812b1587c9d7b7b6e840a7b2e76fdc774269e29c1c6e351da7ed252664744d76ae6aafc619ce63dcd60240d84b0850e90fc365212ba58c2dfcf839f6ef10d38ca09ce5b579f765b910a780c33f0c11baf2992df;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hddd9fe3ec43ef96dc243c423a7c55ed3999780fcb31450d785d526df26983a8f54cd6348877ac48536a75eaf3ddb697dc11ac438f55b703faed3a1e4c718db9752d9feb6c9823ffb6e9399621776b631e8b7daa3f08ca9e483ddb277751741a21f3399d6113fe811e310e547699662d2f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5882e86543174daefc1f347892ad556dc1d60eb9cdb21ec1b0bfa43111adeaa121bc6b31cb4e3afb9cdd077d0193569619774bfc50b12b603bc1723731df9d2c2afb2877d26824ea4756447096a6734e4fc62f8fad007832fb9397095397f26a9a859db056e0c4349b72e25e80e96d19;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h78187f54b562bac0ee14e55b332361fab385777e46b69c50a090a797f001ecd345916f065b9b74252b1837663dac521e4cf5dd25d107c3b16b3d15c2fcd1f45d2a9c3b496c3df07dfe850ba0b022e74628c18e35b744ef68e326f8dbe1d0f35513ab733e30d4cb868d8db1ddd7b2f11f5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8fe84a1cb2d66a5654e47eeeac14077ebc2121e04dc159748c97a063d91a98cbcd55c5c6a3b187c50601a29f7fb77a768a5e7308169a5a46a227a304557a1e87a3a8575f336e70bf72d6444f5fb71b56016873ead069b3d95f7da5b864f6a395729b3fd941d1d0756162062a2beb362b8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcba57e474b67fd73910516ced068f94ee9e72e3acf2be1b8b64e1a8e2239bfd57b66b55e642773a9feee15035c6e5e8186aa1a82bc5851c8063e4870d430b5a288126832d34665581541806021b0b6e703057a02dd084420fdeb98b73ce186b9784d05ac53cd184ec060eedc9d2ca3061;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf11caadb5c793888663df7ae9d834c982ed65bf7ad1a1652697092000f736277b915082dc80c9a02b7b5530bcc1f5090ff0968e5a7446a40c2ac79e56de32ff6756fd7e19a706601b20183766088f8d00c71fdd6acfd57f1afef99fbe97b2197caf9f1d58d81323f249be40d84f53cf68;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd5051a7072bcca3f7863b53ff7962e936407f0d40f2308afee5ad95a090a750f5e85e21739c351d2e30ce0c5d2cb2b2b15552ae939179d41129742f16db11b44294f0167922c31342e419e27b549a706d848c0d4811b73f5fd58a3ad773e5817e77ed47bf276cdaf8870603df4eda4ce;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbfbca31a9bd4cc3c7c2e60d2cf0a40cb5cc37fe5cbd8635f77ded049c13adb5c71f89a4121c3508d2ed838f0d2650172980706e660e4f34bdfd71985a5ec9cffcf5747ee11f8f28bed64c8b5df8bcc0e36ccbe5b5af774cbad71ff1d9bb1fab219dcaf6a0ba44f15e4ca276f29eebf480;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54101ebbc9ebc99b8bcbd710c83d2956cc9b4ca398f86a74bd07c9f886ec92f79cd44172cedc85bc8cb1d3ed5eff3f3e453e812337309cb45b711405373a622e83fb1cf64d34741a8568246196333ce865b6bebb023ea8521d601ec26e98d37d5c5dc976b94c21cca8862e830c8ed9aef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6c727f426979ace6c208530e2d35ccb59803a97873716136965742245f2c216a8dcba4363feffc0166b489bf7740f95b19e421b273d97ef4480d81dc8aa8df08157018a3bb4c596076157756f370269e312756ca954940f6b51684206d523117dc20e69d077d0b7dd19ca9a63b8b636a2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc804c1a7866bd8b0856daf62f7de127244d5c2c723de8961b3996849f33d3ca1fd34ca497999621571ad28026695776a6ebff74ccbd54ae54425d93c610f43f7006bc51337d9345c18e53a9f1f69abff8d5b4e143025aca98d770aedcd1a72c6f014addda0462e165739dd88d1cb97d5a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha9989d27f85698fabbedae012a23b01056ae32f6e2f435fa0ca77f7309a6549b18b447344fd82e80ff953bdd5630dccdd5fada79d2bf5f1365b15f41a58482686363c840b101898bc560905a5424070344ba4c2215608fb65c65efd4e017d2b40875133944e32e07db4dc857808100a81;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h12e3db39eb88fa34dcf5676689b5a530497c34baa205acbb9c2cba4952e9972b5eccecaac84f0fce9554d7dd1a9d311340849ce5730e03e75b8fee6d4e10aded59ffd0534b3f962ed3f8dfd3b168a39bf1d14d190b66c2c89ff0b96b162d3c0da865e644890b7edb9d0bde5ec4d614545;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44c95e5d5d5cb2336f188f41eb311f53a276fa4418983286a55683970a42a4abbe06fde5d052d09c55b03420b0d9daa1a076cf5f34c0ea5cba03d36ebf37889077150871306315feff269da73c0e692dd28a3a7461a056bab0284338794b096ca82c670cd9bb2c3d9e85f1662b23fe852;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h882eb923520d8fac5db11d89e77088009237ba0e48e0601838efcfc6d535e913b1ee99b807f0cd7ca72346272110c5409d5d83bc21dc97da647437846fc69bf160b8750ddd5f32a364d65e5713f9c68230b97969e871e838f88cfadb1cb04f2e66837e70b7b205614921439e4ad43d810;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda377f3af9f366e4c9a1febf764dc332ed3458dadd4c2897f22fb115bae14b47dd989992e3e7c14314a8147db6e5e15416ca08c60d895e2e9195e9aab76215cf3aae88c56b5f2281a78c8af133ba81032939772b2e898d33ee22d38fec29c4d868a29a744b3680fb47b251d20424f4127;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ede277f8aa6a98ed387b4436f6f8de3c0787d08544ef3f0c6c6e3b7045e57e11d9249a9cc09bf2a8aec9b004622de2c04bce0f8457a91c5b17d0d72d4533c079b875336f4b83c78f5799f826848bbd96723ef826e0816aba287e165b9995b1480d31e0c82aad3a7e2ee1bbd8b57876b6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf527cbf42a116661c1384547bf18823477cef47ba6a4bcde0d0218a5b7c9072ba090d81345b270a315c561a38f518cbedf0dee26b658a0a931d717daf0a4b181f174591326ca8627f3cfc605a9901d80504efe220a5665b1755f68854912c828fb88511771a62b4e8855f695de97f140c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3667cf1dd47febd6b1b2635b6c17a85f53c80bfdbbb6d204cf663fa9ef6b1ff34c726958fdb2f96c7a2720e2688dfbd6ac7c3dd7cef7dfd376992107218d46e21c0fc2ba375e31d7223a398e230f6ecdfe1909140c4e0258c599353fec510e2bd2a094b4672c35e13e5337c911b129d3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89e24a1163269ba75c01ecd25191883597c7380de963ca697ef4f30be23ed8b3d6bce12161b14bdb25f2e6195372b85bce029e8632c037f1b666373bfe9e4e49a1aa0ae6969092c71fb65b13d9c6528842e7199a122589c30528502faecd4741d97c77a26c8951e904c002dde61d6c11e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h812228c4af83613105c4f4ef79368ada3c749ba1d3b686b85ef48c465844736812f4b023bb4357460de88d1ffa0c62a7015a6f1b7195f140e25f2eb9e4d30d1d605bb741591418ed82010c4f8772bd4a86e85ee13f1568b10d1b084369507f924c2d4f123995a0fd51f69aad9e641e0c3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d9eadfdf68baed7e3544daa57b84507b28de61bd0ff1f1844c64ff299f4d531bbe8afd4666bf82d10e63d53bc2eb39c58ee035ddac978af922b6cba2d0c53c3e72892a96af38bcc862583e4deb32ffc1c50dee7e6178af578ba1467cdaa650a430bb4d3bd02349adb6f1cd9cd5514766;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb055f58672f50bdd5aa00b9569c50c39a85be59c6bac298baae60ad928f3df240ffbd4f807ad108894299a7f119bc833731fa70efc8c8cc9a0fde3101eb9ab2a9df3ebd2afe2720b7a298774fa94e6f42fc26a79b46632411f15139fbe0b767c458d62e3af1fa904ae199affb9176642;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he66511e87f8b9242de0a4db4e612af0fe15a1735b10521b7dc9963ccc5d680f9a4f42e8a14b3d059a0f170cd09cf7c9e4e15f593721cd7d73aac4bdd00058abdac553109761216654ef9bbf9b4a10e1fd7e5071475dfc0f22d0d793f8efd4d8388d082fb59de9ed7e7093b4a81ad75f16;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ab5e8515c296b46fff2ba9c9eccd2a4d85e3392b25be1fd15e7c796f09f225001ecfd6ac452e7c9ca80f82c47f488ec0ce5245505673bc4de8efee8f055a934105567c0980e16de89e67ff66615bd93231423812473cd873d803e3c94afc018b706c8e1ed38297262720229e57b0bb2d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h77ec1b580f4c5b4bb4e04667639b51e1ed549244a71dbdd42578bac9b1cf531bdd9fcca24ce67386ce17625efd082ea271661cc1791525b6317227f839bb69b2b460353641008fcd8bd363d4c04e3c8fcea3a944bbb8a78a60b429bdeb5f7cc6847cce6247a174a872523d57b21d967ae;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd543f7440b40840e87ffa50971e0110f595e9c72f48470c5a89ee054ddb29a08a3aad489c4443686a596888078341fe1e9cb5c69908af43e05037437c8b6675714f70fc955630a5bd8da11db482f8b6d3a46e74aad407155f24374ba69173ba79e4fc88fa85328f333671d7d90f3318ff;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e7bd1846324a4c61354cd680120882dd8f28793894219f751203d02142db0bec25d9a3e2a1d883d462419fdb30dbb4139df230eb22ea3e46c45b5c392f1640afedf998df2b7e60099169158be58752176a822edda2d6a530cd319030385181c33b224453000e307e68410c78e3b59513;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d0c6997f586f50198cee8c4f9b8436a8e77ed8e3affe3c0ed86eb436b055ccc6881bc7d34d436bf1e936164f4feca3eaad865afcd50d94e5081bce4804f55106e120107c8259ba192bbc404012d958547520bc2fcf1464d158bcc85196a83a8a9d38148d81cbae4caa00862c8ab2c2d7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdaa9dfbfbfbe9ef754fb39626909d94e60b7ea9c66d0faed7235e78541c5394163465868858dc975b762757ee49ddd7022c496ff58562d47fbd3ea93807260e72d3f2c94992669c7d3e1a1c5400093b63671ed07b6c3dd125710e3110bef7c2f2bc3d6e0a5d77c311ec2050c02707d422;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc49aaffeb768b8f2fbde485ffe6bcce5b433ee2ad7d22bc89b405a4b5ec8f179981805db104918ce57f5bfbb60b146ba0ed5687fa1d3b804518975d2d131482542893cb04b4d7864b39a693194aa736b31ec1ab3b1e6a256c9d8c36f9a0d8545a042623a665f98d2c409fcb95e8d26f7e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hee1fdbbd922c0329f00f1999e3a58bef669605852de469a4657726ed2b00c81e5aeb84553a785572846dda695d6ce36fbcbe31180968557766714e5472e532611a0b7be710362e5d16aec670c84c5489cbaa57a9dcbce11c9c4224b03315221237200a6f9c2954497394b4dbce8adf9d5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hffed8460e992b95ba23db5f45eaed5be8093d848ebcf1b156e4701905f0fecac3f4c58a46b55bf10e08a1cc639684c9ba7bc26810a089c375eae103d126f1929e1e49a4e3f091a0a540832410026265dcc9859d6ea7a1cba3118795569c1d2e24242aeef3209632eebc74229679f065d1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf1b0bf163225fec4bb1de61df1b2759801e46d389d8e21f6bce7436cd8ee3dcd4c79876b1aaf92bf5b613a7a8a444605f30ac2245dcb2dbc385b6bdc6e3a19f8f68444da476c36d0f1559a7047341673ef1546dc096089959bda8ab0cb5426f52e13a751e96e28584d93d44cebe35a307;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heb2c63926623e64de5867c41bbd856877503a47f38be0dff17d72ce6a2f9195b30814388afdc515bc31307e1ea3b837631c23f2f78237adabbdebaf46e35c27f49fd54b2ccf9996b239f8c210d8dd867294fbcb7c6978a9def511ace56f50df62e806acc37bf97bc7b57101502e52351;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hafb8a69473094d8d16309dd0b98e4af17700ef4444099cbe8b606b263274ccbdd7d9631a8de8aa4d72b3fab911f35ad62f8a3e27ba2f0c3822081f3cb78a9b767977740a9a50f63d14dca61ec833996a97a3fc61149ec0b6befad1c553165defcffd7b3b8f079758b970bb9d5418d5a7d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc36320bedc08c4d43946ae794cfb0a04e59a128657fb526fe052221d3668f74321daf6b3f386b1d11d6d550bd4ea39930f5890947aa908b7660d4029741432c3395806ed73a3046e49035cf2ccf51671d1a446e25ddc64a31fb7a39a8ed01823f7a95cd8335d6b290d0fe0f3424079254;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8c0cbbde0c41e80aee4a8cfa9e0d69cc26415f4c1dcb5ca63fa91c9e517a118be007343be074a2741677b17b1f77d4ef2293db8e4cd85008858a656c3e7312c3f811fd0dcbbe1844141c68ca19355c73e53794612b208d24c3123c73c8b4c593971d88f514e461911fb3edeec213fc22c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85af97dcce5790b71df3475d43d2af900ee962e8fa380e233aa1c3c6cc0367a279892f5d329294c793d1ad2d13479f87999549f444715fdeddf55e279c97d4d55618bc018bda49ed92d41bb15ed024c72727282c3f929d9192c09b5fc15d94e490cc86dbe8b13d31db77a39547ca3796f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4636feb84e2b2dbfe3f09036ebb79bec35ba989962ff48dec741cc4d3db1267f81f5f1508a8f629a1ebee8d500f4775826e1ea6fd21693cd3b16b8de61b19968cc6ca2326e5415583b60cd16fdbbb3f3eeb6ae63772ff3c4b62407e5b5ed2308dd6dc9eabc38e7ab262c220cb550f451;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb749eb6cd54c858ba5dcf5fc04ab350f03673238f6a9ddc657976876f37f2a56365f4e826c9daea7d3e24923e08b08a481cac2ee814ff62640013c60b4de3173c31700ef747bdcd312770eed9345d22c9327f55cf6a7762bc829f91bca1ca94a8aab2b5776f20a2c69325d4b0f78d94ea;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h375082d0fb5910b3f6b8cd04790b250af8b9fcd2f7d926f200a511427451c6f90180dbf3177f44e0b678385d2c08f71fb72edd99a60ff12ab4940e62196a3c80e1db9bc45050b1263e541d90a2ec12aeb29281e192f0a5283d65025f05aa73598d68895a052f379098189935e8a43be73;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae290f7a85a225b3cdf34b1b2a08dea6fe051d9bc1c5a47af3254f716c780e923753bb361927d4c90629223056bd4ead70aceeff5d3916eaab928d580034e44a70e690061038dcfa7c935e42f257060ced105e0af5a95e4ab76c99dd9a0fbd57461879e6da3d38cf0a06940500c814e05;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80bbd98626531d9d5dad91cbe3bd8ef78c6ce1ca942c41aea035311204f69a6cc6b296768f021c7de6239f78f84aa54a73758ef2cae94684c3d36c8d5218e34b70837206fc5f6efd1cab614ea5b8ebecd9672ffe90e0854f9ad8d393b3f09b1e8977fe7e8373c987595c5e6af0c68c2ad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc9e04f5b0e8c7e4286e878f7508233e262eee3e00c7a04e90b49ed463d7c8d73a3867774fca3e5bba55d7b3c835ad7ef096697455303d83491e391c7e913fe9a2a9a309573b6b35c068ade071d3e426189d76f72d21baaad88c125ea1b232946d893d660dea704616a81e31dff6c43d0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h733718d433781956149adfcc3001cb710bb59c42cbd16e1165fd45eac125158022bc8dc0884b125753af5bb537ba71472e2ee9ede1447132448eff00fee0d4d16795c76d4a41fcbe2ac8eb9c15e71f4d064b2f08f640c3a8beda946ad6371b2e22d4dcb8035ebf4740aa7af0af046783b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcc1cd31194d454c7aac703add8526e7a4e800334adcaf370e9f1da24e67b17abac4755561e85a3ac5525a0dc250146f97c15cdd6c9cc4aed6cfd6be169a15762f78650b6e4c33cfbbff3cabcf7bac0ca9f39de637378121b4a326a26f6c5a8be0639b98e1b9864f60a6f95e7e7d31eb50;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd272f8fe2f9680fc976231c1822f0c8dd62f60b75209fa846f5b8bcc9934dcc0c596a5f6474a65dfe5069f4b0c83ccf3eacba5be10f8f1526f47d845cb281dad9e8b834458f6bd4ce49052240ca77a8551349e9c99f66b019766851ada96b697130b12f2c98543514dcda8d46a54513ac;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd230d990a41c70fa1f8f5b1765e0d28940be011d26550a1e1a84c4386140cd157f5200b2d912caa9380b28fc4ba71da6889446873caf320fe31b9cbd983f5af2ebb93bc08c5e4d2375c6bfb01c26f2ee6f4efaf9d9b1f359e1801f04626f31cfe4d659f271a4677ed908f600a0ce42d91;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1c2b93b121de9c7174859b43aebd8876af6a9aeae96682f5fde2daa9ba10c9b61415d97db5c99148dc48ec1cdd9a2d276d0fa4d66acc4755da6067fe8c3d37e759569de3cd649e1955c34752526f1e421abc5c613039cf99f0726fafbb6c91f544c5a1966e91583e11e80b7dfaf5f6776;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h10f5ffe9ac6f660301cd1467897b9a30aa9842df3cd47278c27e820a0a4ebeeb65ff6432898d9f7206d17467d684e6b0b0c83cef53358d4330358d49ba5043c9fe093353055d650a0fd821078cdc7b326f5587856405717596ea01f3e625d4e48f3cc4c6fcd963a6d2430baf8316ab20e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9374886f43f89c7999508bf0586ac6c105b9bdebf6e41a7c53c4f6ccf0297366dc00c272df4aee84f3f7d3335257196f0270b28f0e11d9777fe79e092549fcfa0de504654c493c8a61daa27e8b9b265a282af7c13ce5c0994853552839badf415dd641898b3d50df10634046a5f7a1075;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he76b4be025ffb11d0c25b99ddcf4ea7534fe2b8c2ffa7c2438e44f51521ea3565c61f6793b609926b33bfe4a7d543f15d30d04d81f7e1017443f4da1c50fb5e65fc79a2fbbeeea97089b794fd358a37ef16b6d946c8ff4e68d9d2be77333951ce42f6b7ccae6b015196264a88d0548fe4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ced2eb412b6d98159d531e9ae2b8e7107bbe5f48d24deadf0cf930fd0f1b8912c6d95667c597a2e3810319955fa5203185370ec58ec6a8e213c87647d584d92f5b6c24cadd3084bca641761a75a609998c97d5fa28972fde0f8a25c0234861dfd05632ab457319f3b667f6aa4ab92fd4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h687defad155980ad3c91fb8408e053d43914e729c19ced073e0aeed9b11d7e41944cb4fab8a1a66fa7a68bad08f2c4bebfee84a75071e49a776362e106ec4f210ec263b1b2394e4b98a616db378a71a4d83788afb3e7d0103f10fa20606cab5cbffae5a1da5fb525cac78a9e08bc6943e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha95af7d926bdb917ad142598e3dd829993da1a34f9ae538e90b143f11e9221df59591b76bfe15968499a923983f02e97f4d0c4f5ba30b07aa17b5f638f5956c773f9ec0267a84c7dca65f4f500eb33d0433ca334c8e284e968e260a109f4401c371469182ed33bf2f2cdabd78a30a0245;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8aa671853c84539bf78ab9c070aa8722f560c318eac04a444aa2dddc56541349500c7555a6803a9f4b1f4d183b5b0f638d27a77edfdfc9e4c07f0def310fa92a6253225cf66f3372419dbf85ab33eff755a965088e432b548089ed8cad87b92a6e4df9346b43a02b3bdea4111c338451b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h84839149c0be69df760e0295e48ecfda23ead6064ffc9b750e5e281adee70de5d3e81b32ec453ee197c222a3555e68124a1e5a4ad9f928ced641e4f8e1a3ad8aeb7a5ef08d9637322d5765b90ab5e22bef743a37ca6a7633e61dec0fd36699d41ccd78fa2a9b6fe98a85e3a872029d65b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h373a310d57a0d80fdd64637918a2da9efe50b5962e68ab220c0a6710322709a37cdaa7978ba9f4cc88ff70fd7f5768219da294aad5392c2cef783c152d18ed157a834fc1cb25fe0cb3be34842a52962c781a2162885ff3e1ebb634c38150fc9a477d4e698c014b544cc93163aa8856d36;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f46bffd0e6765626eaa21661bdd625485e7d04e820018ddc8bb506347509fa2d1b39f60742ce025603d65a2931e5c102f5d093fa81b565320d559d8bb9752f467cf3c570debe7b8b0e1dad8576c5f483872b721af11cd8a364a6dec25af577a10f1145fabf5a10f7bdd1591f21b42bef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h966b1c5261cc83ae9ea8e3dce5ae4e2f564bbee9ed688a86b769b17c061075600f9a61d47669407893e3776b090d3a2baa26ff733343059fe70674e258954e598a42c05f839277aa8860216520ee9d64cb87e8702734cd612f1198d7e6dbfa03895f37b571fccc5bce2ca067637573406;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6e5b4019c5281dcb0f80e53f65eb8dc6df9e04ffa814729a2059b5d1196e0722aee113aaa0d1645886b11ba20d712dae94d428e297604f6ac1b616ac0f20f7692c96fbe59b8d2cfb448aa052617fe2794c9749a2db9284a65588669023d24a169b8d8041e0186c98f548dee71a622015;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc48a1b943801ec501ba5e1f6d3cc6e3adc0e0caf58a3d37ea322727334222c3ce86a80776764595363f761878f0b243243f5908689ba10b62b364d91b88353f535663d605e7baff05394d9bee5e8f73340e4a859b1b1bb2b494fbabe62db9b5212bc44ea592ffc3b4aee232954a152e6b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45bf567224a548f6b48f7e70699a81663d5e3df0b8ba58988a1827b9594630e381acffa3296b7e7eb38dd9d016ef3d95064095ea88416d1a8bdd2cefe5030d4b024aa8a43ea08b5bc251363b98b0d902c4b28fa3ec73d8902ab3b4a1a2d8032e7b855a86dfa070dd01ad47ddf32ebfa8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd59761310cfa45b808b9b0ae15c968c159bad48b08d75147c805df86588970903a664d1260bb17a7d43ca8860f663888c2f9b1d3a90239eeb5ba59a671698ec9ad911d89d3aa21467b0226c9d4f0eb64dc6c00bc5bb160e7c6141fbefa3b6eb39c43c129a5f62d679a11ce45176351e1e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5606dc389be343fb7e4774d1a3142ac3160f878e9c3b1742f2c379dfb6cb36f44fa5bf155c0e5c24fe43d6e3e064f826ad09b43ee8d08de353db983e6076fa127ab9b834910050eb9b2c1fd407876fdc46b8473e900f9cfacb043ba7fafe14c60a6c3c575a8b857787b6a8143c98cbbb1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7c4309f309729688ce347b1d7ea2f0c16fd0d92a3d7597d8c42801b099ef1d87bb3c3dbfd05d87b3426e33202567db3b28568a60c792d2fe32a6f34da6e9538e804214b8058610c80af42a41d1eb4ad4a3415d0193898aab691fd302e4fb2f124d8343dba93fac2971beb4b519f68368c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56cd89d8623cc246287a2bbdc1daafbc59000cc43abd4c6850a0959f4a0a075ed47241375b1424bef63d1f45e1b13a98c1f0c00ad295e29804913e54714013477cba5bee3ece010fbdd4eb4b2442d7b8a2ca1d4f678765ae36d21c625dc81a5c0b70df9fe13eae8b9a266e5c362b0a66a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he5d5cdb68528da8e4959e05b5b1c2fa28af03a5b76b154e2a63ca586c49feeb1b45a341d85088096a6a641303458144cbc43b3ff48ec53f57a0435e993ee3a3b368bd03b20b59945c7b4316aa135d9e7fc33537951b511fed1773edfb7ccbeb00edb8590c0508fd2330a5b8093d6f3c96;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f578b7fe25703f9dd9399b38761d46c95da00b7eb2ce78df6a019bc44094133756645cdde677fd8d8797103c0f1de98ceb5cb2ea9107b525dd5225265203fcdffd1ab8e61274ab74393d34e409c7efe03d0d5b6caf98a46f15f1f888de3a21f984ec2b3411095786b5a920b166334609;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he2c088656123d530570a059f3350872a2b400fdff77512ef522956d43ef36316c5dff4c0960fc6e251cdcd9ccdd4abf642936a81d2c1c034fac12a9c1401eb38389b482a2b8c7f6db05368e5588ad67c90bd805027d44bd5619f88053105a0a4ad7893dad643b9a5e1f39778223f80158;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4937c138cc5d782b40442a8146310b0b5416fe43cbd4f7d2ecf7c37c1b8845d79860bf24c81904add482120862824476eee5b91817705a9c7667a3053fd32a1a45aa193c5677436087332b14f8723a67e295da6d3af127d3b37f98d410e13cdde48aafdc4854b2e90da58e447639f3d8d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb3464fccd50978b67238d628c84d6d6c57224b06712fe17e5b0da6430e7f6378ae5f7dc5bc566b962d02cfd35a25ce2a7f993d363990ae76439ca4b7cd24043b2ccfd363d22379234f1ddd9d3d1d313dd705d4981b7fa2d45e779f059dbf553bb26749f826d516cd898f0cb0917a49cf5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf2317985d8d05854d0575fdd767526464e104add559652472d3e6eb42aafddde261924b1ca1f900e8b6e67cf7e9362dc5f0a4433e16d462117faac2ca1e1ee9b336b0a30807c9cca163c6c5f800dec61cc63fb92b8d91f9e564c770082ef0cbbc346b677b62f4c1832da9c1f3dbff6acb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h30bf9f88c32d38b08da7ad7cbb1c45788281537c0ed7c4b678a6f1f09b3defdc255ed3eedceb6c3cb1ef668eb3096eedc52d3b45c3535269f804137f820eab3e762655d785af0138389ab3365eee88d3732bf9c91acfc6781b037e069290ca7f522ed3d62642d5ef729047bf3c3c2aa9e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfa2c1e06ef77faa969e02d1aaf7658436b8ef2cc3bf6468c313ba93ce5e728cb99edbcafb6801a9698e4c2b12d2b2ab6960de5fcb45fea4e17fe29b750c80694e781aab921f7a48cc8591411d01e8301d869141c0456f4c51dd216cdc266fcc909d97eef5a1722d37b845aad30469bcf9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8eb6ece147f75dd36cd4015c89f23e449f8c48e14503476ae6ac99c8366265487b3f107b8c251b36f4b57112281e586a2f83c1adb3076d4b4952a45eda33856b3c09ec7b92c0cebe42a91441fd68ac458a83ebcb8fb010d5101be246377f274dd9dec33a21d9ca65f4f305c6e630663c6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6700e5d37e860ed3bbe7e361ca22d46f36b27902994fb4dd13678c40efde245ceed47a75ae72559eaa753bd9895aa438c0260047c07fa442795ea1cd5077256740f692609983f3aa876c876f127b4b6186bbbde7b2cfd0bf26073a717ef378f78af028784188ee6b1704afebcdf9a459c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc13e362d918a06527a9b285ec7a6b88411bdf46a97f5cd165440faac098f8c92d9b9a4d5fe17dc981ab784b95f9e5add9dd8c1d1bf83fbd3fa512b59c849ab003a7e70e67e3832831eddf5a4de921a6ba10618be960ea87f5db8b8a30b9a8dcbd2c3bcf9386fb39a7f2ead95ad20113ad;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4074c1740aff2a97f8fcf561348824a5b786268e0b3c6602fb96319b837b28d1d15a5790eaeefeacf068e909854a58a85922901f278ac4dc5b7f170db39932567c7de7e26f4587106dbceb09dddef1471d4ab89e5bd1454f025f0d9bcc94e801ce470d72c00f27abf828a31deab12b232;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a02bd279936ef6f8e694bde112726e1e82854ddbc47c46864b552abc289bb81e59746391a63656323b75116e6ff8664e69bd15a864c868762d271d54f8f03f2e35281a602f093fcc013abbc7d733c784fb550c82eae88c0f8ea765d5959e89aa69767cdc331535cbd1be59bd03213f9a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hec6069da46b2c147c91d4eb57d13d73dbba2e2a98d51373038925b63c5619e1d3184b932061934bf33b8e9dce30f387a67e0b55e81dcc17fc5a2a94be3d9a8151c45e05535ee7a5288ab1886536998a27cfa5890cf1a3159b5cd05b59cdbf1b128bd1921ef2d87375f166b33003187b41;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c86619540ff3848289350df3aa95256445533dcd784c4e6e34631d47d596bb1369aade98c96d187c78cec22caf811c93138aa04d7ebc73d51f0555e9eae622c2c0def516f79197234a344a8728bd4dc2fcaaa9ed23589247d1a07dec70535cd5b76cfb2cc17f18643fea10f48c6ce695;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h705b904d2f19561e41fbe7cd35dfdfc10ecaca2ad23a746e503b9a93759a57f29fbe03ad6ff85a72fb164f151acc17708a76ffa4b63573cc4dcc66fd9b5ab5e74508dafd1398ec89258c1383f7ab9dde4119d3659becc5155b567d2df44a0a124f9e6278ec25d97d56289cbedc2bbd4ab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he497f3651d2f5189f6082c5e0498ccedcb083b9909dc83c93561e7c5a20f9f9d9bfef69c131757c5f75a34fd2b751ddd2a5f98aa012c937bae36728401efc0ed67e11f216f97c21da9e48f2f5c9121df01ccd898e8905ed7fdca0cff71d25513294acc78fc91aef5b0a726e6297a322f2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71a47f3ddd0d30c838998c3b096851c8c3d7b1b0e6df09a1d734cecfbbee89d41f05c4e43e1ed73e504e278d6d89d2c66253c1316cc738ce5decac837e42dc97a1d4b6e04f576c29eedf902d411afc17e52497d21b78fe6c91214e8790fd8079a718d82083b9a8ad00a2125e4e05493c1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f2c75c083a9080c7504b1c54306eddc074a719967bd8bc0e646fd8e777520b2291d2c6e3881a107f565c3d1fc4a47f9a89d918b088216bfd5c9cb8ef416cec1f0b0fd5b001895f8aad7253abbd746e9a2bb010a5893ac4cc36b1d291dee2d05f84f84aea8e5bf4fd9bf2507c0c956aca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49824c31c7683a4041d2e97d7fa18608420bb1be2cce953a2f87f543332781b698bef20af688483f119640e1d626e29db3dc3b54340c277d8287452bd93f1f50917b778f6130f2c9b0b5b6954b544108e63c288ef9b60c67a662a5cff29a13c386567e3209d5c4dc6f048cf9b108adae5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haa6c2012fa78cc4a415428d044da72d25e117a35e05538ba728279217e0309da665c2d864827d8242ee6a6e73e11d9a29dcdcdf6706e251218fa91063cf3d4892f180a74a46822fd955acf97572313238a41868581ff5b3f0bc85da2ac56d7c39dc8d2e3e6762a35b175ef029b0d40e2c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdce2c08b7e8df2a5d58d00d48003f7994993fd17a6c84207463a04341c0484d2eb9038a73345d8a08ed8503aa70c54640242179bbcaec0dd8323d1a63ea52d6c0e82ce6f14865868b79c08cf8063460463d963f9d1d41059a4123bd83b6bb3c6bbbe9493a2e1c8c48b52cf0914b1c183b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hda886a95f9cab56063902f0af6284fb64262af430ce2efde488dfdbeeec6064fe0834e088628f9d3bbf1e5356c968898b2dad9ff5dddaafe9da04aceb6a2067e8913168e1e82a37fbc32eaefa3f097e503559427e013be5faabdf3449aeec8d380d5b1221acdd5f7c5ce901b476e8d315;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd0571ae322f4d22966907faa870e990272a96f35fad8d9c294fd87a9f368b418bc43a8ad918b9d58bd76d05485f7357a056b65b8cefcbfcd89292e8231c1f4726910515bbe601d276a82e9b9b72af8e22929ddf8d89227e4d46b2844c7d4f7a58370a3f574e61107ef11d373b6c7111cc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4dfe34906971df3511601dc644beebb5355bd555c9e1d333b49a1fe1f580822e01812df61aa8ba5af28f463d27c8ea12761f46b48b54c128cdc9fdc316f66063f23e0e9e4616e7b7fc5526884375b50dcd774f1f0712a95ec88edfe9d495652be7094985955dbb27abcb15eaed23454f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb969246d5b90160586e501825d9b1885dcc1c610c2a457753db7a3af99e9778c2608769997b7f4f66f8165b971b1a8a52997eb14d020decdc777af5e6f4688d1e12a1ff92e5a4d08c78b14b0f1336dd5fb8b512766fb2e8db274d6e8f31ddae6d96853acc8617f57f2d720636823b3b2d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2d7786c5d5761ec3fa9f0ba6a3c35340da73ffac07d019bf85fb0465d25e830d0a26c30644378eb03477bd0d1f4fc898a8fc2ac64d1c3ba7357590bb28c15e29e3bc70897c4ac0bad7f6a778fa0716ded8204c5a211f20ad6d6a79ffaefe71cfca17bdd1063b6ef485f2ac228453c4579;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d2c184d378ef8fc41d2e1b15e6f4e6f865725007b24bed184e4b595b8e7271e88dc41f288731b39014f09d9b62562ea8ef7e08e4c97c952b8e5d4737803d67966da39ecbcab96d0c79c832925069f176e68d925d5d1ce98e4fd39d45bb9eef3f520099403c7fca7859796090d86bf32d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7aa5f9bedf4555f6ab3dbb297be702ea3e3dbcecdc35d2e9cafc6962b1a9535f62a0ecd9487e78105fb91d895a30917c38431200b0551bc883d310a500fdcbdd614b0bbd8088fe30ab35c4285a61d4020c7773ce63697eed263ba1fe55d881f36105658c86b9cc84a2fe3d078eab8a6c5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h80520080e6456925489605961332a0cc1fca9ef4a25131173399309fd018b4482f9f4e079007c68165e7d36e85226d9b3937dd44e431fa45116485ae139f14e7507afd9c23ac8f056be5695560fc4e003ac293d9bfd7b58aaa041efcbac7bec5d27e451ce76f74f7b936c2e5de8bd5a2d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8677f3242eb8144ddfc3d4c784cfb9a3ff7efa7ab8314a21b49d5cace2c15a3cbd0ed20ee2fbf9b3dc74e3f65526b23c48cff9e9566bf6c66b7d87ac4301ae01dad0b5cdf51612e2bbb6b3efc17f68b3d3b3d8a894e46be7b89c9200fafd45d99b059c089782f5a5de0fd13f4f739849;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac3f4f9ecb93c9f12782d13c2094d121ff8ab6755a90cd10fdcf3cb0c8ed6673a51fb4188b5a6eb1afdc9eacd5cd36cf535d1b3cdf6cdaa0025c05b45cfb8c21c306c45d7dc9891bed5087b5264e3f2077ec535542519111bbbed47a2d56bb8782b671f80b80e64f041a7107034d3fa2f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h89d10a6f7626682b17551c78e4d625026b39c6c674a7019bc1b04119162107da3e0c576026d3f13454e0ce406d7bdd5b421ff3c536c70e947e0f0d0afbbaa63c684f1c57b7b3def68e421bd3c13085bd756111aa2498c45563b14599d580e3cf8fbfe401b6061d846204314fc833ac9f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf72555313356c0d9c8e0067114062d8785c12e8c0b9abf1fbc9b3b6351b5b5c3cf1e251b6161ce97958534de29f782e2bf294dea516fd161f0701d13787f31104b38be6bbc27b912518d0e9cdc33dc6f1b296b515ecccffdc0b1f133f549d5f27b060de8d9e3396e0499cbd24ce119477;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6270f957430bb8317fe555b66b054002e18682862c1cc34fe014d6c944bd72c47d44fb611125fa1fb0b42d994e02e430659baace723e30ff41e9453528b564de1a3b4bef3486cbee68f9622e66c212f17267d5f9b06001f5d0cbd24fb8051a5b5a09c46e7fb69b2fc519e2018fad8b3ae;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d20edc71306ec420ac4842343f6b15a19c11e7716954f02d2cbf9848b617d36bbc66483aa4df68c40f388215d77a2ff1b8769feb511ed5e2afc1a8e03732b5a26064f1327f2a398c962354c6133765afc1c88c42409f79e776c4c302206bb9d9e56154dce47411f1e130ae9234916ebe;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9b34e7d3996c60ffa830a5c63c24c0da7b6247609c7260030b329522852efde4b6607326c11388767d983ccaeae7b1fc0756161f17dbdd9ec3a0d47065a474f9620e3d4c9c57d24877f5c5bd9fa1daad58618a18ecfd8bbec1e6073585fcc2b444a0aaed62e4dc23c0d4ab69f7ec05d78;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e3c075a6c42970f3cbd6b3e024b7b6fcfa0951c1f903e8aff71c889c2cf1416c6205abeff3b138766a70a1f73dc7886e9428a98461c6bed94b14809eaf0add50f41c9ef05975ab67d2c492db60025b7d0f7132f8cb5b8698954b4bffbe645d2fd02b8b3cea6d5a7d758332d14f810f26;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4bf8140367931250098d1acf8d4b8c30eccddb02f7c22af93cb11347c115369eefe9744842e4b39832b5256ff0a8fda67c2c2878d0450f7ca51cc7c91c568b329a54d3494abcc097d3dcee57c59ee0ffcf5266f521db7ee1794fead1449ee6628240455acf1fafb824665afa7f8078828;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hce816fc6c0681a62f7f29449cf7dba3b74684b36fdde6f7d33b4c7ce03feca43b93aa5de8ea49af36b9f006ae4e13cd4caace4bb3c48d7066fb18a8c1b21ae66b28bf27ee8ac8caf21635ba678091408ee3ed905cc593f079c379723d5d6a43ab689fa9fd2c04aa9e7a06a59da2969fd1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ab90843527f37274de851ba99a9e13150c263dfe574f092faf8f8d9a1b91c32bc42b199bad7bfecf6a01d5959f4fb5c10e3fb87a118ab0c21ac59bcda40e8fdf0f2e86be54411b0ffb9761c7f96278cc8edbd169e732444cb7a296ecb632443adf9c91095803b58261d2c798bb28afa7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde2f872e1272fa9ee12d227546746d7bbd06dd5eba909ed7351666a742dc7eb560811ac922a2461d56f374558b0ac8e8eeaf7355159e35444ab517845c1a2a792392bfe608288b7bacc9996079e8509d148dff5529cf71e48c49d4b82e8c9380bf192f30ba5f02df5f0e43f6bf643ac5d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h886d4bd91876fde33700b602991f86b4af222c7e81a2bbd43ebf45bdc5b7e3934a713b7a038ca113883b15f401dac3386ee4d56a2714120076075574d50bca35d5d5ed55c0c59833c94352ad36b655d8b3938b54c9492d97b68a329089877dee76fc00941c5663affca769777e1a2109a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfae19996994507e3e4d8e24a1469a94418dfa9a0631e9bad6e7bd66fc0d12d488c22b5884a1bf2aee72b7978ed83ca508d70e7d995c753ac34a37710b81f3d0d55df973bad7006d4b28bc611d525f1ced2b8e98e33ca614143f07bf26ddaf61ff7d8f197aec79447f16a76ab98614d61a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9317f1c3f1c1c1b5f13e59f8549e64e3f9ad2fc9856b89c50ab2747776aaeda8c509881b3c1a5c10301076b6c0091f8324419806c6e629de3c3306f46c9ea3813d5b1e1c6ff3b1dd810ca749f65d58111597c0175f6f8dee3b34a0203f7a4e4d4da4c8f2d0e4b714e85cc382d79aa5c93;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2deb52d83224aa3899f3dc4b8ef1e60abda5bc0f705cf89fe80af517b6e18953fe3fe52630bccac40e053549b2a343b1626cd6618619af27ca26a13deddc8d813b0029aca279e569d0ae24c15689372806940a2fde4a09a39f9e7775005c5eedbd6b73bcaa9a72623ce53cb7789635653;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85198ec1021db413b5b42e8b73e8c612146ec144590b9e692e514bf2f5bbc3bd6ae1d6e1a32f7723a2b3cafecdd511cb6de90c2fe41aafef6ae6d8f7c92eb29ef73a728c7544ddf30a8492c4bc93750ade9d36538fdbbae1e4db1edada9110612599f8780040283cbd9b2ff2dd186afcb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he22d533a9bd08e7f113a26d8ece188a6e18a08507a673130a5355a30ed304cfa12c0d3ab959c9ca643473a35776081b782405ee8fff57eaff99a464c408a2d4f62b6081943fd3eacdfa7b81ee7a3c8e6ab1bdd029c425e6945baefe71fae5b8cc234ab797b52de05d0344ee20103dd1eb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8afff0ef5e85a4b2a1fc1ec95829b436a15b48f3e3ad7ab8c5104b133562a36bfd0baaa588cef5e2ddfdcf67e5dc00285dd3c443a2c905d90cbeb8f53a409ca8c95537b4fa53ae67b4affbb6e5da1182d863418ae24983a561f56c0e9b90eedff31151a59256a0368e5e99a14f3901b46;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd2bfa3184bf71eb43efd447533ece46ea1b5b7f3235516055604748eced6813d45170fa18233ad938933b79c6be58f2d38fc3a793f48c04ed2e966ccd87141d3f8e1ae2b1526d9869fcb386ac5f526150ccff98e2aaf41b86aaf079f730dd5b65bba8bad3074a75985ec7ee465b65e9e4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf7ecfaee3a3d944e4ac419072f813d54b3dce167b5842a736e8dafb6ca857a5ef257123727f0a349353170a15f56bc24b625411df51423eda04e68041aaccf7d33b28f48cf653ffd02315830ed3e2b134f9f21a15cc05436926b55dbcef100483ae07c8e08e682fe02c3b7adc07e18ea5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h875b313f2ccad9953296b0b704afa7d3480f277e634a0a9cb52132b35cff0b33947ad3d494a52be6dac5609efc5d52d48a55017b15940f694e6e1f8977c42695c8c2f9dc8e0a4656cf9fc256502758e09d310e917fca74804df945c926b7bf2f6b020c4a379a132a61e35d94d3ba51efa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8865e1fd88caf19b9b67085a3cf242e491874d34d9a2943817eb751c069a7527c6824320b382bdab2b7735eaa0d0884f210c9acdc7f47bd7ab71d668e6f62d0b1299cdfaf171cc2e9fea0a57644f5a1a75b9b4c2be1f6c37ff6f40268fd97c3a481e42d3c4ad83ba10c282af1a7f72f45;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he32ad155622fbb1d7b7e5897aeaee33bf600bd3c28af5fe93ea16471d971bda66b770250ceb0ef88f531fb9cf1f0a62617c3d084ed8d4fbe23370027bb7a81872d3d2160b15919953d7780995d431fe09ff5f53a920c693b6bad62f028dfaf32781da7e4c97903fc18d8126592f5a7294;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf30231cc1435a1b95c074000aae32b90df5f33232d45a00971d9288ba50a9bd0f5b3080a5e3493979e9d09be41a22f2041272ce6049b5ea00c2754ad5cb9ec85faabf646ab4e4b931de82ce74a40c21c01a9736631f797511b2e501a3b8c6967b8ec601651fea8ff217b318318795a250;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had105f6ba1388a18d28746398b5c4f949afc68f1c4c2e3ae6f7be18fd918dffdf3259266a2e2b49819c8ee400877bf23de70d90f88a2e36aabf0fa804805679d7fbc9935e049b9eb93aa14eb8b6da5c372dcc8efee5d29be27a0e93f283a8a85abb4de41a1009f6bdd4fa4660c5026ac0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h75496b12c4cf8e549ab7b4ab22b2bbcad935efb9831dd07e4690f78daf3b7069eac64484d4b101fa8bebac8382be708ad0ef58039a5577a0931dd68133f410520821df6d5af90f8485239c011f8c4092f16873e24ac5d7a6ca75bdbdf9ff58179ad04f7196a430d5c65f272c4927fdec3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2a90439fec4ad3e9f7932a420732c02eb5527526e50414faee13501865e03907c82d89264229d6036ae0782542936764e8cfc63c4921542fc9723f1e019a2e72f0df53f02ec139da2112f8e04291b78aaf7d17d80ddc65d55048408e252fe87604b0b8a0668edeaaf6ef30d83c6e10658;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha45b9a52e5c38da08e34b7b8b26a780c635e27d6a3166e346cdbbfe5685adc0507b6fec08a0963a72967277bc2f657fd8ee11995a0e57a55d7d0c6c083f727a5abc47f7627ca0b0134dcafa5122cefb0ad3f96ce424a371b336be616103951dbafba21e660b0b5c10ba215fbb3a024839;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he4b8a9988bc9d5c016cf5a2c496f540d46f3d336abdb1302dcb49cdd15e5985ae137dd3b99ef336f3c706c3af5c5f77600a57beb9af700c6c79303d76c0db710af2cdc0253c9e56011629fd4a2d498260152af6871a358a0fe2f56acf67e6e2b24001a5486ffef642462b2f4740d2ce5a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a80e94ba6b3e52665eaee4992c77b0cff81cce2b259eb72c4b08641b045515249513ca469ef3d293d7aa8d6c51ed890e2e0390c8d46611dad97c40af2c075ac1031ccdfacfd2749448e49dd6f1da77c78f420b4d6a8122950539635a0508220793bebaeaa5e8dc7181f7cc5b85e36c15;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd77a8c16cc03e89ea7d6c4df21d9171884914fc85a69a92f6be362be5406a6a3a475641e7814eeceeea5bc3ae8f5ebc14c51509a2c315e29346ca54e6d27a9d78dc73a7057615b7de488cda4a9d6a18039c4883a57697c98d70868128babb2c8d2989866055a22083135f05c87166ebf0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3fbe2d783705f74750859cacf770d7e11ba61c9f10b59471c8bfa9909d600842b61d6a4ea5f4cad177a7d2d5b27e7133cfe112015ec6d11f1a0da15cc40115d149751dbb0c54306d115f3413025f62fbbe5aa164e757f8c42a3c8e3a280340d646749197fc11fd94eb379612fa6cafdb4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8ce6509e68ed349ea7965c8250d75794e7236f01e0a29a0649bcc258e6f5180727374e6e60a9da6348255257bdcf363d4d635ed4cdf042ee8dd15ac0c602613c837d7cb7dcd5b14b946bd3300d2690b55d12d8597df490ec5fbcafffdc53144f838dd9c6666ccfac18f2715d3fade065c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9049349f188a504e0191290c7000a907ed9c0c5f24b260a5a62b62220bf12807ffc6ff2cf2bf4e14f093ad67d371252fa4bcfb22b624c1bcc04cde4080caf547a0a0aef5c2d019e188cb9315ed5c4fb795758c5299837dbeb97d837acc9e51cfeab341cb1e75d37dd33de32e1aac706e2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h681618dd1ad56930052023a1a900f6f48a56ae816c15b2d38e413fc4bdd3e18087fadbb0ac69d93c2224497aba36168b4898b56a53591d1cc881cef2e70bde1e05206faff2938356104e196ecdd4de7e7167b4bef04decbe2961a180d629d35ef725c53e8a4f2ce46d5ea9b43591fa5e7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h809cbb1b312f6a8e8f4e7888a9e25544fe17474c5fa23fd1b87da0ef427704b221a0f4fbb1b2b070a3a05b977782ede608fd200da76ef3841b1a8b6100fe7fee43eedd531d22f30863b6cdc4b97f9f05daccc2874ab8250c020f34ee2a9ac0429d52ddb55726d188501b9decb08b5543d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd9ac7c09257f74ddd52561ff7d94b42891771f6a41277050eef8ed903887bdc55d188600c3f992683d9ecea4be04e88bf016e65c585764e05885f5a884b874340099b20091aa8541cd395291e4a61dc03d763594b8f2bf97af1d5dfc941d8a337e4c2685e34d82fb5864468c48d01e19;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0f009fa8d74c26c9633dca6bdf207a0110a49ce3d9c271e3954b3ae6d38596c6eb1b3f41b1562ded8c9026eba5a9a25734e091c19b8a931f1a7ec4f6e1f33c4ac960ed1c8d330768d8166ac0b60675f66239497036d6cdc3596d93c85cc0b815e1407a73a72b3c310d8197718e234338;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h33bf48a0f956b1f9b930fb712310b1f11da19603d0f521ea0e5befdf111d483fe513d9df52f34f14e276c96f70afacc2deea311085ee8009a668229a30737dacf6e49a01f48afa42e63e9fd461febf6fbc60ab274495f89fa6bdbcb75cca5e9d71b871a0c385f9c53e310ed9c3a8dab21;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d4899586fe69dc7d7952021651355d24d7fdfa58fb60c6470f61ed2c5a30188dd36119cabab987a1dcd23513a2ba50362597c4c455e62fbdb0a1c3911d0a963252ba7359d5e3f1079224716e8acfdc25cd9908fac331ce62baa36e5fee46843da6bdabab53443e7ad46796acb0b4955e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h714026c5f20d708d45633519053916541d184e3fe8f65cdabebb5c9ff22730adfd8036939c34168bb260988a42bd7a34f5333bc462ba1b1adb34a69e0d2bcd0118eca19bc8eca97ddc9c76a1e2728f36bef217b094fe1b189d8ec89eb43f5576fa53a748c660835f2c58b6cd330ebcb2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d8b70c1fda385c73af87efc69569503cfd7eff2711cb06381ca1aad00584a9c057f7f5364157cf0e57e3202eb0f6c54460ea3a6d7cb196735bec00309e49ed5be9b3260ee9cb0b5d733e93a63ec352f82ce6a7bcff405220e053c90473da047d431b775fe93fbd4c8c606d52278e8f6a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdd966ee1f48a34755783239de9ee43489500269e2a5214345384aa3f5c7a1986d16dcd99efaba69da88df236ed9b381ae746692dc9e106a2e0ad0abec7e5326cf7fa07896a3f9f2d41ab28955a690bfdaa9c2a35b2469443eaf75631d87662fd680440d842a972ab6a07abd1987cb7f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he489014d4c38f54cfe4c4820825a5c61530b070066286825fbd160a95b69b9eb1fee1ab7c425be615ff023560faf5b10fc0a5d0b786e5ed1877db3a6cff1cc0f5b3abee9aaa0b90bf5322dc4dc7b57406bf15917b9cd126a553ec6b39becbfab5a7f5602223ead0da827b757897bf1e70;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2b9f85b055ab1a195018403a9244352c670d6757f01cb4025337e826d1379c94d502dfc0c59c72205caeea8d9cb0cb24ef4ef36bf864946cc5cfb3c35c6286f4403e1ce438ab7ac5cc70a162cedaa03d642cf24caae951b53df36ef4d522a7cb8437dcbe099516efadd514446f81cf3ae;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d6838754318fda52f437e9dfaaddcf123b76a9dde1e4b157199189dd2eb54a0a0f424e32250da2e348556b772784f0994ec58dc4cc14ab0c0d67993c97b10bbf085f5dd9095bc52d3aeeef73d10a7b8ba8c895f521aee09c660ebe67a01df3341464f2503ddb8384027e8ec2dab1d391;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hae7fb561d0683b9489a81f280c061b6dac9b0ef4b7dd053cb81ddade3d415697982591aed0e95fe44a629a4ccf4ee9cc0de1525a7addd60f87b219121e97e657174d9a62ab0a5b9a04781d71fe87998515a80892b86cb1d109fd20156bc252d6cdbb4b33401f64b409bcb0c077a58897c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h56f713267deba66c87e9f380e2c07557cc7722e43ce78feef6c1b41a657bcc379a6d242d407c7024ff1ecdb0c75455ba0dad5cb0db7d002bce9b01c17d9f0eb52203cea7eb7825d25e748946b9717161cdac1bd7ca32183747e865b35b1dbba3c536abd5999f9bada943a6bfb45f6b901;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he3e16c20d26d3eeb9127d28d77767e7c06321a8cc2014dcb76c140d6da3d1a8ba14b96d000a833efc5f46ef5106877f202c1b8bd421444f0eb91918530aff6129791fecfdf1270d46677023190d9ad40b782bc52266e64436e28a98f2dc095c607b4bc8283741930b3ded0449f5f96b8d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha7bce5e55cd0edfe1dd3afefe6e475e0e0a662ee938346a8df85f8918698db15917260d5fdb12b4153323454edd0f6fcc6f12ed56e10f99556757c5868e2184abc34645f87d1be1286b107cea787615c95d4610f384fc10a094c3b1f557c2f5b10464fcb59be290296763424d41223a77;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he79ef8a73ac4a17ec540208fc8b59c0ad95ff58a8979ec5fc283d382e092dbd2014e92100e4531cf688a21e43bdf347be1dd74ec8403791b1feb69b08f3dad8a502346f7971f33f2cb0be40a8dda8b6ca4286be14800e90e41518714c2bf88d1e5b976e047838cfe5975e72e575e2a449;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h454c97b4fc6a027f74e027f62f1be2d3ad8d5527d84aed60821cc59a999ad76dd7fc3e47a20a505f1d3273a093ac48e4e98a144f85ad04bc7f9c9331c02dd70ca7c5fa7866d9ae8dbc3fefb61420aabf3c9058fe21e13fc3243e93115f36b4fba2993904d95e9f0de30fc85b4932feed1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9759aa549d168be39724d799a16e58cb5c9f701828e4e05aa4249b93a9744d4affda3dcae235df4d79e072af28edb6483ae95b4e09cfe6c261c0a448dc9714a789f2d87232ab0da7add32b1d18fc82f7c5089863f9714a1478cfa3e10a3257ce4bde4f233d34770870453cabde0a2d1cb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h403f0a5104dd161ed5b44c4bd9e8904005e80ac6959360530dc2de2cf45f79dd39dacbbb6bbcf0bc7bbadf65ce8220253d943ea659f5184a7069faba55384c07ab37d2f240b709caf32d4971e26b491ab2b1810df113fe9c69d2d3104758ef5af7eb57d874093e3df391d4b846c4cc09a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha01eed13a60471e1f7630716eedff9e6d605fdd6ea72f5a384cf4e299f30116ea7988a40ac1ff9c7357151de223b9220bddef966cb18295c73e692f237469e8e0c16a941b1b76d06a602b60cc9e320579026e1544b17c93feee87d328927d4b55046490ec521fb01956efdba634599664;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4b69a796344d731b5f378f6ad98131d492cee9aac9ba848844f285eac9f3e72e4fb36a2d635463ff2be363a6d54b4a7d255efca564a1a3f7bc23534eea549921600107e43b0c01aa573ecdff2abf6b3e1ea7cf5d0089cf007767a6637328b800dc83cad95752d390385facbc30a9d62df;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc5f5324e59ecbac50182e6be2d535054bac4568803c31434bb805c9dea968fb1863f94ba4ad465d6943050b8724071cd2cd02ef5eddecfd071f4e65838b2d68dbaf705654221c74cd8ca24821b35d88cc6b672e48c61123e9cfc549154242eee2f5d0c8218209724a1959205567491cd6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h514854707abe4c7e568b3b4720f0ed63ba23d05f85ff09e8d609b34398ced36807bfcdbb305a3df4734007e2f6615e8b36b2fc3f59e203f935b14c32498ecc179f78dc1c05d5e6c870d8c278d2297a8f627e501220c8d106a6597a0b1685367eb8ca2016e3cb2b06170afe6b99c7a3ab6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfe0a9eba44d783530082bc2f854e7a6afce4c2f94fba4415e9db6dc08d9577ff536023bc63e2191757f32ba1f4df2fcb76d32e13f91c4c9cf38fde1a021d9e4d54d14ffa1f267f514e08bdd39b26e8ee5fac569bd68b88c9739a209cc0a97e426745d3a4508d5b8b66b8b5213f762819;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5fac33151ca82477fe4f4870ffe3113aa7ee6c72ac9b5ab04bb3b6fe19aff54121e6aeed4977cbaa499d75c1afa5041e9a00b925a8c62f63d821a0f9018bfdd81dbcbe4431dcb037364a49117bcc5f74d92e06a0f9a36274c8696aecbed05c8d7f8d5529f9899dd393958cc51507224dd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ccbe0540a9b01630c3a7903a238b2cbb53c5dd295ca0e3a6aef3d08318ae04c5a0d45c1b0d8478889858bdacabe3168ac5d0292f7be62f53cd3e8158dcdbf46df58b59820aed053150604c1a5c103f5b3da08ac91edfff6f3410eaccf85138ad50435c5430f436d7db184eda273e34be;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9d40aaa8b490cb664d0881cb9e537c0e7c9b28ef05bfbe90ceed5aa93003395a41bb3ed35ec598ae660410e3e856ad3f7eab59583f8d693c2b4b01ed3058bd1df1a43560412eef116a93d015fe25f36db85abf7f851aabd282e920e343faed7fdfb5ea173fdfd241e09543a91a7e4d77f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he57544542e944e6ec4df77d6405e6cd7d82b5f05b6fe25d57487e1225b234f07bd0fea0c21da8f35f72d8c844bd2770d93f0404bece109983fac3ac4ace0cae3922f470bc2b1269191fb955d764b217e7d9e0e75a4b2580cfd2674a6af1fa403e7883b105cce6a1c2bcf149ec6d0099cd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d8272e73fef74183b601a19cac53984987cc56fd3cbbb95400702a8f83f5bfb8603ff9492a65fbbd08dcd9fb2848d3064793441a1ac004b6ea6b16f256e980157e656e472eece6f30ddecac0dbb813354fb701c8bd31b62407be76dac81092ed148d3a74506007cfe5f156d41894d8a4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c2a4e2f36cae1965316dab9ed2b93186ac357d8db92be7a5163fae595d27fe82a9d91f01037af3cfaf3e0cb92df2afb7aa701b83123b4e24ae79a0e8729c513cc1886a994c2480a1dd4894d0f3cef1e88525d0df81b7b76e189aa0b5ac6fa729e0d49a71463c90411b8a7287137180a2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f356b36cbeec4be3055060df458ccf4be7f1e698cec5070ab92cc0b4236782317dfaa9bd081b87bda29edf1aae33d943d4e3df1c898fb6556a917f6d75032322e4e20975e10bd079dd34a6f87f5254be899ef0d001e95d85b6955e06822cf06bdd6e089c4461e5082e6fb269a91babc1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ac56eb882b611481ebba52dd87d2683ad65e5c0a345e9b1069c67d78cff66a76a4b8a5107eabb9e8ccb3e793524307925c51faa288e165dd6bc264ab9491c86b859a3675e1f6dc2c8d8f34c685459bef207e233ec6f2bbf44c0caea70152e46db0aec7282d55233835649b8ce784714c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32218d771c984febe4fe27c0cea5c1cf08868caeb5686b3fbefc4ac0d99712d7a8cb0be136062ab573527440c3ecd43a424c06607afcca9c54e6ba768652cf69b12fceb6f37498a1da48a6fc331e646c1a9144c0102acd2d02cdafff7e3d400010966c84a85dc57ecb33afa77e5ac1407;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7451ef5a88be4ab495e93f777ebffff7405176dc7d59f2c8445cb0e272ec0623c82e83c831262187f8353dd18278e6bddb220fcfb9c9fff8bdf689c41890fe4851cab7464f771fded454295b1a4d18be382ad0a9eb0fc6aa47f51a86503dac58e15aa1f1d2c0794b1e5e38888cb4923aa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb98a2c1c310cda9a938edc3fa47189d93aa6a86adad71c37767417ea8db7f4950f7bb1b5d6b83c81f07cfeece4f6e6c336cac9783f2a257cb5ca1047eb892e0b5707c93e6cf51d9db2679b5ba533ec0aa170306186d3402e24a720d545d778c9aa018a530ab9995c1375cc14503c2d18a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8df337a9daa48d85e74dcfbdff9d9b15a156d7b3a3d033ee3b36e1819df010f5311e586c9f30e1c5c29c9d7e9dbedc9bd113b1d06f4b66c7a6f4025c3aa5adce24199c73d1a077edf509d42aa7cf05f1e83212fdeef9f36a30d1d05d4f72d78e6b888a456b48705a5f7f6ee2863c75145;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd6db03e8273bf2f3fe8910c915f0fdbb870678c11ce4fcd8b655cdf18a99c58b6efcbcb38cff3815877340eb54c537454547df27e3bb1f12bc5edab5fa3ecbe0e3e792ca6ccdc0f99e108f0ae21ced4086cc440154437e2c31e10e5144d4c7095fdb193e05aab215063145d0944eef99f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha145748cec63cfc3c9767969ab9b6bfbeb2a76466662e1ab757f6155b40fc80dd986ce659a2265605309e11e8368260a908e3a7cce26e07d071743dc45bfbeab414c270796aefcabb92c0fd2d548f652762b1a597d1122cecba1fa9a09e06ffdbcce4396f5c9b567f201ed3d81a7d6dbc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd5e00fd8e13d0b8c7e778afc557d333683bf636553dd1268139fd411e78aa9f89c3e5a1d4f3b9aad3f2edf374065ce67f4fdf0b87db7d68a73b815e1c1871b0fc98ef82b2b5929ec19d23ae444ab13c14cde4fd712f13d9ee187890d706da53766bec790e43145c44b1cca957e51f2777;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbcaa2ad25a89bddd948256761399262d5e339c8d667cf9be448b86c6fabfe2cc76bc72846b99c534ab87965f50da16ee90aeb35869d764fcccff6e3dac4925aa997355fdfd1b1f0d19efc305f5225ba4cf510d05e5089d91edcd749309e38fce5a4b0d57673aa4c02a34e4c21cfa1e7c6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8a860268c406b912e8130eaeaba79db1fa33cb6376e4442c6c0fb896487176c8eab43b51c7d9241f84a7b6720e1d7e09f19c3ef2089213697fbc1484ac93185d5d7f53c0887e2d9008cafd2c508b593e59d79e395b076c800daf2e24fbccd3e073933613816fbdc3c6eec7d9ab0871824;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h729538e366e390c896f410d606a395709d316b6f83b53e1958c0221abc1c27b5c7d6db6ec006421f706ac2e9989cd144c0768181133392d7badbd21c407ac4436c8c3a265c05712d627fa496c2bd1de52934fa69435e67801d1466223468de4416451caf0195319a01edc6474de3322c9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he4ebebd96b2deffd6100102f01d83159e30bd5e413e47e30ebefbdd1e950b31bed6ae35dc5811ffd4640bb35200420d6aa5f5957e3fdc5d2cdaf00c1f91d72ba2cdea301bb13390813d42ca56d9e39b063a9d9200369a23f77cbf31aaacd791e210ee6fae5bb54133be4c780080dd308b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h677d01d887e9047dd5baaa2efe6afb73ab30db01be92e3fa4a45289873baa63c7879268409420d71808705159152ae4dcf25eb46fdb328055d66fa0b5e8252400bea40ad2745610ecf4915eb7b5a8cd11a7839f01b0100a52163e7df863521e2f486f946014c49b557964c6dba7197c85;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hefee426cb7cda0943d57706c124263544435c8787a60986405a11544a03e55982874286310a75be8600d8a7ac65f36dd6ddfcaf58a3e3d4f162b62ee13bab702d8936bba257044bc0d370e74f517b2575306302a69733ff27ea71787b7e2a799440204f77820843c76e5de7c4602b4fd9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfc93b7777d4b5f9600ca98ee58bf48d9b1b004bfccc0960e3ee9eff84f3da38edce61a6ef45b55d9c57bb7402b80b69e0edfac661a97536b9c20be4fcca2506602b06a4d775ff04a46792cd97428470fc33b1e9b0734fec28e086eeeae865f5ccbf3aefea5f40f1afe179e54d378331b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb2376f827abc684fd12514a124544854066d2920ddaabf42b2dbe3d40329b8f5f54f25a4d631a4c028aadd8d209049431d4eb6e3d1cc4be7ffb655e5206ea49474f973a3ba6ce3e85bf586b504fa693d45cb8c49fab99390ff4e497d25d27ab27c7c3f9666048bce3f93e9ad18577d51b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbe46e3ea5b9c35eb1548587472d496358cc76cef1891fe53c380c6276a9538006c972b51b217999d75c2d89cf8a846ca1bbf74437c9421428d410e7b3e19b073c79e61438d5ce069b40bcea36663ef4e56d159dcfb4c39c19dc658b305891dbd8fb652d37aa1d0370e62818a364a795c2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd0cacbdd1281d18d9efa874dcb888f1840faa7a7446f74c1c57f8f761d6ae4b831b17f8836274531fbb872147bd17d3da0f88a1fe5b1f6cd1d8fe2fcca85f2e8c13a57b933e802dd2249fd2e4ed903c0afc5ff35bddbe6be80c7565c698c1c1e6bb9ce9ff4d1d802e820accb8ebac4c8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha54f7618bddc140afaeb439e6a977bd667199cc17d71b03ca6eb96cf869cfa944378486b15b583da780a2349c7d54306b618387db9bb993a043f5c0185acabc132c68d1d21d4e2f5c9dafd19c13618134649963671a4e969519de7185dc96d256dceb5594685da3b4b629259f32e92e2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7464e5aa101fe5e269afcfafc7bf3c6ff186e21c1e6d70a9c7990408bd0a9c959d8ac40ca9c4bfb935482475370370d9174122a95efed5a21cdaf77c9273505b7a50be7e153300318c37fe658b7ed3e0ca718ed19990c87b05c87d6723efd2096b5c0a703006004f6fc2f2d5e1fb30daf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2ff2252be5fd8bb97d895ed5d439d21355298e7bb64f4c906c533fbb6a0c9bc94a4c6ca1d2c468044386af082d8e4b0d4297759e74d4587ee7d71102eb36a1ca196a80f9b49226556ddcd81d9c34eaa23488e6be47cd8da219f0145751246598cc01944249bbf0a939ea6ac0c635fd2f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2cbabf30a16dd32aa364de2a0fa3fc386ad7c6bf5a57e27e12784281055cd168c35ce73e74edeb838e9a0141dcbca1a48404c5e1c3d3d498b6019a85b5634e21d62d74f07a65e3ddf4ae44c76a8d9a5293b7dafd64c82510742c7c9803ac93b3a655d548ea2588cc920e57436a6bcd47f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h37c1a8bbdab3835e2738453a017a850381cb0414056a238d9af2627200b7b7932350b269725c47407770fcc20712a61c7733bb8e3ad1243a176f119d19fa8bbd8b422c66b268e1927bb1d2eaae232f1bb64d84bcbaaa06b420edfc0c890dbf4fb594013401aea6aeef730f0b177f1fee0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h41063d3865f07d87267e10e8174f0171bb87eb4e1f89f3d1e75bc1e14a9e7e249e8a0818605f5da5a861a24a96b27fbd37ff43194883c8c7520c7c3f638c706dc30f8c97b30118a8945034ae06c86228188ad14767da82bcede48ff34ba04e44a61625c7c4e3749338716b0c4d1aedb8f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b17757e40d0ea76010f7ac707f8720e81b114072e896951fad3cfd8b8bcf35e1132280e461db90ba9f09466389678332104e5b3166782c9b858f8f2209c665a20b93ccfdc5f1abc5ade00a261cff9b045b6dd0cd5126f9e8266ae747d75f2cbb8bfb18a7ba9201dd4ab5aa3238caac24;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8465fec6bff0145457735ad7242a71ba7d472b08761eb34d6a57813ea9968b8af2a9012c34d5747c75c1b2ef5e799ae7e15a6dc030ed6168af0fb90dde3c89937b973ce94b385f3b2970b948cf06f3f0d454af57512b626f3675b06c72616c5cef75bf5239ca9a425fe70fc3620b3c249;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h43b30273235d319fd625512ce4b8faa092fec8286bea9f967a84e2d32a557ae606994341edf2ebefe9bcfb2528439138d93afc3ad6720868fa68ff8b297781b1c8064b437f5d0af7c8ed5c0adbe668920590f3709b66ce64f0c8091f190d5686c4d0eb4f68bda28c99d5b3a21a78c6c50;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb64a89626cda0997d044e03758101cb2a084aac1f815bb55304391a1a4a733c0f480c08d3eb1445e7545a0fa2425198eb169bb93ec3cd75354094136b38e2f8653a418a056e064a1c29262f988f13014c4b817f58ea0acd983f60e314857aaa7f7f159112c54fcbca37f23c0f7a0520d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbab1abb980e02fd57e930e0a299de5a54c1dbfe1fe896b7ea8bf08e1f3c5c02070c3a07fef9df298d04f5656118815f76a61877689880e449afe518d5515f9e0c2510ab8ad685ae8236b18c4548fb36a9166f21da158be0f8bae1efd742b8f21d550fe92382c64dd83e920566634907e2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h566f48fbe1807e24ed22b7b00186d808c2015e41edf1e7918c5997e0e4b38fc383a460ceec50dd5de1538567beb3b17df8b973dcbfeb9ba2e480ce1342e0cb12f12c5cd75ee9489be9eb64ca7c6d638dc055bf4000e53d86d07513a5e8b439841c33faca2e9ec3bc424a6b9ecd2b1c1a1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h896b4c3654ea9cb107ee5305d54980e725b16bb7060271eb6b077ce5c0971f898c39dd71ca499b537eba92aebca419775e3942badabf55b373ec2936e5a84ed97692d9913f4a1fd0137136ab801486e507d4176cd6502de741b61667e53275377f8444f02d0efa2d1e4111cba09450282;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h779b7562e9106d41e4ccf0a132e48d6a407c5d6d2e989b5aeea451b5ee4c16f100b1888efca73db8a3f76b425d5b0f3752944bc97ae4a24b4b7f42301d5ffc11d67eb2acee4a8fdaa0be13da4837a9d67bac694d40ce4d5af63503e2db94b7bc01cd8752cbac83769f217c1971b27d150;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3e536ef4119d56961c61c39b52bfec273807e60f9d11d4c23a4ac528f06120f9c1f52ca99646f0aa0ee3a4db96e4a47e1dd127605f8a07c213dacd72b6a6f6ea1e9d462be4730f4794ab95fa9f9e8b722af7d6a046615cafb0f74f5b6916d941dfefaf63c816a57fc1c7ef8a67726c9ab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4c5f38ede399d4c662920ef922ce990800d9eca89e4fdf7e67235272785122385f1659136ae5985a212e3821a9b3a8f333f921e8fff36abf780cf1a67615ebd8669b6e1052a0f51895d5cf5d4bb0303cc5ee9eabbd56dd9cbd05abe5fa3e48f4da114174c58d98a64512cfacb9a1a1830;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd86c58dedbf463115a14a086d065c0ae53e8c4c05e517d10ae92ce182746d4cd98b02fa7c03fd69c731f0994511e33fd84e219f19fbea2a710343679548fd70fe58175130a9bde9eb99603be50e017f5c7351b138970ac9a544cef3023e8f44389f3bd9f04d7874dd5814402b749fe394;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c4e35fa08babf8f738b6c7f0f55ab5f88c8c572d8138d9ff37292c0a6105abf64407be60d2d47fecaf7a3b29dbfe975df3aa86810c55b42eda42e4db58a116120ae1e7a0b27735875e8537e208d1953146c9a73f2feb98a5d6ea98996076db1818f27e0f19ddd7791b0f9ded619099be;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7ddcbb2cf9daae4bccb6f79d6aa0cfbf5b3f5456bb02be30eef4124796e1ad4b7c7e04803a5e58e6fe4bf7b09c70a57ccc68e5888843e599df1f87282738304af2010802e0ed6f42e41df7aa5cc694763bd41cdc29673ffcf7656b85da27587450bd652d47895c9eba76673240057b893;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha03f488b72be02fc9ddc6f5032bb0efb4576aa832ae20afa8d580d05c023056a7fd174b80b52faa20db4ef252f1b77dc6c60956ac16ecd12bdfe114728ed16ec7c166ddab8338262f775932755d0cb17ee6e77581c6c7b30ad278d8c3487d0b451a100a549f1226aa6dea58190b6d1ea3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7dbaa8748e29885e9fa4e48f1161849c4a7a28025cf52daec4cc6a801dce40b143fdb31b71ed7ffd7d1c052ca58210852bd961cdca3dc5e6f11a9fa61236e457bda8663cbcf32db0acba658dd9d8381d8b7ad11d2b2ed5a27fea544d581815608f5c31716917884b0513a6dd141f0270;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc4c6727e1fe48e7c09fe436ada3bdf8dcc2ff7b63f9395ae91b9bd3bb60a696abe34c8ff33849205d822796403a23776a0e02096a7370c9ad99866f5e83859afe4f88026485b935eb09af96b4b287866d8f61e223ef7141eeaf8d176858cca2d4e342af0701ad7116aa2526c3d190f423;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h165a7ff9577a9200ea3d29b8efd57d6cb1935871e86744bd2f790a1c113db4fba4adcfcd6f29b1b711eacfb1bed31533f5023fdf53bb8b69af95b1f2e625f565643c416e2327ba2afde7bd92dbac38bb31bdc65bf8fbcbeddbd9d5ea9f6e39120ed2269f4745c056a0cf3db9e4b5ac850;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8e2f7c63ad13706d1ffdcf0a6d7b8907522c7e02e0b155bdc4b3c395cfa8ad9e5e68328dd7f6d70c3905e81ef1586d754d4efac9ab15ec2d62202a6b47a77f02e92ce096d3ea5af7560ec1f77539b7bcca7702763796c5cb3794d06d649f90619ab018b160c612ef31c64823e83de044f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he65efdb917797a1270706c90b7906cc8dd15d3549275b0466d4ce9ef6c8efadc28043a169734554d1383d06a937cdc6f89e421f269bb28d6ff0d0707f5572c1576418bfd5e5586bc6bfeada8b1a6386b79775b30df983772a27f2e74c064dc47c591b8877f612a21febcdbe5bad9cd70b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe706c450be8f8a5574fcbb755ed487cbe62f0343aacfb0655caf8321caf1be05e1a307457d236ce9158769852282b5b1395a373d5418ce4fbe371b178385904c912e7657bd1251dd6a2415f942d4df77d90633d7e21b9623fd3305ea511640f665db903021894302a6c94133528292cf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h38376c8186ede0575bf8086473f797cdc3775a654f4bc30b11de69103235c724cdd49e2cb9261fc12942d31578aa901f6fb52c1542bef357f94161c299d0da9c9437bb19dbf348066386eda69d79815571ce15104567448a5b01c58d22d0428b65316aba50dc804042c45467d6c193a52;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf370eafa036a7163192c985ccaf234565d83fa468f3a55c4a447653e272f7934466be815192f88e963e1398483378b40d12a12e5eb2dfd664feac9427d26d2273a8eeed7c6cd123963464105474e7dc8fb576d6be5415d6692531dfad4dc58a9f92333b7520a00e0950b109617b64ecf7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc1159ff8373206761236becddc4dfd42bb7e806130cbd277baf15d2f3d69390cfa06fbbdde5b76e5b4f19a669a1cfaf7d5307a9df0127c5d87e0b5250084cce6583a126352dd32130a047c2c785f09a2e3235a1d663ecd70272b76397418532dea20b703db286fc5757b60cd6d3403ff2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47ef2e9d59409c17362ac6c60f1bdef4a6856c225684d96e72704b089c525c8c2f560f5a3d63f327a69c2003b5fa4b0efdb23be6c764b5938ed27132ba70713778da331f22e7bdd34b02bf71d585a50e71a6ac8218e094d6a7795f988ade93e53ff8bffa23d484a7c66899693c1c5d934;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f713e0dfa971581433a00a36322cab2e37087bcb005163bf4bf27681a1eece2fd6ba1bf4b35bb31b59493c1a7fb52fdf5f0f4fcf154ff61ac040edcb3cc2424923df3d19b62334a67278a4cb4072c9d4118f1e6b1df33da0423283bc26f118fdcc87d713797400476c1558e0cab75f98;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f531181aeaf49ec55d8cb87473dd7240358c8a9f2e25aac46b374a98b478b341227f1cfd34f4bcbd989b4bb268f81ad1822fc7336a7505fc94d3835d0a134dd8d81db1a989e42ffa725df516207e82daabb7cf909c4e7a7ecb570d20d2d57cf33785762801db965fc7e551bf17e621d8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6b18b810f35c1eba58537dea2984ac025bb8e7475f62a2f859472a819de42f2c201869888fdee71b1cfbe74792940a3af23eab29dfb5e7286b8ed3a3ec2da5b204ff4285c656d683e786cd474198534e6cb3f47b54d370bede387611d22b946e1b705609665e68fefd5d0eb8a7c210d80;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haafb10b33f12756567d7fdb63d3acdb5afbac835016826afaf810f8a1ee8fea2d7614a60e78704f108ff29140165485df8cc2d4fcd84b81c226f59dec7dce93478be76a62d76fe5346f62f901e207e0fd4c27e5e3ab205581d2aa4a45c2614e14f4929742c214e1a96508e7ef1fc9a937;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb7d30a7296c8ac7ce25a52e86776e34b2344e3f3e900bb7b53b2fec9e1db9e55ce4c3a9026e5a59dddf52a92502947081eadd3844a00e5d845f8e61782776d35a8d30fc53f7c06e040290ade55ff61a143ddd341115dace766b67940aa785745932b48974f5ea3a213363aebf6ee92175;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab3ddc3023379a354069bcd3f9f69bc75a3548cf17985207cedb7e11d9427b17b08356ab74ebd69069c4723390fb9e81834acc8acfe9948163ba3999c32a4b8c885e1cf76886e9146a2e0baf6f6a78b86049771e8d0f1b730841dbf388bc0778dd9ce18b627d2415ada5d3bf6b116f722;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcde0bd9f742aed677bb12664ba5af68994d61788d4a114844060723f84aa7e723dce8167deaa6f3b32a6250846b0bdc2e114136b2c150d6436865f837c8fd22600dde54a4e9d61552ed42df2f41f8fae5cd61e0ae4727af0ff6e9b29750a2079cdaf02d42f2c73e887cd5c01345823c63;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h58db5935e10b94f2be438fb84e5428256313d0a26fe5757abfc7a051ff6470a34d2a15d08d54738f243b71b329305e510661fcdf842b9aa25ef04b3187c02d86862c10fc67359a712271f2b17a3cc40cc39c0ea217bb860cf0268dd1e5735cce4a6402a6609272af7bcd2192f48435029;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5f348454306e824582e4ec70eb9a45d79121287dc39c029960093929d57c571da39b8a50a6372fcd4a91758e1ac2466c7daf25f8a9779d26259c3b1da3fde7f98c8b32a3c26b98d4937398f56a3605392108ef17332dc34ce2fac03b3842078d8827e74c343b1e5144b480a4a3f58ef3f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h70745a7cf045033d186c3d7df6271b7fefeee8a6f380a671153e418728a975fb9d68e7b28c7d89f43c4a724511012f305c49e382172e7b1883c4eb25c744107067d693fcdd79e11e8a806ff169d23fead3a9d05b9588d3aeaa5498681128c5e19630126a790ea41c7b7b105eb28593abf;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf338a32afb99f32cc2d36b27d5a93dd209bbddcc360da54baf7ecb58d65dee135e284e2feeca39e55eeae0635e5c711fb556f4957575bc9673b916b20f84d7a27989303434d30be2a5c9d9fb48d095383f12a09de1828dd3fdd14df6b8213f5418114342530bd162f1f73e479718f70ea;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'heefd1145546f90fb780a845ad1c9f5f85d4cb0a7e72f5d53754b7cc090fa3c74daa63412195bacebcb4b0164401ed88027f2c6000c34bceb2e2be1364b0795db229d42d5cd0be210e6f2b354352a8c48ead918acf4180165b9bd731f6347e1f5ac257597093b8fb1f313092ba570ff43f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h854724b494a6ac98528226279cbea1670c2c1eb9ab0163a678a122cd4e9e38be98cbd02ee0a1e437808cf28e8b50e7283c77429c2549d3ffb5ec8b5f286bc8d83dd06c25be6b24f75910814efc332bcd4c7c11d2c5172f873b284bee72aa6996d7db98c98de4bdc7482335bbee06f74d9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55a0878f38bc958bf3c5ef4f87a15ee32ba719a9fed9142fa63630b9050e1ab95a6f797239855d89c81e0b6df158e34ef2b74c5cacf7d81a59b26d0fff96676f2b1baf68e1339fa1433d1e3e45991fea5bcacc6706cfed5a4c00ee28b45f14b11b7769b58296406a4bd034362fc620fce;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0b77692c9df72f590312853166500b47a290f37eefa0a9fb709864caf85dd896afbbb85f36f251648392065e392d9fadd8af2bf356f763407d9685b56278e077411b21e5a2c8a2223366e1f7a5d840d1fa1162b7a8c73d5f096435dd66354df19646c07d6a286afec24a9c722f2f7bdc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcee5b6242c90ac6ea4c6219f69c496707d2d566bfb9e98d56c88245a495350974cade72bfa42b854bf5e08e4efcee051745be46e8e0603195171c71bfb879c9a32960111a7e09ef3b6c4493f7c11f7910ad575c6b43711a0d559dc8f72df7a3e9b04fddbec0d98821483cd34098567f16;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6dcc5c825b1b4118ab9bbb2d591170ecdbb81e16e5df9e542dbb15e9eddf843ae657d7487dfd737823a6d5f6504b9eef116ab0c5c06ed7560f1fe1de0e65c89df4ecd076c8f719ef5792814aa00048614314be0d036ad620ccd4f3f8699b4ec86e8191c453fe4c2ac7065efdc3b28cbba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2926121032eea5865edb266459bcfd0b452877b8ae903201be2cb845da0430a77f2fc299657b555bb1557872e1579271fd31fc262ecb81fc530e5093039f9416248e6eebda972ebf6108c00c07f00830afc3391b626c5a99b3f723445d426f7148882c4a42ae1d10be6c072bd04d8823a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h548ebae9ba5ee144bd76db6a101623fac6082aba58e1daf3a8c58f8e212425a335c123ebe48b690123565ef04b4251070f8b2f3414163ddb4b2b52e9750c98d7a1306ff631bcdd830af27d7991a2f354eb558f1208af6af7f2010ee3060567f688154e2b12db4eeec2d0380cd7c62d3ca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9fe1922414f719a2372db25042dd5fa51f632e7ce7f25dd4415187b1e6749f31d56da45a4c755d6a9f3c0eb9f2e63c81272045ccc21642b99a4a73c5ad9d4c48b5b88b10168b52f7112a69926b48961fe5d876387a8424950e716b5c52394d04d2133e80b57a53535bcb00a1d1229947f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd9c083c86c6600af6d047387c64de4ddef4955d740e23498e578579101fccb3f8ab2c2982bffdd0f32ea4ebcd32503e4a96e1394a2e107338d854d24979962734a3e42a1632a3b0c109bdeece000efefef93d8b6af0af1440687b07a450077a6cc61b1beb40096a5bdc11f0a0fc9f5c15;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h529607b535fdcf1e2da1a6ba8e760a63b355fc00d72e45ef33b821562b6f34fd5f1de9ea38ec0b043be6bc89752c3d937762b892bdb4433337e54ea34c72792dc5a7117b59a3a0101aba0b2c483997d62617856d37f0a4473cfd1e56a0db1260e8466f471767d35f2c51aa3c4bc8c1241;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc492a0b84be8c8e75469ae82c3eed9e314646b4246e021ce065a729f2e135172327349a71a239b8589ab7932d8fab23031a7dc255fdc1f3dfd710dc5fbe7f38b26649e4a6eb352c0de3e5c949ec8732567417aebb326381a076183c7adfd3b1448ce7e4d637b0131a6ab8c58e9694f394;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd3477350680dc43618b98ed1da4283e9e9a4011f325fc59ab42e38bc8b6c68a2d1671895c837d9f2d25e52b7ffaf3adbe7f6245753598ca3876769672dfd437ec63490ebb0f22a57ef1c161ce56adcf993dbf68af5e6b9c8987ea8b98ca146a8c33a594029958cd1e056970077a28780;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h180eb885da5978d8b218b2b262052efb47648bdb72be54779320a574b0ff1c2fcd9876278bc9143146ba202a3a34bdb6eeab5921cff4afe51d131f02715ab3b1096faba030bc2f6c00a25e60c202305fa34db05e884d40ec4917bdcc51ce5007f21fd716fa320f71d33b00e927b0fcf7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h691250b0fdd1a97a0c95ce0172705d22d77f53c6b419d6b1804fe2f17d5b46a6dd33ce30f7cbd7ea3bef0c34912d2d2b2094703990ab744b9adf9b970ab44823bb835cc58776db5a889390308c4902dfc9fb9dd9d3e81565a98a04ca855f5a12dcc29dbfa5dbdd02f2b7de9af1ba1a815;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hccf91e2a0b61c49227ebffeb52df80735eb5a82366bd4c3de2363444e2721543cac0e1c3e5ec76149ff6e6fa1d941759bf94431e33c34ce94935e9e6a9933c287685d0afb34ab5b7cd91ebc9422bed2e422ecfbe776e91a165c711e54f98a54826b721d4229a79258f734a8f535c24ba4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf0f5467ae727dc50bcf6f40f3c0601ee56afc94792b76d53ad750c1d0dec68a9ecb9edd8d577a2646deea2c3d53ff8b45a2dfbaf46249a766839c0bdeb77115329ddc0961c762b77c9b8cf14b976250bf76158581808ce7033502407dbd0020e1e5317341a59a2389d370f843ba2f434;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h440089b4d7ebaea2bfb3752d7beb700c21109d87b040a77ea433dce977b18f5b4805a0962bdc05539d8f2707aadbb25e770a83d8beba33bcf6beaa5fb295d95b95ca232239b3919ebf500498ac025d1f3a1f6e37ec233e24346b028faa8caf94f931e65a4fce4557cfeb089879b4a13dd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac1ffb7a7703e1953a0a8f7f4b4df087e174d7250288d966620e2ab5680e6d92389056a87caeabbd04d561e820bb4ea66a0080ae9f494d45d9a05a6aec8e5d26f874870c99f12cfb28496e27bf854d0d7b006c9348c424eceb4e13f171459d11d9137def5e5b3024d1f7d4a331b8e0660;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f239ceea66b25f8c995084969cd3d5bd1003e2b1a111513d10be919eb39104594b95b8d5f1cb5ed04410eed3752a8590b06dbe8acf0c9cc73fe0c6096d80c169bb24c99d6681c85dc209e7133a3f345474b4fda5aa9ee7c2bc4f206602de18c0290e734110d88133a39adf4343f08cc0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h447e739daf7562e4f0b3decde68021d627dfbb822f4ad60107b936d2badf27b9bfff8b02b47f5aaad5d89d69e3077d7d0fd07fcc7f02c9ef72e0d69ef399cb8d7ac6f598ef6859ae881a075061ec358e62d7717355e08b99d7125e11d1b77c32c3843447818907594a389f15b89938aa3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfaa7e35638815fbf2c166ce2fcfbb5d444b1877c88d2714fe7a4ad313e9180e8b1b1fe491a822157b027b000d5c1f48e4a47fd4da48343caeca571204d167401b3067f76d71565a35c314fbbd5e12229d7c0223d0087751758b5ed692b35d1c45f3aefdb04cf5969cabb221628488e638;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha11dfa876cbe12f9d3bc8aa2c7dc3dee327c3a7c74ae0188de0bbc6d2d3ad94cb2f13a2d5f9cddd219ee50c04199d431da526f2494f65504d1d57aecb553865fe9f303f65eb8f044d0fba42d36a3c5073156cbebd2d77c6cb7654ee9d1f8e352a0d8ac502bc5aa5aa923fd165e797f92f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h328cf2399c717d87336e2cc78169b15254cce5da732840c8cf33e38998e04e14d73cca05c88591f9067614df2180d3848a2043166423c38cce49ad1871036bafb4a2de9c14ab9b5d9c7bc2925bb57675a5912653882df7e6f28cdabef9046d46e58497ad001ca3a6156d0cc97874b7b51;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9e13ada25cf5dfaa304df611612efe58f849b880d06cb1c8e1875614a5cb82ebdeaa873b900ece1032a6726a7aff6855f839aefd886790bd3e263a5d1cfc1fd0a00456bac62ea83ddabf01473e731de24ea76a9c92df42bea0b0030e490329708d54fd0149744a12cdf41e74bc73c1254;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9804acedec388e8b426779056e69fb9df7b8547256991463f761ec5de0e639fb236359ed844e3c0808f684f9c3dbb31c48bba5ec1b3c98ec64d5c7add2f902ca1369eda3df9f50896ed444cfb48be400ff93ec43c28da29b068597dd319bd355c01e378e84d006f7a8620e24632103b01;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha46f0c35ba811fd4347bbca595cb55e7c7d1447b5aaea5d4616e6e605cbf0f6102883b24c1e2ac6889c9b86c9b8a3a8f245d3f983c0ed094e5f0d2d36b58dd1381d4bdd284a9a76b9d48063feeaae6d9782f0c293b23324ccb7cb75377d3f094e8cc10d779c6b7e337eb6320545ea351c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1054156f674ffd7339229ec109accb3c453e83aee216a13525af408a192f5861a220bf5ac570a158e1a1df2c7026c20250aafbab537a30ae459f429737740b98d9240c503ab320976728f4f73569cbdc9d0f3687c605e7736a7c86402ccbcd17a0a854ba077a5ce8a735e27adc2635a9f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h88a6f13386c6af09c03ade492392c2acc5ce0b1d2f4d7a2e22ef2f85a95505dec922d4f51e214a9adb8fd50683218ec7692761e43ead3a31f01f6255a5f82aed1ca28567ba7d4603d7a0dd38c46f78015bb708b82c8ae9fdd89e9b7e0c311582be7dd8b92b5fef05be7384ecae9157010;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hed7946df7671502d85e2c33989ab2729a7d47540f77a3e1c28c71ecb992252da7e30df9f90d578b9f0179aa3b20ce0d18f20bcdcff645dceebff6e7e63f35c2be84beca639eaf4312a432ab0f02a44cec672f355cfa4fbf52600ae2a398234a90638b4935aa6fd09427e5629372928426;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h248f613eacf425c09d0475677ad91696464f189697fad846a64068cd5b92557d56d3ff3d35a464d6a88f5b51b0dd0b209a917153e2fe6dc235e80812a63c71571850aa9855a892e5c7d4bfcef84461ec6f48a5aab5308f96182b613fa073a1ab6e350d6873cec99d239013fec0777cada;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he77338fd58c623c1c3f3e6b0dd49ff4700ba566d85bf3ada3c5db280aae17b303ea6747cff95383818c13b3005c93a158900fbb0c9adc14e34c65e77e8d9fe1307d6d5bdf543ee673394a8dca15e9b11364e8f1d877f010e8807e2123a0e0a6703c3518be11550e5b0586a5987de7af12;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he301a1ed42356efe187fdf8987136a49267da9dc5aa35c576aa740fa91cab5ed28a7ba9cae9f82e2fb112958c9c9959d6be57795b0a7de901002eef0183a501735c1deb79361a4fa31c880f13adbfd16ac2c4aae328757d1e1f2b9dd28ef959ebb57ebbf946ccd76c485afcce6b7eac68;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8a91390bc2ae99beade086a312b58fb364be3d32cbc62e3eeadc84a15ec7e9337d6a3e0048f2585f78808ec137a91feb50fa4cc9808a97934370239e731bca2c8119960b46b42d894f974d93b71677b3fdf82785d4872b3eb32b0cb943eb567d632aea949ca6fc2f3b7cccd5cc826d70;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'haf8f6d129fc7edbeae4a02438bf8a8d008085de84bff650c4a8fa9cb415040edbd25a69196e6045680dc3bd4ecde38ef0c9303bccd071041036f144ea246864f9917dabe17cbbd58dd31356befae54099c431c5318f8e231f0bff5aaf4aa09176697c86fd5b9a8dcd20f36c1278c105ef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd95dcd1e857a89ede98135026b6f5d43d3123905beece557217f9751c4bda5a0641c5ea799722db07fedc8aee70231042ff0d27ad16b570021f5832709d6ffb056a62bcc6cc97d8e8f2174adaf89b721a60726997cdbe35286ea18fac6b7cd14c683a46cfb5efd8119f2163fcdd3d9864;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d3bd8ad65bd6cbb4a3192974b5be2eb53082bdf46f622c0afc844189ae42a692674e24fd22140803b74fc3f7dd97d3992a22c8c7f8f16005fe8ae7d8a11737c6dbeb7f8589f578b73a57aed08d02713727001a5905b7a7ca4bba8cd33930ef915bf641ea1db5cb7a1f65223d33cbb0f8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbebef852b49b00c42da596601769969cab17f74b81146cddb4ffedd96d3ab10b879db65e54f3e425a6f19d9b4f9f9c01b4530f7ff2e28bc5f70717779d925315c55abd123e06ceeaab97b93ccab24bc289b0882a729fc8115eb02b04fb58be71a53c3e0cb75b7e839cb18063e29c764eb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbd256d3641fedac0807d34be22c9e91555baa2f35bd1e99fc08d9443bf0f816887f36e596883ddf7c68c74314f0a5d6e75a4491899fb5443a3df76d413974cc29ac5a2379c449edd18cee2ab3450f7f6261e0834b282051cb1dad4407d9724bd9621f2d352ace29ce4980df7b56e7a49b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he8eb8eaebd6135a97145ab0cd5cd606027eadcc0065afe11d2d99a95148984adfba8a2c19c2325c6520ce8a21cab18da8a1accec4b8c11f7e4b30a3b3d98b8d043a827222605d0aa29386076edfd91555b6c4da7936c5827cd2a23b1e7b6bbdcd6bc764456497b2baee19a24b39a4ab9f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7d854a27ead1a904ecf8085f72be768686ac016cc12c682c12a0d4292bdfc43071482b948b32b578de2f4f1d8e02518a287d93f32fbc2d44725921e274b5891fae9952c96d8f8d380496d1ac10bcbe92d6f27c447a6aeff747e81c65d3e8930408b7066471d16478e079c2f89fcaa8c81;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h706889acaec42839ee88180e648a0ddc094c980b907c9c7e9078ea28fc351785ad62af24fa5d7e69268a1c1fb0482edc71d74f72fae6cf190033339849872cbd154943777fe623b23c00bf431b6c1035eeb3bb659578d78dcf5f84913bd1110ac7c290588218022de354f4a1d895bb38c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h93649c75cb1573f4f71abe81335f1effc981e089ee49cf1b57d660216036b5de272b7b9eaac2aeaa18319bc639ef2be0884ed1274e0e9a031c5cbc52ae332b9d5a0672756bfae3c85bb0fc513dc46fb7a20b0c905e3a030120e8099c18b9496c446ae1d34488456d2ea40425fdd765f6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hff2b0838ee45e7b680f48bfa46929a551118c9d21a6b225c540e9ff1917280a0beb2e5e8e5e3e9629d170e647c46230e24303397669a4b4aaf8e17bd31b54ce89bbd762e1f3cbae050edf5eee0f967b24f07a0793250afb544290099f635e1a376dbe92c63776e85584a5e248397e6732;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d69d7905e7ee6f6d0e9ad53f997d14c6135f123405e3ccd5dd96563532b28fede527464c90f677bb8fd8f03236b682f44564ed594137e7680f8f618c9aa0574b08250683c8281ad942bb41cdfb3865c828d730855d417ec1c6f9cc0677b110b4ba7ea72a8cd8662b85ef8ed90603ffb1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h234450cf3a7ce138dffda4f6cb8cf4c680604841a37e021806be8a063cb6c602a03c17730305348b90bb2776f4cb19515a2660ec9422d0f611e31e66ea98e4347fda0f4339bfa526373f6e97df60d52043b09ca645edf864bb05f67a87182eccd983b281d0903d93141e50c392dcc7948;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9148a10408e1dc9704de9806d1284adfa92bb318bc321f633fe43d3eda08b4ccfc62ee8a10861f1f8297915bed54e37fbbbb32c25a0c7e530696b4511cafd9dff2eda945ee1875494bb841bd9ae92b3baa4d9afb243ab0fdb16069dfa026e8521ab458c267e0de90eecc64433714a7934;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb74ca7a76261b7b84b184d89fd6bab93450c7ad71a890f9d65af7b43bcb674c286bbad0c1845d4876738ff25e3e6c0235a01ca90b0923381525d9acd6e62694eca8ba76a9c0a2b4eae96a6e494dcbc4ae995e86b858e7988e2131a636c1a098023f123948812fe742dc094da8683d982e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25737430c8fbc84183a6d6f583ad63a80a4357a072956476fcaac033109b3e450e0613018834c1103a63342e798f3d9e37efc05a1d4d9b8c4a23ebf0729928516e509364266509f4f621b839c7b946361efc50548facd77ae926ebd94598baa0f4275fd639176f060e3ce6de811ce9d09;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb0b3faa4060e5bb95f4cbe5165707b4b0bfc214e2338c3b054d25b3b6d0e5c701de6ff680a23bc00ae72ef8b154cf245ff3c23fddb42a4dfc034ebc0c15060f434181c18168cdc39eb9798604b06dd24552428f2208fcb44573629558b52d15eef7a65e8adbcd20b7734f48294e81f14c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h455185b8b472cb57f43010311ec6c839ffaccc526406df4e899bcf30cc06e761c39f46470964f4f888db8c2f778b70995cec609cc8169951266a123305116563c7016361e114553f20945426d48541685918815264aefa9538ed5be0822b65e779377be26576b9bcc9c0c79d4c1d9b6cb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfaee09e3f15fefa47c778cc03ca6eb5d44d5f141af0d96dd07073e336fcb39b839411e42887d523974e46fdaaaa1e98bc1300bb411dc45ed5638b6e6ccb276746cf70d5f0f52cd108e0b811668e89bbeac17e7716dc59ad19f4541c4defe36726f6039616aeeea97a420bb61aa70d2099;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50beee74aff9456d4eac5138723efaed8c6b4d4e9bd2f86f0387e6be95ad31b39ca30fafe4f64495b20475be946dc8ec42be0d7f59395bb0e1ef9795b1732cc12362784166131c2758ee0bdc8ccf1f55eb71b751c71effbd3a8c7d3abdb11757ead4302f0f944ebd634d110dfcf8162e0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf9fb2677381505110e9647b0addea949230c334fc7f1fe98df631b4b7dcf058b191260939437c8a78281c947f49d84b97678108b7405ca797a6500d52e61d230b813550042f079df732b52ef6ec12d3accce017aaa72c527d97d696dcd4c0779d99d8282e9d362d4cbb4773dd6d14788d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7521ac261a88c7079ffa54cdd6895cbeb03c658189f5c2f0d8003fae494082c214f1d552ca5fa027af2e02ac21c928e19c8879e29487e837a652ce909f93220d7a004be90e993f4e69d77d90c4405697aa5759842d56c3f531e03c89052e98be67839cb6a3394ac7418e33c017899dca0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f6e170b47b907cb1e185a38fc55f605f565a7421a755be274bf21e052e69d483ad746af156a3c2377405110524d7000279c50a2005349e2fa440f450ac4a9c9b3d5123eaedb583839149a10477f5041ce592de560886ba382f30ad123b2672ddbd1296d2144b9d8581079e6495db2ad4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8295a2c61e4f50e9dd1fbc2e2b7e88f3d0ef2a77f46dacfc777a1f05245d89abef38381fce8ee9b0bc1b029293a91d112b896d47d1e9f16ce0acf30242e8f091568595d38c75f204eca8a6e5b971788923ef010aaaf297ff1f76797649b8fa13188b1c350d4dfa719d731e6db1e29c63f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h116058ea0e040431fbb92aca8b6a5343376cc6942ab25e157fde4d044973b6d65430439f9922c209e8c9c70a4dc16982b3c4449e4815e2bc1ae61f74b0d1c2c21ed8c2162616e7658694f59e1bcaa6b875bf7a57a7a148666b036079f1ecbfcdd95e9302f54dbec566b7533b25c07e340;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6127404475adb461476da925ed69e0c5d02bcd8a9b10cdcec404103e803df037e8cf0716c20e69a749921ff2fba5136fb2eeeed7ad26b692654588266962b333ec6f10057f159754cfcded7e3070ba889e91a93e712db5f98114aaa05d6ac4fb7da9b9b9fe816b72737151332d07393da;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7439d4e847ad693cb5543d53c0c2be301efa4ad9e4f7d2b4aced9e30eee8eac12a658556ef8becee32cb23513b6c7ba1417ceb124269f06f44c21f981c0a3eb93973234807de0bc4b31d63736d5dbecd6a7b56b4867d6086429a5563664c6ba67daa79a968b8bff8f987f8468c3eaccc6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48e9709b269a054337da56cebf12a71544c5f42fc998ce9815633dff949884b87ed375bbcea022e7f484ab4907d113bc6219d04dbe5f2d4c2ed5d6fed4511c504641db7c3cfc48264f051610557af35d7cea1c9d26c22d22dbc373928eb9b537f1ba9938a00fe77df908eb3b6b93dfa3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85d73c830b7615b6951129af4cebea934fa1e0065b3ec50cf7f9fe1539694a3cffdf8dce86ef63a6b43b1bdd83751cfab87273038333c0b0e51aa5b8f6d170c5365a71ddb0686aff5ae64afed253065c9733d5a865aaf51077a984bf26c1c6cee87908c16063b3cf4213336d2cc5a27c3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h85ade3a5d5a18d147d8ff0344e0bca6214f7ec430f23c61dc83f5b600e96e816b0bf3a51ed43f6eda5acb4cd2e6aa69b44e3dc32067bc4a506906a98b8d631fbdf959cd777bade5bd16262d2768da7aab7ccd41b3c301d913b7b05609059521bbe0d8b2f876c220e2fc985ffd6f071177;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h151ced6160efc11a19a148d238f32bd463e778a261622d5e38b293867f642f7f02dcbdde47d27a9848e440ffb87550c29c1df15745fdb1b1ccec64f659e87308cdd101cb7bb45e3be89a54db2c866578f1026c3ce963aa37054c187bd05ef40392536ecfef9481967f1b7c7d7dd5753cb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55023abd11ae9ec0a5fe6a43efff7a5c01f7eb9ecbf162df2d2d28f036aba8a997f70ce03ec625030df9f1c5e04d8f4ce94b65d1a0a65eacc892d7dac684ecffd710bd33f5aeb7b76ea90ce26de42febbdf6da13478e8400d702a78bf73278a7ada94378d093295158251d73560e19ee8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h94030665c5d609d7f9b587f7241d7f0a7485b0e722087cb1b44a38b180c53bd853290d420d4c0091d59a0ec09b3e63321a85442891b1b7cf640c4cd2d085c1e18fe433b881be4692425927bedf01ce83de5c15bae26e87e27d4620f14d2ccf477db53e0f2eedaf517fbfeabad45e32700;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbc73ed3a0a42aca9c399621b65a0cdbf4b5532a042c37549c19aecd9528a6819d8c9ecf7d2d45af1db5c9e2f4bd5985eafaecdcc4f96ac84685fa397065a5cb0e3f17c9afe7e21b67c9a3d9c487a08e96a873ccbaaf40c08e493f6dfb144f640dd13e71ff4e5ab51055ba7b8a5401db59;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h904ba9f2b72da4c066e904e7e9deb6b71c9ad0a928d06db1b1025fcd115024877daee1b13b0ed159791624040ce1f6cf1615e55359e73ba6671d6f681791f36945325a8330afa268b47200e5975579aabb124f508f4db1a6514fb92393dd89c6d45a42576a46eb56fadf7eb7020c67099;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h499ebfaeca8cfd9bade43a61f33c74ea24f31bafa9c38da00a4e21c40f95a70be7d26dafbb2ea9ccd599a7d34759e236c1a4e4394694f9b0fdf715f90d7cdc6a5fb1206b4301967ce229cf05dde40cdf94cafcbfee1d24b6da79f05690e3250dc5122020b2ffb5eae81fe96f0f174424b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h11f177c77bb05ff73f390d9f727dd14f840dbf4a5b8c50f159d04f40742027d2a835a4bf60cf9a62ea213b3092649c64907826730a4eb1a291b4657c4ada9c1bbf057431a0d931b1f23b184d9f8abb446492a9483c4f74dde7860d4e757447ed88b8058f49e89e17ff31e630cbd08ea8a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5ddeda9e99530360c59552285f02cc7239e0577c3d5f13e5f0de9c8ce7a9d9b94dc3515355fac96d0e73ac1510cbaa5bcbd8fbc3527968dbf9ac5f40ce8401dfdf7ea76b1701baf8f1958b745d1209990e91f88a867354b25dd412c1fc89c7b85538a6ac691e5b71eb42442bcd42f0d5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d13d18c0728849798d2a9b588501d5b050c5228e2353969b50fe37596985a7b9bc3d77d4f70f776e93d62b32558fa1f9a8bba8d848be7f428b54d6fb6159ba75c2eae5abd834821dc67e42c2ca1e3671a2d3034c45509870980d7857cd8a83856e8e4f6f4a32a3e7cb495621cbabafd8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h51254168152151215623cf4fe7f675d700338ed43628d75da4d116b3921597603e993543e31192fd4dd0e5b9627474b8706762672c1f2e863b99ee5a8f0986b97971ab310383436b7f13fae32d4011b6d7a8182e01309cf4dee142d845381ebbc8688079bc2ff3b60599faaa46deaca05;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4323e7d34b8bc8c790a1df7cd95ef0fdd26d72fbacf1e2152db3a1a01370900cfcea522e92ad5f77d3481b7aa2cdd434f67dc1a7cb603b8ddcd3c324122c547eb592f2c30836a5d2c4caccb5de6c65a5ebc863b61c314e0a97221530f3d3cb047b9de17f04df4d054f3f54226e833ace;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc84a2c0296e12bcd1bf9c0f6ff2c97b54807b9ec3a21bca21c43b19150eb1af67f53c602aa786c3ea0b92615dd807fbbc77a66aff51f5f88e055146cfd9973a1926c5dd559c056dae8781177f197ef4f8c43042d74637aadecf502c379a247d897aea08f991ac907d04822a18cedd63aa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h297a7dd27f23db81b28f67df977309985c6a2965b1fdd2665f315bfa9d5bd42fd1c834e3c5707ac8a5fb630550ba631b233957707859425ecd7a0cbc42d322e36b3ec709aa71dfe8b6a1716c8df4090330d589a1874d720e899d192cdf91813e990389f28b0e9c9475e09f20af87092e6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbe44f58405ed8d960b1b2fd5dcd49b289ce36f29027acc5626530646b56be028017d45543ee549a027fb361f9a514fdb16b59cd85b41e6d0106e6b0755d4ac04aa9cfc6cd5a4dcc7c2b0c10560a1cbf7b4b0bc15b5a22a23dd1ed8e240cf77251a90673994bb4005139d513ce43ab3e2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcea900f9d5f42b0b182a0916e2f9449576d4a0cbaa841a955bdf19a0b94a2f4d74d24d4c2ded836f63551c8cf6b96abdbf13c52d8c4361fd9b0a739213360fb06ee947faa6235388ff6c8cdae82ce20118167e07713a8efd7c87d1abbedd208e357cbf4b4f3b64a7e64d24ee1c12ec890;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5eecd8c9a80bb96be2ff29b88a848c5d4da81a1572767165ffcfc7e6ed9b74db11afca43240b9943ec70239b21df0fdfd07dbf2bd6009ccd5f6feb4cca9921738f4eafc96050bab3e0326d92d2887eb2ab956dbbba063ece7d33acef33bf3d005c1d5bf466ece64bdb55f90f8dfcc39cb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2eed1a2c957114750b23e4689a2d86e40c8acb3517bdd80a417b805957e28c389478a89adf4c5cba0cc1a254e11eae806a93996bcd3612fb19a0b9bbaf9ce626eb71ca08a933e493d991d87cee9da581a7e973ec0721b953b56fafadf9d4f033cc490735a40d67b07ac2715f4cf2ca7dd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h108ae6e31859f41f696ee8bd5a6b96284a56e56ca4c5733541384a152632e2787b8e8f6b1aa8d99304d4ea76029ae1bb1998a54c2687d6d6bdbea47a1fbcd2710aac624e4ebd7f0f2ecfb77973e37c5ac2c1f65caffda4fb5bb045d60b2aa98ccc3c0d182d3f5000cd6f69e3f2b1591fc;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9bcc5b18c4e886f32c94d36aed0b3fce0ac032e826c327f66275d99da41aada1026580fc8b17b4902926a02d4e8c366d8a33124f83223889eb66daa146a12b8db1a16aec886072e948820c973ced45e48d9e6b1c9cd84fdd5f168fd2e6f9e5daa98bde39f6380dad3db861cbda6058adb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdc5fa02854736d22db18f450c8bcd20837a96bb0f88a96cc2c52796f691622ac87c57c97d53e1f7f1fa655a4a540ddf3fdf7c946e1c3e02923f20ca3007b65bc47988c570d68d8c747806df60c37dffb5e2e612346947a3cba59ba3af3002e44c53b518c30e7aed03033db21ce8586d05;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1949e05838fa38eee540cbb1e61f9e540cc71841a8fbec142ca76fbbf6b15122484a8fceebd79365bca8f615c46695ba5533c769c21104dc742e817913a1a2986c9fbff1d1a6ce89aef117c0884d80fceffa40fffc9222464ac78c8f36141685dd74dbd8a35fa45177c820270757091b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h57bd41cda4bc969435b7dce2a40fd58d248c73793e621c3d6deeef18412d7932d244b247a1940c9750e1a74fbbaa3f6c473f5eebfe5830b20b90db627664e04a8b84d48ff12fbeb0de7b1bd0ab0c5b3da2f43e887d96420490193498dc9296bc74b7014bfd976e62ee979eb5011e0a3c4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f3d4d855280a98e16bfe2aca6e12d19aebcef0602ea856310bfb88dbba79b37800ce8096ea8dece7a21ef92e428aa4cf50f014106050edc99e651393907712db5343e4826b8ffc076c46ce9f0d15e7b409544899f8d6764d1c2cbcd7e30768f4bb03504b16e567d3422bee482b6e2c75;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50e43038c0b8551883d310f6c2871a1f8989195ddc6c206bbdbec6f06277e12976855a2eaefc4c56ccd1a47009f20f79cbcbae8c51c9a8a16eab6d216417844d847d283a59ad51787a97a22064293ee4a0c0374b35035043a56e2d2a632e2c0d5ad71306f1f9f70a1bc978d1ce6edff68;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3530bbe8e8bb4f0c53003548d540ea11105b478a1623a3d5b6c566e8ec03438dfd56d93b36f57cdb53b5fd94acd569d55ef41472e9ac8817564f9e4c8988708f6a26326f6d884e8736059565ea19983e7cd7330e87fca20869721e277ebe48812ed0c3cc759ef966ba4726f0597935d31;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb020ca5bfea23a4c644120333ba5f338d3b02b1caea3e02fdc23d1b787e8426ee9b6c825db2b7bd83b11b2b3613feef930c2a28090ab320c45f2d97e8bcce33852b4d5dd32e523cbc431cfeecf69c6bfb8e757d7ec65c258c3823e704ae644017c66cc6b1c387367ccb91515148c9f207;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24e81a762c42293c30ca2cb6351223bbb941c1447ecc494a1137e87ee8ea94545a0f657863dca545f26afb64c787d08ad428beb5b884d895784c12faa86029b1aec3fd16094279da969bc8f022a989dfbc4d4d847ebeec4a169d6ffc625f0b95db8bc1da102b3496e42fcbe8bf83bb296;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd4cd97a8bf9d4bc82e581e0fc2374d35984d37a396ad1423beff95888e260ae811699246398ebcfeb48dd3a2286f1a485d9c355bb2e40f74356e116d6dadda00cce26e0549c4105049bb53711378ff00a7b638206f8e69ba7d8000f44c358e61d2ddb0b96f34f28f31dd6452a46fbf765;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7760cf9a288ee48e4069deba6613b4ba9d66236ba139486787361f22e47f851ad029cdcaee12fc8c555b144d398796c0cf47f9e2ec8b32920ccdb056f6932bd284cd99f173617e8f3eb7a8ed280829d2bd0f795974a4fac75fe331effd220745285045205fc156f65be681b8dd15d1718;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9a3885cb9074c9616b241b542174ac3336d45d05c8def7b388c6681ec710752a18e17e426a17c3ca2512b10870a80504e01af6e533b97e5e87db0f03cfc4d8bb7f3a0fd853be1a588d743c492c820241073193b7a383f0de76326e70ffef454d956e485ed5aad85b8d3be5df45a2676e0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h563e2547524c3c921ecb59e51096cf50a3404a7000330795eab09fb667387dc4ba19876058fa85119d3c76211c33fe08f339f8a005642cbf79612d307956ffe0bed4774e07bd004c74744a46ecef3211b5f0d83f992282751fe59c9f7828ac8287771a0c0ab59d88025a49c0dac1c2c4d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25c0d39eff0373da80f7166a3561381aa5f9bffbfde8c35a0f0b39103834cb3154f6a20ad570a89e07f1c1cd9f0c2c7d6f2bb7fd0a7f78d15a9f6448dafcbe4234d82225183570da933d1c87b7ee8675c69662c82fea0f26c36c2b44bd793489ddd8d57834038fa09a85226aee0f2c561;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h83867f8e0245172462a1ba10ad4f8916ed664e47c1e17881aea2ada7b48b23cb82b9af46f836e910b0ef3e108b874db86e71c6f18b3257e225b5bdc1a6ac1b6740610653593213008a4bd045fd968cf5ee9648826886c8cf1be49a9ff3753612d061d30380480e64de852147f79b590d2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3c77f95778e582610b5bd361a46820b426b2bba7ec32c43df3da2e1dc05bc312f75df676dec5200f96c74a271d4368f0228aa36376771fb0bd0f60ccc68f26d4fc2b055d628581d5e4e788fbb3036ebecc628a832abf9e55fc12c42fa9b5f7c7c2160d0d27ac4be44dd2b06747a942acd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb901f1d8d16f0dab047451e6d0f74b6f50d78b57baecda99aa4873c735985f394b75c7717f31ab94ade7da78675ba4ac2a07013198c53da8edfc6e2032112a4b93f7a5dfaa6499628b6db184f5a947b5e431b45a59b70440e8f69822a947a2d47f9050dee22bce55fb764bb7add91935;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hab1633c90df8cce761af1eeb0e4a53f33c2feb00f8202922c6bb97a32e791d0a4e5510cf384006032569e79f4f6787548196f60ae5aa2f3eb9514157d77c9436fc44d324ce9cd611164f647f6588198f973f0171c9d79df283311c58e2c3266152457e52f44861609a45c9cc062c83b2b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b9ba33b7444020e46a66cff5ea7553a300ae6392019199a54c8e2946e4a1328290e7356504e23c89075990ce3fc275740aa51f1c18c82ea7bee93efdde37f2979841cee307a4fc448b5732310c07298edfc3e343d4606bc4d2100e0074d5f89f8921617a29c0659f91d7d7984822885b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcfbb1596164bba9a1a3a8983633162c9a56cf343b207a64541ca41f4d655097a047477331dbbc05d111428e00328d77f7afac95799e56330da3f8fa6eaafe0012cf11111502a97a7e8f00abab63835c976004976f8f5b318beab30f08625efeb06b8d66e39368243034140622ddb95217;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3011139fab9f4a16fd8828fbd7f58d9c5fb6d9d47c3997fe98c440eae03b47035f52accf825ebd99e9d94f97f55192f93fee555e31d5c9f01f709ebab835f86251553b4b5b2e1e137c9981abc9d02d5fda7b48b6e2f5e73df7441673fcc9fdcc189844497b4296b0a07bde2f828eb0dca;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdcef1d2f8d73320302bda838f487270c6cc2e823fbfc383951e9610f396d24200e563dee1d6bc042164b9557cbaf820b275be5bdf0743e69864c10a226668d7339482d9fff4b462783b2d8b22c2f22d4314f2c572a9f486872c41125ca0e0c87a3358e7967f3ac1e2e4f58cc957b2c306;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b5010c5e683ea07473a5bd294fd42cf0df96adac2cc1fceca26b2753c0136b39b6940efaf013fcfacb0581752cef13265561585405a863f62654247c8ecdb67eb940ef748fa0ccd3c78c0d2b0f612a6f54dae62c6f7321f1c9c9065c599b890fa1620629711673a6af3d7d651497f803;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5befdbfa885169417bfdb005ec43dbf476a48b465d40ddf1d22ed754b4932310679f2a2aad7a1c87924f14bc59e1c776e820e58b6663dc24256d3d9847c9243d8165c41990ad08117f073f89198ec132c53b474ed3bd38146e86136f5209725e605378f4546cc46fc42d0ad35e42ee7f0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7f289ac63df3b504aa2e876d6039b229c2c32c57d18166a61d2167d0a2cfae78e025405f6b4eada63400ec482210a1c1f3c476c7b4964b0ce42982d0c25830cde0521f476b40c2a7970f62a12de1fb061b3fdc3a5e87a128cc4c063cf6d4b98997b062e0b54802485d9e88bcc9197301f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb92b6af31f4697412ab362a8c3f7518c1bcc642e197967e4439f3edaadf425ab3e24d726baa3fbac62967ca1d20e898933d9b591fab0e3198fb75840a0dd550c7f9640da1ce31d9e061ec516a357967361cde2b5142ff2fefb30e8fedc14d4044032adb37affefa5314109e1040b172e4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1598cc7048aa5f741c25cd04eedcf35fc933f24e9575d988efa99ea97c01c76e6c0e008ffbc2a5cb6b4ab8551df7f0e104808ff4604c75c3c1910d745b1ae6f3bf4b318d64f07f2b178b08cecfde5cf3a36e1efa6cecae2a7b9789764de99edeb9ae76375c39482861e1ef07d32430da7;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h17f803b36bd53b4ff039b493fcb23d383057e45dab62cbbf9ed4b26b97418d3159f58c8f242d7ec8e8bd83275262e3fefc2cec99b1b253ada8a59024fd877ff28ac824e7860d781f46a902a40425a4b979403de2492e0ec1535ce477625c04e2be658c2adeae7c279bc9022abc9d4d740;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h13e100d0a45bd9d8b94e0d3959bb0aae153db51e08aefe625a26d3a5533f86c55a48b381aa8325e7d5f3492f42cb0d92f709d86e66e892d6baac1b284d7075924de4ccf0d3d0c992fbd7a0a44647348ee0384a040cf4796c88c61558b94a8155fa84bc1ed0c74eeae70bef01fa15d01db;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96e03bcf506c803ecc5c65823f68395a96da142ecc45edc14bc7075b1ab01b58534df74c088e8ea931f618af5d45a2a6074777fd5dada8b2dcd6b410dbfb93070f2693282d6c7779c9286c04dcb2439a9756549724781e41db7be42c9e12991a674e8a227d2530c14153fb237eebdfa24;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1d069572087cc2996d230cfa339ad24be7846dfa5140aa3c7bb6e0365d690ee97524f8f38c1c27ae9cd4d501103a1202841730d0b0b81ea17f9d0f397ac030bf18489b9eaa577138683472027ba6d94f469e8214b658f42ecbc676423e3a6f3eba4b951ca9160636866764ec7da543ae4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h92618daaf0cd6cae7bc286f26788b05a1b8c6f0ff5826d97fe25155c2e80be9f12cd31b56028d0b829fc01f2469f48363d4120bcff78c6e2ca44e2bd71ab5d052e1cee41d02a867c831070a6da2d8247fad63b38a683035f82c6f9b6607ee5d5002e86ef5da69cffc14134d9658899e13;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h944dc52c645e74ce34ea8b1a9df6891ea2d6a5873d3aacb687af30635f10b000777894b607a4afd312ca68b3af5ff7da91f6e2bbad88c8323a021944ee9974c28434812889362fdd362d257f50865989f7f878d9ea08142a55a2fa192b6df0e9783bb4a1a2ca4f1b7a719900f78f7345e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71ee3e4c38dc1b4a48899914fcf818c3f284d74e8521a96de77ba6ce8ad6f743645e4c25079a8aba4edcb938b69287d24d57bd445d86e886018cf8f150a5c5bb331e336bea65908157f0705050cbb66e166299c9d9bf658187066244c147656cdf5991c5753c2482a8df6af0b415c08c0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h2cfc1555071373133e8ab0836382a2e8e06d82d5f2213654d65d8ffca366f0f8a709afcb890c67b0697040ab930b152e633b74a30e819f77ec17218422900e7dcc65174ee2713d942a92f4f5356f37b78893b6d6566e964c862f848fce790452836cd6c0dd44e30c375097f3582e5e4b4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h76ab01195bc8b50aeabd69e25bf42bddb5f842f21c46c599dd76dec560f6e0a98ee52576ac1f34690b298b622f2f76b3a8d44063c6cab6f49871486a60063e762a1b6d05280fedc1f9be2c96bb6d7d3e919e1743c90d55e1017eca3a36cb2c472ea1c4b5844107ca84b0dbcf72e928e92;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6f96b283df15c7a32b7a6511c6f368ff1441875b3328466efd28fb26cc0e736816fff9056cfc6dad6933ffb910c8dc0ac43013484a8aea138453364f01ad02cf74b3a4642b1f54c93464febdd005ca21a4c206f1d09ffaa5a9a6451382fa9ab22e346fba8ee28bacf6468d6f6bb9d05cb;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h26d649bb5d842dff090f16b3b2140fe6b59688c54553bb92cb81cd7d5fe88019e0690851126f0c41ae588e45969762d6ca661e4ebad859df73b5ebedbf6ba25ac7f387b399c03fdb461296d81f3059d93252e282aaead4475d44c736d41bfd53512cf1e7f5193c47dc8e0e799d07ccc27;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8eaaf6dcf0e696556f413066db1166befaef29a8dec9d17ec3d67f1ee49f455fe98e261fe0e9814e3464e13bdac9a623d0a3fd8d8758edd5cc0ab261920ad65f396986b5952ae1257cb2f85a6124af26fa0717b97988733ca56338da26163e9bbb034d94a8a54d89f61bf42de87a787aa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hadeb33c7edfa673f57aeeb4ab70210e5b97543bd5301eaa0a622768b6382771710e248995b46f881097f9a88f7613c5df5ad6c23571b524be5a1cd0fca4a366188029b5e44b933f959888f4b06d9e763b8bc53060a59a8f59b10138093bae452817e63f5a0f5d51033dae7ac52e048f02;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3d6f8f2fbb4d8888739d2e0e1c2436410aa13b097c4f1efba1fc66052366e7ca44fe497d83377b40e035eb97f8ca2115fd1bbe0e2c20b5670570fb40629f3f5ec10a32323a595e808b986beb59769c7c78f36b957650ec9a48709da1416d8b3cda76ca6fbefb56393e01c057f27ba3c7a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h48aa3868a3c5fa98e44622d0519463cb2cda38d9cd7542db055679d628f9201f5c7b316dce0ccf55070e6744f257ae9a56a3cb6fd0b5f99b8e1f0363d88b83b2fbabb5e22edcc47651c893733f308055d5ab5690ae8c74dd7313dedcbc23248e47a223e4db985e7fd20f9aac77de4abec;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47725b6f09019b16a3087146566ad4fb49cf87668627a9b8394ab1bf66d0496e495c5081b9a24678b8a6fa66fc30bf46c958acdb0d9e85133ae415b2d516ce4d716f1c9b299dbd9c49b68b3c9ab3acab636df37d68ad7ba7ffdcc7a4669b893910258f1ff9f62a99b881135dd58eeba81;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h55112dc99f7f1f99aaadafd67933d143cc28b871becac34c0c8f06c2d7dd0ba17c1cb02f7ebe2ad817c2b09bafcf4d5abb57fabee84b5c8b589c8e81ef39246918e7e49f4579c73385862cb0148e68d00593da1598bccfaf1740727f06da6ec33ab7a2bb19f6a7f10f92b284acbee9400;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h54a78185fc85a967dc6b233b55b08f97075f33071ee1790b3300f84bbea286c1047bd351deafb0437bd4e2d5d0f77b104019158801663f0a71e70d74d02e8c596771c9e49d80c8558ff67d6e393a32d8e794dd1e18b3e52975d56e05531785c45a5de70e8ade53db7ed1a95b61168e40b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h842a6bd7fdab89aa0816cfb083e3fbe52bbf84d49375429b7dd26e0fa249ac1811478adbd5d84d09a6abeedb85056bc12ac720198ed2db6e17c069fa1a093397d6120353bc20040844d04ffe2e232d89da9eccaaa2b70a1d31c8b692d38bdc0732c0b0547a406021b021c458ba6bb2941;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7dce7822836f5a9ca13338dbc46c2b2044a3bed929c82696396f3bb22e53e642b1fb86f09b1bc93c3cd443173ed3bcc175e100f493c03653a91969c5d5a7bf3950b8f5cf2b7dff538264fcd9a20a8a5d6ec19772b3db706e2ea6f45321a5b37530012c7b5eed68c2eed022691b6645850;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbb35b2015bb8d199999e6a6f23ef30143bdfdf6be949eabcf81c239a27483dd56c1ec343f29d09154945ce70e77f58c40c4df907422bd5c41154ef90e5f2aa7373ad8a61da662870f675dabf63649e259b06e18d90092510dbccb3335ad1a4fe8e43cf873b1ba8cba2f29db95fcdf4b15;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h31972ed0a503b127fabda8ba33fef2169451959b20695f03edeaf369711a7a376cad5206daf4f22840b68bb0a1acd0a34f7349cb851c8127d5e227edfc49a53580e14d36be90aa56fad186a7ca4b7d1cb3906320e586489bedafcea382e86c15c1d3dae88a6ed7eabbec55dbba1d6571c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24aba46eb9839203021d17622faa5975623da26da282739b1f6f589a719e30cf1c0d6ccac0100d6134612f077b8f009275bccceab1c89fa0930824d63902d2ce0190beaa703eba2f8cac7e783585d7e77d2d611e4b2e7e52f284d70d0a48cb711aa6f4e2a75e2024f990f4a057991969e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66b1536c7e3cae55027d9f57cef72f2313ec081c0eed6d5fbde42553e358f45ee24f3a8c9c772ff65972dec5bb8e233804f7de0d45f5e7f3e3b818ef1aed88b533efb2e2b55254b8dbc59ee7ddc10f743943b96894c1320f9d2fc7949a181c329420875ff8b21176c8a7685f0cd298117;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h645723eb1542a714302f80c7b0cc7f3c595c85df1b0343ce4e61ca048c99eb131762db9895e0b00b00aa324e10663982d6fecebfe3a255d5b10601230f81808e5f66327f257cd44febde864b5ee3f7f8bc7e186c2d9d4faa84550c4ca4a8b6843632d0956600e73ac3597a18311e8a14b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8d1e2e18948ab454002a7aa1f4a654b5f44ec17945e0559916dde9ecbe166e03bcdeac55de98533f35490686395ace4a62dad3e7c975ffd379ce9481fee1c6ea1c13b6600d9ad4c462ff607c5b24d2e83a0f009575ca19727c8ff27949079f99ded89ef1bf18281af7f97de9362169e20;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h61ed7937da6dbd05ca6de0e19d7dc6d614084dcda48b14c340f3b4247a6bd74f3a5b7320ab06ae5186eb2b4b1e50be726a9dce76ea066dd80b7c7826a2aaaa60b63af02394923066be11e3bee40b518f5a37c27dc304d7166eea85039d242b6af872f0b6260a3785dbe1b89fff08d26e0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h77c79850a8aaa3bc151b956cff65762fc4ed599c19c959310e36a5d21c1af06ca80387bd049d1770dc19b4a1d004adb1fb33570d302e20dad28e3a2c9d787151f73c0cd31153754a5ec7cd69880d2cc805d3ac0e06958f3450642bb183cb4c0923d2f59d2a5a3b531ec88230f7deebfa8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9c04c589b955060f07d44620f54d02a9204ec53ef896edecd899f2ed55b9d17b9b7843efd97bf321532e4d10ebac48e2e000a6438c11b51c217e8b9432a2bca2e7acb8a92360c7a25703f8ad7ac1cd1d9200f95673992ba4324739509911a291f877e1be62bcc0806b2f11a3225aad801;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha5250d5f0dcd21443209d7f2a03e18af729cb873406c56a88cc34d2973660ca660ce533cab46b270004dd2ebe1814b8663a87545b4a04f40eedf61cb49408364fce336b28976ef7cc3376a1370fc5a893466ce4df7815e4b27f80736b9a23a80c3dd8f50ded4b8e29e52b18ab69a63c45;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h25cfcd933204e0291cce8959491ba136eaeeea5852f1271d4db8a84e7070ae3a06add45c93c5413932fae9b2db59d11e2787df8306a0038f57d3ee47e5b690f73d04c4a59e515aad59ac0f3e8bd3c68ed6ae6b97ddabfecc2b39bd2539cfc92e462b6bfa3c1a1989312029d9e485d3636;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf02b4e3bd8e21dd269737fb8da4cb884920ce9a4cfbe2b7f65a2fc66b3a7006c3dea6fe8508f3f89a581949cdc036907e826c92e73b0142e80711317e4ad855f11cb0d0f1b576266a89768e8224b566664ca45fcd4b6b75a892c00f75631a59abaff525a8858f02bf2ee4fd15d0089e57;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he112c37f2390c491e97ae372d58d22d13171b7fee0c4f52283d8bd96faeaf0a162ef93cab64c778bd0af30ccec1ce4b3b891813d62a4983484c6afe0dfd924d7b3aedc58d45f64b9c077c65a4dffb86fa594b61a2db14c52e2a846449986154f2ba6d8ff81b6a43245155a2955e03a1f9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5b385d6130fe58da37a773dbdffa8d1a3bbb1e62fb09c622c9625b4a3820fa458bbb99d4eed52e2524c0122af243c770fd04ba9b4050125be60a3302c02d0b4e44b134756a68adf17b0607d7b618dae84c7b73186ee41e195d964e2b5d589a2e9a2a94ebe5ee7ec2e8a74bcc3e092fa80;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5c85aea1e2feb2b970d1f605e9fe7446ab7fc21ee38726312c64d7945ff1dea47c65f09d87286e2e62ca1bcb63ce914618f122e55d81d57a13ea14cf84a32c13972cb87d12eb55ac240d88db3ad01b78ccdfbebd5f4d1c16eb707a32d4aa27fca72e8370f0fa79748de84f18b61dc7f4a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h62785a3199b350020ec113763a9d6085abfe7e1857401ae51ad09bd99c289da6c1ccbb1159da81b14ea9db09c2eb20122bc469a75b82cad35b8f4e3099803377d473c66914833b7526ee792eb5087181a4aea45c9ac6234abf85c210bb908501caf74838f36fa3777abd5cc1dac1f5980;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he164a45827b350175b5272358bd73b19a9cb60f4d848bfd3e80754688943fa97e8bb616642df31e6599c45447abdb1b1da5c8f9d4481073fafe3f8a12a201c5039e43afed5494dc6e8b8fa31394ea17f33a190ad8ea97de4db9b7003def600d70d94f671e004838813bd3ccb9ad906f8e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7378314dfe6e8de126f882ed8bfc77e3bd53c0d2f7d9b0065823e25e0fbffb14a61f609abe7ea2fd2aa3b8c99ba499135ba68c4b5383e5bc0cc6d56fdcf9e1a928298bf56da2208ed7c1bfa2e143a3c60de8ede0c811740409dea8bfffabd3b46039a63a199b222bb784e06300cc1648d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb9a982a99084fbd5914b384f87fbe4a91076a5e1cffe4c0856afe5777d991d8fedcdf313797779fa23b55ccb1321a3566d02751f474867e675f1baad4820d0533fe33ad6cbe60a5e0b21fd84bfa29dffee18122d218fa269bc4207e1546d0e3a4434712ccd1b0bd4069f3c4f04d95266;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd3ad9254d584a60db132d1dcd6a3d9ebbdd018989058f3c5c16e6f5d50d070baefe89584a2b253202ea6f5a7cc06535becb1f6532c90758b63f7257c1ad5266aea3d16293f48c4ae51b0bbbe66d22f7ec04e3acc856e66e5e3c6370903ed0664252ceac7ed415df60e770e6fdfc58667f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h44cb88a5b41e1505d06b42e09b1346d1a7bb65a3d40fc34d4a8f6dbce0b4ccbb45efa9d9c7a7d2fb528221655f76e516c72ded32f196f219cd29b7c15720abb90ba0fe0aec16892e13086bb341cc47cf0584757431409f3bbc3c0643443f53d28567bbc06fcf4c021a332ea5599372eaa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h144602043b2b934626d1c143d0231e02b05817cb9da99dc6fb7783420a37ed4f5341ec58f7dbc97fb1eb71acb0b17d8dbf566859bac3d15bff3e647e707e741d60e15615f777a571e47de895a2153b03aceee508e3577fcee4f5ff89d994787f9e6ef5d496d1477185c94caaba50f602f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5e3bf14c1540a179d4ee5f3d84f6879d53d803577f60f637e6e749a741f82519a71bb478d398bfbd2f242acefc07921b0226b39a38335977d56e7a39f5dc28b21f2b44f916def418706d26e17229a63e9ba79812540777c3bd56619c8a2aabb415d69b12c6349e27e1572883506353815;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7678b672d4d863082dc71402602116cdd9d60af02ef0ecfb061e6c079387f50e9a96a358b05ba1a17dc06ed1e0f56b2e48387a55338adf0d2a6b085f1a6e6af8ba572acb460d8b59734016e7e08134c9ee96b6ea89e3a9ebffc62c07500c7c155e76446fc0a82f2ccadee8c582e4b2451;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h63a6b2bf1f34df50531b3038c36b9a8b8f4ca8289d93e3978f42f57fb34d8866195aef43d830ae2d0d2ad2b71f0db4de028d47dfe596b24f9e9b9972a451d1df0fe022358a28155dea0237881ca0bd75c3dbbff789875f09ab94da68150eae7ab6dfcaab25ca48952d94965cafb27184c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h90fdb5de752e71a5805fd10f5538f54a8b3f713f76f2b80b5f0affbaa0e8b653aed9d7343f8f914a3a405708655fb75942aabf349ababdd934a74a9d4424a849b874dcd0139c2e10445dc983c5a9b8f73432073400a9aae583353d20d82ee25ff0fe5157169a3821a34f3621d34c6ce17;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h402429cf3f54eb7457b8301c3f3fdab5b1fc2bd1ec5d216161958d99ab1d84de33925ea7996a0865e965bad46197defb801fad2257b9a5065df471962394239bd45a9951d3d86bec75d09a67bcac64dce7d9751b4f85c53853f7277c2cf6f274bdcbfaa284b7dd14e5e07e5bd4788d50;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4d41822faf0b74bf28ae76e803d21a72760789279797c9c169279dd405ccf7aa926d4beb2e8a599f9ac7fbd8d31b36b03f9ffa8b79187781b4775da45eddf703d7d4e3db9f33ebb69fca1a6ddc8b1824917e9cc9ce8f8a7ab1a4080c152cd8516b988beff971d31d8d8e426a7b303e629;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha4c08e3e6ea61e815a884f7218d2edbadeb459b8031e5d1078c87cf2772b5a1412939cdf46860fce532bde62b1b7c9c76f33662cb3340dc83edf1a7cd95250782225c9dfd292538f030a7dd3943bb112a1c6cab969373eb3f26c9d1717e7f9a62531af27af0ac660c18e4118e227035f0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h954e0d74e196b4c973b5b2424ea8bc63d424ac656f1c68a8c514ede58b04ed60c12c3a652b0d6bae6c05207ca6d1a526c8438c99cfe0271567af3d05642ea8175f7a9a35e40c2633538498f63219dbc416c3bea009e67ad2296a87d526bb81355052812cb236a96a0952f2f85e2ebd434;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h69a0199b75731aeebea56271ffcff5cc37e2ea2cb501ba9d8d18dcf25afc6cca58fd15747c214b2eacd234eb5f6d84ca9a08ab6ba0230b2f99a2db4ba3a3c94ed70dfdaf66c77528ec9bb6d22467e43d0e19fc3db6c9791828dea4d70e9d981ef737a7770ff6335a7233b531d23c9a393;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h458cd1fefbe4e5b31a32f98f472c843add67a013d99925160c4acc3376979630b15b68cc79477344f9d271e30fa858db4d6100bdbac717cf2d5f425e3edeaeecf1cde9851fc65d95d19bf8670fa4ea50174a533c4f41988000b084477d70b54650a41f3ab13b14081ada7a8dec5ca8364;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4a982699c23405f21a8b4514f8d6ea02dc477cd73a22f15157bf14c8d36d0675ca13e27657f88d2e805bc22fcc34e22e075dac593d32de1c270f5ee5a9d529508fc3394194c99ba4d2d43b26be1262a49fc75fba05a98e20c65bf69a3934257ed47882f102e1e23f6a2c18d3d2085df11;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h365c32d2af085e17816b540d15663b6f064d5b5d8703cd03e230089095bca9659f08681191b0ecc971c9408cd1446cb1b7d50d491bf8905de276047f2d604f9218eeb363e8db351cc5558dc15d609050226b561d9c278e7a8aaade7d739c177943c215c5f6de858b3d56ab0dde0bea15;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc219ba3923e459d81c627d7e9cb25813b027e56ab428cb4192f92bf39443faf9b74dc3e71ce5aa4ffd824f3fe9b6d07d509cd6ee402411e74bec9a1bd54dc66b49faa69c7d41830a17e5032e71f94239219bc5ec10b4758a005effef025f14554268d6a94fd81ae85f2bc3a0a9a95515d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1dbc8ba1a4d97fdef3f6a50e271471d8ea3613065278e9200ca74dec806716b0f3cbc8ac1d3fa37c76642e899b9f9dd981fcc473931ca751b7c8ce73e50bfc63c45f0811214731ccde4673d28f36b3c1af3e192d760181aa7df0d7336d0dd73c21528d1bc2421907ef4d8c57fc6a883a1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe79a4b2c1fc5522a6bd348432f585aac7ef91d4df111e2433ee1d627657e93e7e6345d239a0d0fd9d669f48031db2d9681dd0213161535d516b2201d77e3346a432a2c9501fbca4fe496d6b92e6e3df712863c1d8e24fc440b75ff5d2b62fb9596ce8ec4b21770c64bad41446f0faaba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hf40a34ee72baffe9c178b451bbd31aebd5f8af021f7744a1a41cffab1fbc74e199e72d382308fa49629e67ae94cbd3bd8dedf709048ba3579dc4ca0302524cc77a04141e3f39ad3a9661bdfae7f60037f10e9afbe72586a61c400df448b5cc086b433b34b4c967b236f4093dfe3b7f3a9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28c0d182e7037ce12c4524b960746d11de4f273e4ba3b86cd08aabba68901c249fb71c3a20844505bbb113e306069f09c97f9dc3f9d87e539f35234af3352600893c4c6063dc46969001575ab1381234dea1a12c3437a5c4528a18201525369f98cd1144e5ce3e5ecd7ff92f89bff5f58;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1f7f84799ca724f565cf519ffd095c1f0850e883260e2af871c003d72548275e5d26a8d92fb63cd3bd5acb1a0692b08b5792e3b29d3260e21fa1a45b4e61b3457db6105a41bf4191f39139a972a4234d1bc68977855acbd55fe71adfaefea3390edd8c456e5c8d7c9761f1adcc61cd08f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f014734be58cbdedd8ed1cd04d4aaae788eab73ba1f9a3894c96cee61d2112d085b1fcb9d37a4b49adf5cdd4fda429ff830330d7503f485c367e60937391fdd2b6b6c01f82120e4426cf10b2623eab11054a9edfc7d57258d30d8677bd23d990d7495840140471fa72d58375a99d45e4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h118833d950d06d8ace05c8adbb097a6dcc8fd5d9acae4ecf1e7d0b7015e1a0a653fa52a82523f2a18a95a427ff4a6126484c3dca934e832ea486694996c7fa8a95f7462cf777a5b64e4cd177e92319476273f854ff687e1aff5749c80884cc82628f6816f8ba5df6ca800f4718ab530aa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h150cb2be1445b66ca63b9af7fc42a7c77044a8a927b162ce8e087d06918c1fb2ecfafbf0846d60fb3c889b998593b87ba8bf7843b1c075de750bb2ce237637a329a25560362fc237a1dd37127cfa4ea4ef180b9ca34c61399c3371a5e3412c47e8297e3934b475880b23014593a259966;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ab64c14e2bbe9a29047b10c68d4a127c79518057dc5a715343cd33e06c52cedc0547eb9780b99c79c4c3123a9f29b5e7e910178e8bf45e67201c3eb6ceaf7df8cd353d9a77a8e6cd386e2278c84bac4df6147727b4fa8fa27a92ca2e15778936feabbfc0040da1b50ab5454ecf9432da;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'had9843ac9ae1fb4baf20f0e9e171fede1fcdda761b9891be4aec12a1d215c389f564d80139e338e89646635b0c9a655649516d159fcb5255f0b02d852a18edff85f50fcf881e393a7f7c1f536adcc6c4d248dca1c274d963d79dd3dfc9beed8f42bbacae424f1d09046dc8d997311c35e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hac22b35cbd92c6bcb2aaa1eb11d6efc6d049f18693a43a89e72f4fe87055f37f6e792f9f7357c31f54214d1e363c2aa80b15c393f9f6045141f1dd05561a0c997bf1ddee35424d354ac62a06ca35050c43820764053db111b9294c403b5ac3cf352753277db1915fb4ca1173d57f7ce39;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9ce1dd010d2fb4637a44e1b96ad7202bf31d0b17e918a47b194cc861a77429dc2e79277e6423ec130cdd1c2e411ff3e3d74f6ba55180b6c08bd86122ba8ac94bd33b30eecb007dbab89fb5128944b0e58cc828202f7f00d5068ebb60439f3d570df7b03ac443390e5ce1ff0415129a609;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h71c8fda9d76d4c8e8e142860d4d4a4e2f0481003f0aeb80ce2c2f89227b1588504e582c6b05561ac1d8acc7a587714c31589dc57c972a74a0facb51b70fc3f1304955996d05229e14db5ecda3d99c28f6839ea6010c05725607cb1bf0650aa65bafa0a885966aff42629752c7bb466813;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfd4a4a6bcd17a9ff370158dab6e6f5db209a0028411adfce930c05060887f3c9d2d0d55b4a9a3efa71f938dea9403cb6526f3037db95de71ed1d70eb16d76b0d2e3098c0478eb9e67fcc57aff852b00953b453f241ae9ee91c579efbd55bf37f1fed8beb42e8c99dcbee392d3bf02c7d6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h47d39d87695d7823a037f4caa5312dcc837460f0cba334e1b050058c8b1eddae4823f55c864159c4739ffbe7576b843a63fdc4106120ec4b57ee001586b7cfeb4b266c8cf9ab12524aeacdc41d4c63bd715532a38a85f13bc9bbff069f619b14b4684d07498bc78ba06c6330ee79add2a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hffad869845bd92344766e751df97883c0cbcb19c4a6f01d491c29bccaf88510f43b4e25027409895f94de921063aa901b8e7946475f0eaa5a209c42df006d543076f1064f4bdb35ae1d465bab5e0dc75e9eca7ab8e1862f7aecc76ef31ef53de3775be66705b43050a44ef852a1d9b19c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8784fcb2e4b2c955b1bf70e9d82d66fd1b3aa01d84055f8e1111c949a18820127f763a1901c89fd3539d21ff5753639535067a984916c391c219d94a97f28eadb907d84d3f2c6704a0f6582cefdd2997306e895ff064c05fd46208a99012e315a3e88e6bd26e74036ef81c95ad8a6d64a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc30dd360b83c0422a690d2c5f24f017357a71c97f88da9d0c2fe685e0b467b504b8900c2e07f0316726d504fb4b39f273aa3d7d6d56b5971e5d2671947476a718e2927a6bcf7ac5f33aae43bcc49231688dd29a997bb35f63354297e9103a506ac200fab45a732325a8d3f700418ba8e4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha7d710de960db7b98420c88931398128dda65c7ba1d5e4eafc903abc52e0699290d8df10d25d54ad290e2b890d405dab2d5d73a26213744fcb26d5b79897b369397bb498e75064b5d5a5c964d5d30fc79ec177c1fd53e1045f4af365dba0450195741edfddfa995d5caae012803453fba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50bc86aaa76ac76cb16f4f71d35b3ab561c49169f9353a3e9b4bf63b327fada51bd4aa620440fdab40664e4f57192520654f53a894c13bdd34de6352e41c92da48d80d2c98600eda593fd95fca0a1c170f5bb8fc8b2578eb144f54f2b23b1522bdff577c4af4ef2155d51c264d0a2c300;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4ad006bbe2eef412a1cbc06e85bdcdfeb6152c5117eadb05fd82aebe709e5bd064bdd5c464dd8c70b00af4a612830ab3c94ba84be7728405abd6aff0efe816e27f2ba873bf3e21b3078114dc203707330bc53feb5b97c976fe4420f834ef1f1c0eb4cd05f47eaaee438b2b0253047410c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h954558521c5f631fbc8645ebf8f2b186bd822c3a8ef4495c36588e199c652c5e203297015fb10309519779ef6066e1b740089f8c9862b21720145630ffaaa0d91c7910bc5ebdeeb16d11bf19d6ef82997db8a41e8bb3c1473f6f84c93f6acfb5c9fd29f5103685029286780d34b92af6f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hefa1436425278f417953ea49363779d81ffb4390fc832cd154d6161931fcc00b98e6ae60c00337b698d3ccf85b6773b30c63eecb86eeb05183de6b7ae17cf2f1483858e9cc6239dee30f5be95cc355dbe8a219f43ad0bc15938e2be4ca514f5d2efc1d820d3a9b434a661f8666d7b061a;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha73845f53be2f3f2d08d55e99c00b08cd9b0000b67d0ed3b7865aed824bd492c705b79a87c656fb7a9f20838f66270c29bb00d490cdc6d2fed7ded17b1469a28edb17d6b596715e727e61e955c531420593eec688ca2a412afb3928fc5b11d520bd3733e6053a2aadd08c82171aebecb9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h247f281ce196508bec480c3f269731875ad5cb54fed7671b8ba075a78698329bf65f4ece37b82932c8fc5e3528970bdd5aa3d7987e9f98853627e0786ade44d4aa2dd793b4a7c820c3cae274b526402c820863c84a5b8e4da6a8f188c10fef7827c2a4bd18f335d6447d45c67a8403c22;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h513075e5d72be06a98c3e1b274d659a5f1cba7a476267da2282ec58fd8e4613a200d16e2e149254b7221710fc82c1f4af535fc9cce54aa16a34f23fede6ee5d7c2528ce61652cca7ad4615522c0832915c75a16e696b321b841924e23f2ad06220f13173f26abb86d55e78c723b6a04e5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h484bc09f1ac8fc4da324db6eeadce3254e0388a1b737181f7e242d440f2ca9df3dfa03c5d37153592d01f0c1386b342b8d08408ce4a8b25a4139904156a93443ef7e7dd0ddd7d2ae28297d001e7cc593f7c0de797fc8b3cbf12d1ffb109f4f17d439354703fb780757dcf7819b075af8c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h64ec2db751dba59d92d7c0901fcd1575051027c133ad90a5037aa207920d435a6d3fcd28db7ef7f96ccc0ccdfd750b87d002fd27602dce5bef2dd62eb534f53ae276d64d3fd4cf06b8209ec1d2efa9bf7a75653d5745e11b51c73208599b5d0298347ee4b2450a07855eecf40eb33a36d;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1e7350b18fcb427e1a95783f917765db4820bc6cfc684c04a6715f7e5decb2638fd63d03268729ad31e74aa724059322c5d6c4eeac129f6ed44f98df891bda31a3af6ce08f0e80156d1b3fde277634b34d2a69f788c17996075768b0b5981c4b82a68c1a1abea2c46089e040cca87f4a9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h67d1a5a96e9cfbe3d7777dfbdb784ae3cd6da38f818455b2a7214d6e64a58a5b0cbeb8156000cdbfc9c873656b3b1081680c9f2a2ce410bb179bbc116d6155cc2cb37898e8d3382e2b280fd1ad3c3a4526105cb6e5a7aaea12079a1be52280499fcc062a6ca71791584404cddfc7be23b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5162a840f412fb990897241722eb858ae5237759c2c05c53f5b43c1325734541c66e9083906232db3c1f4cdb48babec67c25a0145301d3f006431e4ae3f571ad8671391dffcf8eebb4c4234cc50405e5eb0cdc3fdaf0f50e63ddd07ea7130237cbbfb85c1349d9662872d790e7f5dcdcd;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hb93e7a7748d784d27ce24d2b0c8bf97fc6cbde0fcdec98cd08416dabfe156edf78c7ee1346d1a09803dc3bee508a841783f6bfc9a3a33543bf3f9fa5edc46e6f74c6b967420636e7e5d2b0169fc6ded453d90e56c6563e9d96d4c976c4db30764476d74eeb6bbd242961019498d68c9d6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5dfce06ad19f48121e06a34bbf08438098eaa2dae744b79bb68958f969e2662ab6595f63f8870960883b0fdda84d9b38ecb958df8b54d9edfbb742e236940ee1bb012e6a6a557f6f3b7d9382069c414cfbc1ad5b9b128bdae6e5fcc0ac474e6fba97befe5fb126d3baff08ce87c7cd9c;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h49bb1499cd65da213d80858a42c83fa90113b21a1493468f5202d9f5746a4d813fc8dc1605caffbb26da478fff927637ea14b0874b7184cba511f3308feb6b6ca85c071102f178b4a403870c1b47efcdc26153bb889adfa22c72209b64d8977ad2b33e6d9147360992646863756580057;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1cbea575fce69aa858d7824815b630b5784bdcf59995ea15674c3d4c0f5642c1026e6abd2dd0acf194b678b1d28bf27d898097f47c543188efafd575af4daa6833e2a9954441a888929d53fde500acfdca8675bcab31f611a780c54d648e3fefbca7dcc33e1882895eea55dc37a417a8f;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he1ab60ba2b8da285247ce2c6075bf3968eaa3c2503a5ba6100140eff48056935a1426127a4c526a0721810e3ec847837cfcaf524a7cc25f0b57dc19f11b1a0afa630bd71c5a3f404911ff4f5dbb09fbce85c9512ae739ae4561885d789b15264b5941ff5023ded71f66de4023255b1ed1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h82643e9fe79ac14743013bbcf13c5e6255a427590b2196c36b59eb0f9c469f2c83fd21ee28be6d7748df7cf8c8b68e071771d0456b3884d064831ebe27a1fe8602586f5b1e03f09204e20e0a724184b77390d394a6d7acbc36daff37a0604fc05a232d06f33048a9e808ed2532d68f0b5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9940c6a9660d0f91ab78f955669688d1e5eda848e917433498b64885d5842832ef781ce950ed8cc7b25c6654dc42eabe1132a59e44201bf1acb01621bc04f1e52f78e874998b63838d81dc0fc6a97633f2df733ab3e41ce5b76e9409cbae4727cb3e43248f2c679d8f8854368e01ce9aa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h46c5cfcac3b49102b77dd7ba8497129d5f9e8ed9e2926b738b96066686c4cad8cc8582d7651a12b27c9dce8583f3d2ec443c2fd759a8a4d35b56458ffe5cc6d1e7ecc59e60732fba38826a1affd78c3d546c82d91fd109d1f5aa6514fa2ba035163ef5d75af1b5242be0f696dd25d49ac;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfe6ecc7464d4140f601a3d135e6519ff1c6b6e9ab0b1b0eeef62a6fa3d533e545694694b1786a2436c0052d3de799f26555cef8c5c88b0d69f53a4adf8d37a6b2dcde80b476335c94190d52d606725abd4ee90892c06ba2353fed9e67db93cd10e8cf0a495ec047da150ae97d37e085aa;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f30359c54e3da999d80f5c1dabf1ca98dee41ba79ed841c5dcbd764ca539bcb2f226155b7b8307dc1dcfcfbdf2ba10dc3ff640ac95a9571037a0dbadd85a5ba8abe0e57686ddd1c7e145fe4b2309599879a50ffe62e7316258187cbbf196d7d6a558ea11be1739f78790d360cfb7f7ab;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hbdfc76d6b5e9b517752abc518c4016aaf6ad75197c2ca2c3b3ea10f865c9bec03ef8ad8437e9e34157f70982c53bfae3b8b9fab416b73240dc096f4ab0486f650016089938a71a3e0646f12e8ac78e238e0d3ab07e1d44b11e0cceb61f4634b06e7bf0506b5974ea3a3fabe12846ab26b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h901f7da34d9581f70ca6809e8d31b8780fe526be48e650669f068d00b023234d9b4f49314a17f814ed114d1c6dd0d4815e274c2e265339169912b0843a0caf33901997b1e26f587310d62dcdca24163eda1e05386e873bc33a6f7e9fc3b56c591bd5e143aed01044eac22c1c2335b64a6;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97cbbe5c3a5f02be110f8fa48c440b2ea02dbacdfe440542cd905ee4d21211ee7ccea3b38d3b2e4a8a9af10b08426c0da6da75ec598dbad38ccdb92ec8c0fe7e6837d82ae2686538868c3824ff18933b4cb043109e8536765321ddc4139a0fcbd183cc42dc9a4192ad34626df4ac6b8ef;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h24baa7d1801921c4fbba79104cbcceee765e480679062cb25c7267d97260d0364ed9e9aec4e38adaa14ad0d287c0f5b59168d6c8d43e7268e9210f52bf15bc996feabc18deb70e124b53a9d2f050c5ed2da3ee57c7ed76ffe2f82381cd11a6d6853eeb8080c520b9d6d534523677b43b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha202a838ee2c41c0b13b050d42b6cb8de1ea5f3279d0565b405c37ec1d80cc1568ea79d651f7caa5c82603f0ed200211539995ef619e77217f4c8e6ba6971867528a851a8ef306bcf3a9f4b9bff6f88530244a642ee87e83ec7c1af552d0844605d8ee20ace7936cbfda57101b3645515;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h97f814fde7eb8108307f4ac56cec19e0fbea609bc5bf363a8c9db51bfacf134316df73dfe580f8c95de538c42572a9fa62da1347337dc076ff9c391111160f381d7c24a262da65758ec9c9ca7d39908f93c546ea39431b3e42bd10bb86ccc58a323663c901973142d5bb4531a8868428b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h578894b6f6c45ec473bed3c29abd25efefe3210cb1c96997c6e295d6247fb5227a8bd663f48f9fd08f7b4e0990041d59cea6ffc3a14af90ee2c2f8b2bb80ce6eae53cd8d646b607400b04f1d070fde2af6e2b425e3702413d309f49dedd6fc08ed96623bccdc32a90262a98f12d2e2c40;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h32687aa0ae8f9b2d1e0278c5e1773b2486002b689ccec38cca218a353cdff04ffd30b62d123c694bfba69b06895c9a07658c8380ff30a1da3f2d4e122e87a61b8ae7913e4b7e485a5a2f8cf372be8f5ec44aa8d5f04108a0f4ede325f488c0861730db29d9a87a0157483d00137dea7c9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he44bd7635219c0960edd768e81f1a23a0993a82ad86ccd4b26465de3b90d3c0a8d34109ef478078189a1ba734bbe58c8a7175a4b67058a5ce2a39afa685c9144f920b0938589c9b7efa934fe051212afae404eafb5b2e67a096296b835d92ca9c0b6f16b77f210bec4012a7eae6749d47;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'he7c92babc0e779729ce47287ae3febabac1567fc3e558909b8e20050cca74bae3688a7a00b9de69cc1a18bb8f4c765e64efc0f6a60f2806f1c7d5ec9fe87d84e526a4b250733927fe8d1ce500eadd6b59fabf386e2c57f1a0a7082b6a57e452449dba52de59f4e4c52c4812b07ae3a2e4;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcce5f36bc55aa34c104048ed74933d826e03e22f29d001ba428542f1d3cbfeba359760c0631da91d17866d163f734bbcf4adcf39656af48ce23771ee80ddc1e82ee4d446ce8fe26c1f1e6fdb33cd11d44287773bea579806ef5ea025d146a98d775872ed2888c31370d56abaf444ae548;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd8373a3b742b3dbfd4ed896e8eba455151af3ad339e749e2b55e1ee611822fa01cc563fdb7e926c09956816e3274063d956cf812a2898f51a6c747c13f2be442b27f43c0b5d8e81b2c5df937bec99c8cd4568c61c76f11052afe1164db054b252e5283d522acfb2139e9c381d1e10a016;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h50d68a1727131d0648a57a18ece82a47555d34ad7a5378751f4f920e743ef4e7b49a0759c9112be6f5b4fac9b4044908a1b2474ac8930dc67ba13996d015c85e369510095215f73fbac86341b3e4da6fe3f78cb5c86c42908cf9dfd665b68ebbc0bc80859d4be90123b342567a152c69e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h95aab60bfaad821ac0dea5de6756a2ec0a6e8ebde450e843202b9a5044ce74715f5ca15be45f7d9b4dfa2ab7820edaa7895261c1b61c565e1ed456758ebddb3682e0af4e2e10fc191b93c1fb465135f1da3cff336d98e9cd8a78f5e998344f38847b74ade21dee98cb96060515ae3cd07;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h5d1d867aa4604e4f118888690a09eb653e9d8429e0bb67ea8d5aeb9f950f3f1310d92b6e27921d153aaba9e9cbc5c7e4654a8c5ecbab90baba2c02a614fc73ae8bb910d4942b1b8119642758997e0afb6575a6995588bbcc5fa0c80c698a6cfa102942bfa29a4af1ce37ae87f81be831;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7e85bd7a8bf23a0729a73a5172e61fb94eeb644dd76ac988f5fd4c957b037002d58422143a91d1ed1168b0d818a7aa45e30e8883e21fd08470d8424193883863b8c0a7c6647f841636699ffb423b0f8f5ecdfe85b55269afe878c15648d7c33046da035157157702a743564b53d9e5427;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h485bd7e2b639a4dd7bd7cc689dacc039146aa82c9145c3db8fe4a6623d94e1f02094fabbd47b2003b3c84612a8ec02f43437d86ab1c5093756a670190e727ec154adfafea45233b9e74acb44564520d53989b90713ddc06c0a0dab0c8f0a07677063f39f943ff1cd55b3de5e2439c620e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hfba0c5e91d78d6a3bdba58261a107c4d3f459f45ed4a0f80f4c2fa116d90591f83224a3c59277bbbf7e03f7fb25f797f7a1a75c4b999bc41de58050fd3ae9dff30424632c2a98206516e2b40f85fa18e6f09901ecdae7a785f8d572277c8b55df1e6a7caa4313692b24082e86b72ff6f5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28f0230bdbeb6b29ddc4744814f4920153a4ee27dc3ae9d1de3ffad428fc51df3e311670b2443b5300543c81bb23c4ca2a5271558d3acf1700148814388a558ba22e1353e1e0e35de07628366a60c457301962b85b374c1ca06a54b5b1cabc6e71e781071ddc9c9cd1b730e8ee72a81f3;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h397146c90759cbd9b4cbca4f20a4d9fbd13bc109401829b0da19270b336b836f14be8598247492b0635094921d2c520f2be79f232579fb86c02619e375e0debf4fc87fe0ac01dc11602cf4496b4962d1feb15269c3b1273c9d67910ebd95046dff11ad208d52cd79a9065613bdd779df0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h9f49a1079547356d6a48adcd407f1970c359ce20a9a130cd05b20c7e3e99cd387c7f79753c2d93ddd2c3972906ef00e0dabf2dc446a581fcc700c509587306b7990fe768312d6f2f445163f86305f8692e5b8e9f29bd7837c630e9173417c1fe1a0be08db777514f13e4faa44f1cdbd8e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h526572d2bb50930be3f38dea28f0801a3349a30e77a5de6a4c716b2c91ccedb1cad76fc68c9e8afc091e5d6c484e1e4b9d03f502f02c00836bf2c59535446b5d7ef84256498616c31653167a271f82ae2d31c6015c852785c5463e21871d4154f440c8cd8f587f270f4502d73b36cad8e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hde61da52a055916589e1de2ced505dfa96a10ba241113f4c4dfaf41434d60b548c23d2c88202c377d988d0371a3cfc4b501a9ef54b695ffc0a9840dcc3760b77234e763ca54d71a470e6fd83a1fc066f309652d7a7397e9809d817010db960fa4c64107c2da77ea784e9c8ed6930485ae;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h14d2b39232576cc884c419d2c576c1515f4d4ce50f5cc9ef2919616f6de6d6696954c2bbc00b2481d234625159de74b087a91b0435c740564b35648d610fef6b255e6f48785d65a5767edc8523fa5667236acfdf2a2ad234343c6e62e811e915f7408e193533b540d44baf854ec683f37;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b6c61778c2d26a9cdfd700ba70dee1892738e68bd5b5d15cabe94b159c2d8b2a2b312ec23054877668ee1e3841f558d7d3d23a28531e72da16787a5cced2c0aca98d7c2eb86d765751dab9d91e95f21511adf8acaa6c6f07451b2afc501e0de006bcd6a7aee08a7928f7f7a1a9be4a82;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h474bb028c1ca8e447f6df0dfd19adcd5a2c656a36e987992f9fa2fcbf3a23c782c89eb9fb9242faee4bab279d9a8dafd64cd673261d975f8f59cfe55e6067a1f5bed751cb90f6479cb90a562423376af0cd889190709c599b1eee759c1a5961813a0e4e7f6aa9e9c1157242565420ef63;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h13e7701423ff699bfa6dbca60a26a291ed1dc39aecd8b1dab75df763c9631400813eb57a89481d220fe988d2e834b4ccd97400622dd1a71a95162bfe2bd9c62069984df0be58c5af33f580f35e614a7f1aa7bbc194276fac00311aefa2ac91bd9a60e5b0c90c6633acbda0e9dd4ef9ef2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hc2d83b9b5e2624943dc15ff94d824cb91d68ed1fb1a2c93c76f9e1623a209bde96360345f5187a11fc19b540ed7d1a89d21fdfe294e037b95eed93166c878e0536773e8b1c287ce3de60308eef1ab80270f1765ac3069f6a82fd3cc5eb144a3679039372b162f22137684f29b161132ba;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcd69e63e0267522568b4e34b2a3ea7a140242a74d6fe58b4477273f1feb13d0756db80a92f042e7e02f20d6bbe4f39e303bf36bf3a402200dd730f8159babeb9810642eebd4a507099cd521d2957189af159f85d36272c968b58c83b8dfad387af61f7b6777c0628b47d986a60b70a026;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3a37973337c1799ec11c487468fdc141fbd5279f03de59c04ec3167346c8abc625cb2eeeafea832041b97a0955bb2f95d4cfed14c214c38b50146206bac13383bc4218ac640cfee0964404295a71918c2ee9c5dbd3661a625fc2cc31a1e3c2c02ed977301baa7f902b9f6083f591c0231;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h7df18589675f439e72f89d0d1d79bab545b6c9061422671b10868ae9f97bb71a90afcb48cb9ec95cee0d268aea96c45dd63532268457741e6eec2f9cbbd1ab78c331af4014aa1a99f47b82d9f661defe93b6df36c6805ce14dcf30ad533bbcc29a11ebb94a26ed9878f43c82ad5165961;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h812f1c546da7b360ec1a2212b36796153295ab4fbd7b776a5020af70d8843c6e52c0f648a8a04abaf732b2a4146685f61178db0d922406950baa02651947591c16d6984adb010f5d8fadf62a35881d2d547d6fe374b3e7ff4495e8059545fd34ae440b9c6ed1190a92223a3c2ac18b2d5;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h45dae9f0f090d83371558aa84243212d986a230f075d3cbfb4f977a68a24f8076faeccb03c2e47034346ba0b835c6cb8b27818d634bab34fa99cb50244a78f67d7fa201e2306e19ce7e439fde6451a3511e5aae9946c5468c8e812bffcd2bfead7c678a67eec7d9d8c70f1c319f0ba2f0;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcdcf42b4b5ab5c94a49542ebc1ddd7eb450424821ca2bd01ee21563466ee085926cf8111e99dfaecf93dfeb5b1e36fd7bed799ccdf20cec3a42fe539b18717528548e6d37305d3c87a369423db34b0c35b3fcc446400cb0ab1cb6f3c7759a9e6c69429de884d42a3ab1ac0b7d93c6252b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hcb2bfb6a6c730745c61c549fdaa73ab6eaa3f0465826ab0e6dba458a10e29b8b0029a3fc0b0db71b39dd50e91323d250fd7c58d7ce6d0a4ef134aded931b2c3406989a220b04a0eb0c98af61bc6bf516fe73df9b40b846e0ed2a684c87990b7405fbf2c6ebc9d69ba35663b0e35b0cce1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h8717d9d4d0c1f5f549575c3d87b2707fc218b5961a94254f94ff20c30f9a840a9047d8d1113794ef6366031a4cf5cdf4e02b65a997f97cd759b8380daf3496b88b6f8a59894c9936f08c7946cfba997c022b95ef040129872c3691226852fcec0abd97e159563fefafaed375aef6cc6e8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h66319e4b4f0aefb363949fadc76a1795f5b0334a18578d5c5cee94cc168f6bc327d772680ea145e16813af5515245480d4699d8b241937cdb1a454f743a8cdf79478a82a6c2bdd8795cb8ff3642dbc118845715eedf57b0492364a049e707553b5f57a19fbc41f2e0684fced2a4f9aff9;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hd970203f5651f6159308966207902c1de159d0287a496c75a9be0023adebbe4af86c41f09eecd3ce21846f79e881df0f201222a6f3bef811d662e9f0c040707567b859c0c8bb7ca11a2733c5de5271610a84de0e2124bedec0bb90f03451c494eced2e05f5bcdd204e54c43570438202b;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h3ade343dea51b80ed3654433cd42a32993697ec3a1af93779461e9c281c1037ff507d7b70a46d59f67a3eaa5f6115a814933bd7fdce1006fd97c624537829c7932494f2c4a5a7ae35280217a4d29089544aeb7141a48c1cb0830b22850df51b7a68638a5bd479834f7004cfe683dc3076;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h28746ec061dbfc6e4874f3ed8cff81f36a4a5e3ae9f7f34cbdf3aaeee82a4d0b79688ca0077c6358bd1eaf57a83d57d0bd05d7c4c9d3ac88c68e845a463e385c96f90f704bec4efa705b70e2398e17f5142850db0e36d4a572b5c237f2e1d129f697ef617018c814fb2d820d05dd91517;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h1b457a3039d929f76c38df20d0e1792fb8d223db58f01ce1616bd7b353d321c7a4803cdb793dd4d6999750388ef89b61c1a578cf48f2c79face495c4318d00602594ce61e89bc12f0ed3f0d13a192eb5663ccf10e3a230dc35a3436d54812ae1c0c197dd91aeee8da4dec959280684bf8;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6ffbeee2e433bcfef6dbea837fcc05fd313986409a095b9089b5f9f4001ceb2657bfca58b7d88d4e0ce4a0f5a969c0d89f7379bd8b197b7aaf07695da4d095a396c7edb5bc1308e374c1b7127063502bf7044beee5f77dbf22f6006fc00c519a35735b8eb8ff555f4e142152168dcf11e;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha986ceaffc8a01ab9a3f1a87b6d7c90f9544389b1424dca6d9121dc32e73eefd6aff7cbd73e574a8450d3ca1d6368e1e437adae277b8b5b2fdda56583b2d407ded25a7576bb4f66cc1eaa7b482801671a7b8ddfad81e6d77904dd2c3eb1732e54576c9aa82d94acb9bf75cacdd7f97b81;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h87d137158020500fd6abb5c727c6939b64bf0c396366c90a79486db0dda9ba8c5cc7dce0eb5171f86b0c6b077754e2f16c6f81fd03192891579a2e90f51e3f1fbd8002d84ad5643f544e5996975163d4ded7db836b1312e614b2f3e171c0b5cf373967dd8268dfb980ed29c556368d136;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h4f7ffd9fb8c45d891078cb5ef04fb619acd661d290362bba8cf0eeae1b395ad234b2d7727beb4c9918e277d54ea729b59caccc3f0772c7f04b662bbc1bf29c156ba02386a7c540f8a81d65591487bc518be2cf4506884b4897aac52c72256695b76117e4e869e8fffb6ddb007a11a2642;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'ha1e0a6afbcc3b4a2fcc712d2e9c33bbde8fe0d5b1360e61cf11f8eafa11a55a64b1e5f357459d04422cfb2e6077f6fe796bd8873e218fbb1edd7ced432f306bd268e54528358a58c279a1e483a17a4f91c0541b25e0054fd3a43e174ef56e75bbb44ce2bec6f3b10e99dfcf3ccd8232e1;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h96db55a25ffb3b52a4cd217c5d148d36009a48c0b7f422d23978272a490dbbf6e9008622d580bebc42ba00fedf1b65894ce84b9e42a81067c129ede7064bf27eadf2969666969e8d6ef822dacf264ba64139ac431ad4ea7989d5e5e05fdaf66bf1bfea8b58c566e8eda28df302f7f1b71;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h13b7fe9fdcd01e95973ba09072f8fd332733536c56db7a58d89608e2e74e543ff6e154604c0b304d54346872231f2008ed5bd6495f13555428869ca07fbbcd564c247b56b89c8d2123149a2f0055308bf1c060ac067dbef3de1c8f7595c50b15b19dbb33e6565c3465659a6f4e7bdddf2;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'h6cf1acdfd5e5d923d3a18df17c5e04856ac0679d0a79ab047a65ff2057b35900787bbddc26a9ffac0f62b87cf80e92367e2e6c018601c0d19d254f7c10039716da6cfa6fe3e30467338680cc37b939e2760145971592f2742607f74e0fce7dfaf518a7cfb5cadb4154a436f9e96921232;
        #1
        {src29, src28, src27, src26, src25, src24, src23, src22, src21, src20, src19, src18, src17, src16, src15, src14, src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 900'hdfd5d1844de441858bc67da76552790e2a1d27d0aba376eed8eca732d422f2a95772d85351dd07e7888e2319266b26d1145c4c1017a2c599dc50448de367d58119cac96fe2283800ca6292e7034eb507911cab4fb9ab854063f7f4005010273e20ce2bbd8fb3b2a01809d81e00e7d3bd9;
        #1
        $finish();
    end
endmodule
