module testbench();
    reg [13:0] src0;
    reg [13:0] src1;
    reg [13:0] src2;
    reg [13:0] src3;
    reg [13:0] src4;
    reg [13:0] src5;
    reg [13:0] src6;
    reg [13:0] src7;
    reg [13:0] src8;
    reg [13:0] src9;
    reg [13:0] src10;
    reg [13:0] src11;
    reg [13:0] src12;
    reg [13:0] src13;
    wire [0:0] dst0;
    wire [0:0] dst1;
    wire [0:0] dst2;
    wire [0:0] dst3;
    wire [0:0] dst4;
    wire [0:0] dst5;
    wire [0:0] dst6;
    wire [0:0] dst7;
    wire [0:0] dst8;
    wire [0:0] dst9;
    wire [0:0] dst10;
    wire [0:0] dst11;
    wire [0:0] dst12;
    wire [0:0] dst13;
    wire [0:0] dst14;
    wire [0:0] dst15;
    wire [0:0] dst16;
    wire [0:0] dst17;
    wire [17:0] srcsum;
    wire [17:0] dstsum;
    wire test;
    compressor compressor(
        .src0(src0),
        .src1(src1),
        .src2(src2),
        .src3(src3),
        .src4(src4),
        .src5(src5),
        .src6(src6),
        .src7(src7),
        .src8(src8),
        .src9(src9),
        .src10(src10),
        .src11(src11),
        .src12(src12),
        .src13(src13),
        .dst0(dst0),
        .dst1(dst1),
        .dst2(dst2),
        .dst3(dst3),
        .dst4(dst4),
        .dst5(dst5),
        .dst6(dst6),
        .dst7(dst7),
        .dst8(dst8),
        .dst9(dst9),
        .dst10(dst10),
        .dst11(dst11),
        .dst12(dst12),
        .dst13(dst13),
        .dst14(dst14),
        .dst15(dst15),
        .dst16(dst16),
        .dst17(dst17));
    assign srcsum = ((src0[0] + src0[1] + src0[2] + src0[3] + src0[4] + src0[5] + src0[6] + src0[7] + src0[8] + src0[9] + src0[10] + src0[11] + src0[12] + src0[13])<<0) + ((src1[0] + src1[1] + src1[2] + src1[3] + src1[4] + src1[5] + src1[6] + src1[7] + src1[8] + src1[9] + src1[10] + src1[11] + src1[12] + src1[13])<<1) + ((src2[0] + src2[1] + src2[2] + src2[3] + src2[4] + src2[5] + src2[6] + src2[7] + src2[8] + src2[9] + src2[10] + src2[11] + src2[12] + src2[13])<<2) + ((src3[0] + src3[1] + src3[2] + src3[3] + src3[4] + src3[5] + src3[6] + src3[7] + src3[8] + src3[9] + src3[10] + src3[11] + src3[12] + src3[13])<<3) + ((src4[0] + src4[1] + src4[2] + src4[3] + src4[4] + src4[5] + src4[6] + src4[7] + src4[8] + src4[9] + src4[10] + src4[11] + src4[12] + src4[13])<<4) + ((src5[0] + src5[1] + src5[2] + src5[3] + src5[4] + src5[5] + src5[6] + src5[7] + src5[8] + src5[9] + src5[10] + src5[11] + src5[12] + src5[13])<<5) + ((src6[0] + src6[1] + src6[2] + src6[3] + src6[4] + src6[5] + src6[6] + src6[7] + src6[8] + src6[9] + src6[10] + src6[11] + src6[12] + src6[13])<<6) + ((src7[0] + src7[1] + src7[2] + src7[3] + src7[4] + src7[5] + src7[6] + src7[7] + src7[8] + src7[9] + src7[10] + src7[11] + src7[12] + src7[13])<<7) + ((src8[0] + src8[1] + src8[2] + src8[3] + src8[4] + src8[5] + src8[6] + src8[7] + src8[8] + src8[9] + src8[10] + src8[11] + src8[12] + src8[13])<<8) + ((src9[0] + src9[1] + src9[2] + src9[3] + src9[4] + src9[5] + src9[6] + src9[7] + src9[8] + src9[9] + src9[10] + src9[11] + src9[12] + src9[13])<<9) + ((src10[0] + src10[1] + src10[2] + src10[3] + src10[4] + src10[5] + src10[6] + src10[7] + src10[8] + src10[9] + src10[10] + src10[11] + src10[12] + src10[13])<<10) + ((src11[0] + src11[1] + src11[2] + src11[3] + src11[4] + src11[5] + src11[6] + src11[7] + src11[8] + src11[9] + src11[10] + src11[11] + src11[12] + src11[13])<<11) + ((src12[0] + src12[1] + src12[2] + src12[3] + src12[4] + src12[5] + src12[6] + src12[7] + src12[8] + src12[9] + src12[10] + src12[11] + src12[12] + src12[13])<<12) + ((src13[0] + src13[1] + src13[2] + src13[3] + src13[4] + src13[5] + src13[6] + src13[7] + src13[8] + src13[9] + src13[10] + src13[11] + src13[12] + src13[13])<<13);
    assign dstsum = ((dst0[0])<<0) + ((dst1[0])<<1) + ((dst2[0])<<2) + ((dst3[0])<<3) + ((dst4[0])<<4) + ((dst5[0])<<5) + ((dst6[0])<<6) + ((dst7[0])<<7) + ((dst8[0])<<8) + ((dst9[0])<<9) + ((dst10[0])<<10) + ((dst11[0])<<11) + ((dst12[0])<<12) + ((dst13[0])<<13) + ((dst14[0])<<14) + ((dst15[0])<<15) + ((dst16[0])<<16) + ((dst17[0])<<17);
    assign test = srcsum == dstsum;
    initial begin
        $monitor("srcsum: 0x%x, dstsum: 0x%x, test: %x", srcsum, dstsum, test);
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfffffffffffffffffffffffffffffffffffffffffffffffff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6141e4a295c3f113f6348655725a99def75065017e9d14bd4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hebe47e5e2b239122642c5e996d51c56d98645458d54e9fb84;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hffae5e5b011dfac94e722a2308b6c54a0d94db89ce4e6fefe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h743f66ac976745803981ed9d4de0f77f1eb4e72988fd3aaae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5907777ab499dadc25ee4456f284e533561f5f6defc117ab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86494a1165411c339bf8773d573c7b3918ba35de1c91449a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h445ec90a7790d743a34a9a13ab6decd5ebe2e2d064a53fd7d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc07793bc0f55cc9394b0450f088c9310c1ca83a69805269e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a1791d276706cc8680e40846f5d792e9b943662582b902f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1c8c3eb4e8dd77f0e280955bfbbf026ca473f91f3a73e72c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h615d7e3a7f8acb6164dfbd5fa5c1218f692555602e809cf0c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32daeec63c859735fb8f6b302d400c28e2fef5d4372e63b6e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a28904b32d58ff883eff0e21cebfa5d7d94aab5f85d9df6f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc10f48482ea48fe5afc13ac593e85beef5d41661282b4e137;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1aaa5c151d2ae4bc749d593ea1ac1456bac5ed8d6eaa4667;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14493a7cb129f554d02a29968892ee7486a065ff262291e0b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h939716d209b9ce4c16bd69be79f7374a3681f2e50d7641db7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h350c3a524c1448c74d45cfc60a87cc7e6f688156e27fb506e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b2af5793ce8a7c5bdf74982dc3c96e121b358c86258344e4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h142c27372243abce1d63c8929a11e6f9e3c6718929344306d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hefc620cc8e721c497f55632998c6941e2a98dba3384319b5b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ecdf6ab1be840171e4e08b0013754759feab262d525198a9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7054061f3a1290be8807232e7c988180a522d69a901f1cc5a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2d54b9be5b316e7b09a5caaed2c118aef9a1fad434c62b4f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf22a824bde399ec2bb6df813ee80eb9378c5468c6c33709c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f8085ee130e293e9c2074468ff4748b16634bb40596155a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a32635bf1e160bd0cf268277b3132480237457f3ce1fc9f3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfde1c1ab6e758d3f6ea848123e66d5a19a9bf5d7c930163b5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd88b5520afc8a7ec9283529a4afc76a6f42b5ab1cee964033;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd6b5ab67614f8cdd360aea437b772ba6a311fcde31150a085;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a42d582850cf609321114a5403fd988c94bb2256525f83c0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e0757caea46ccfdf21bd8155132930d117be1fa33d71db88;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbea999cd2670d94c88ef206381c2a9e89fed394107a678922;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf146d96cd61b2018ff1867f90d011d9032cb29c965fa9472;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h687446cd539ab7ac35caa0b54682a4a682f8cc3dd289e675d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdef2b3753f4b115f67eb5e909447638056cd118f7068a8d1c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28577356c83e43e16ff2394ba25d26bc3374dda73ac5a549;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h385fbe8f3f81608fc45398a20506ad722bd6536d4c4cb3c84;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h592e7d5186454fa00cd04c07745243d6e69efc74927f55d14;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa9433e0d9cd54521c54feda0b92eba292f64cace20e86ba7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54f766255c2fabe420a731ce402d3165d161d64d3d3b581e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h580a7ccaa9adcd336e0587124621f0119256927e36acbd0a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6de06ba98fad6a19723e23353f031deb83e7cb1ca55f36e7b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e6d3971f81d2b9af923780e7e74c2bbee7d343903ca26ffc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hacfdb383048fc3e40228191b909c053edb5df56c7208a7a43;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f47ebb96e7812ac083ad73ff7112f7ecf7003989e6adce55;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ae8cd1632f263f6022010c94cb0c4f8bf5dbba1e9079d614;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h676f6f5906b7bd4a02ce3854928c25f1008b7782a61cd37f4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f82e302564ba7fdca8ac9f990459896bd39080b05eb8d107;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h42ff2cf4657834638f02220acaff1f2223c40741d18f69a68;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2690466d8e15a5000abd53ac0962a1307502274e3f115c31e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32aff535cb21e8d7fde9a3772c3761b821cc6c955db98fe28;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce4054ba5b256532469771811591308c9d1d075f8fe915c89;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he515e7b1de207ebaa5ce5a8f9dc297e2762cabebe18b3e300;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h945128ffdd2b08be9fa02d6bb5642e5054c3d84f78f5cb9c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9461cc7ed82ad7835b6442bb121bb2dce9ca004bf7f05fc48;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8ec011c2b7eef7af54d4472229794d919f4c98ecad9cba8a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfafa2cb65b5380021f004873c42fc2aad6f16bb75a043ad35;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f85663820809d9bf6b5a855fc7623569a439705d742fc48e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4bcfe6c01abbfb9f91ab21c8a13d04d145a9305f99f0d955;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a9160f18c115e74ea5879024ee1e31d74e6879347067ffaa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7eef16210c5d12bfeb1203c7c8759b9e84527530f38fab3d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h603826a49b3b66245d6dc68cd1690670ef846638c3217a73e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf036bb150cb2fee0ca6203e6192c62bf03fb39d631782c629;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4487c00476746d7cf002e01e1e54af9b5ef120a9be0e9ac20;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2ff5e81b912e3176edda4aa6e4a2347ab4048052ecd44bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c0f6b1be19707665d465ac7e0d89daee7115998e3571444f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7e6c8f240a1d42444a119a8461ae8bef2f72305dc19af54d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5d50f1141c730c6e6dd0af4fe3a8297070e56cc335e6de7b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c15778d76b8bf012677a37d839d352ea01d0c8e535914e4f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h388ad590845a249fde37baeffa14b5422d352bee7b31b265d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4fe3f5be6904dd739fd4a85a67854cba62b663fa9847916de;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0dae57df678a301550e15f174e6d8636e2ed8566c5bc39bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc82b148a8d61c6c87b7ca0b4ffa8740f8d9952f2397ada61d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ecb69a64dc0f209b710071b43c1019ab8c5e8bbf6a8074f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha952324ac8ebf7ad67dca78c6efd7cb43e27ec6d279192625;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf662f0691f0c5fd4010d5c0ef43163d5fe9df6c9eed94a576;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0186fae73991e0e4f9af13b1c5001792dba9c0740a8d8b0e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd61a7d9122b4f3e197842ae1bad6873eac3a5458d36f29a97;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd035a837e773e0c8195b55fc1a797897aa9da75810b71d99d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha5e2193635deafe6c0da8c163a370b54ef0799a88a1a2e19;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22b207aa9f70733cbe48b8af90d71210ddaf593d0254d6520;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a934f382177ba0bfe16265906a94f3ff2198f6dbfa31fa8c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25e248ada85ef44921ca5095f505ea2f1b5edf2a55c43e71c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a89206ce14925fe6fbe3096aa1b01e86a7e65b36c33805e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he8c7b349a69cf0dff14c81c55f38c48400dfb41adbb827dee;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h723f3782b57761246280b4f8fe2af1204b2c34a705dd77587;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f3a6eb476eb83ff826b71f091646cb55d2a6c07c0ccb2b4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9571a1f2e570622c9275d89c97b841534198a5d5ef385458a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he6dcb284b52ae1ff944a815d6ce4a091af47427549859232d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c172ee1f489e6df04cc77abf9fdd560db8196b566ff7984;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h51d0b0db32be516b72b9f747cafcb6a2be3623b657203b9bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e223dd0c4e4f3ffcd9dca8592b34a570fc66bfa495991c33;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b6f3ed6579a98432a80f707456032100d09264eceed79855;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he020c45f76181e91153ba023473d13bd60486321215df9d1a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a86680401a940bdd89c26de9fd6af02b5572632bfe6d9a6c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h835f555fa617a927b683d54a6a308d27778465d9efe55999d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h338ef5592cc043ab68aea709649a5ab2ecd9490c2d4f43d34;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5db8348903ae0e7115e3887b660562630ea1ab16b3655389;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd388fe340c8988dc10d58aed80ddb9c220d645ab02ca657f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ee31f8e7c72f506f55b751fac97f5ac254ba3d3b240275ca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95320c291a9b44b02b3aeb495cc4cd729ff28535f16deb001;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6dac9d4103d7122010a9aa73430756e2b8543822ff1b7646b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa24e3d8c75b958bf72c78e6cfd9b8be6f2eb422ad7d01e5c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4115e18d7c8d07d447802f9241f9d574a9deb8f9c72929afb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha16c6e1d85b00013903f9b0b26672c2f672eab13c5a0c1e3f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96bfb1c840d30d744cddb8f786e29b634c627cd1c53a178;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c6bb2d2e9d66bfd5d7caded9c9f0efeeddc1afa4e884336f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8321aacb0600e1fc396b66d8459eda9befe665900c1bdb307;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d3e790af5eecf7d2f0628eb1f6e244f49e309f88e5f5ca0e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf683e82189a97c4c8b1277f391917b1a9328f3e17aa75e9b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4201d61f4c7aae057cd781207dcd70d5dacb715c392a21c8d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba0d1b4cfd4a5f03c1c073c5e8d79b3561f8e91e6e39c0ccc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1a86aba568dbb31453fc81f36c3a5afee5dc29d0ef1877148;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8a8938a40211aa6ca5ab147f9f63e9d7f73c67a36e4e4e1c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h43d04b18a6e157a672930b246148078d09a5461750515d92;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h352b88d215f1e61693dee16d92d6ab29e1cbd8d7bff9d3fe9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h665b0b4cccb2421e278f6fb1b03c702b8e41f929be6a0548e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4824c986a2ee2b06d1fff502414ae0956f237f46049fd2b04;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7145c73294764a6324ec7372ade6e3c154b5475f161bc1517;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h672c2acfcdef340daa80a9b1c172721bb5aa3a0831fccc6c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f0a1206f8162b04e0d1d1aabe4d0a95c9e09937800f1bb5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc1eaaf4d736efe0bbc251b7d8e3ae57ac5a0cb8d32fcd5cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf98e4d87cf7e5e19ee9415a84f876595b1c900c2e46e05e09;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9b4d2ce79d913a701002816d0ff8214d5808f134ea73da0a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf150da82a5daa079b8f5456a22b4858ae1391de7c27c6a8c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hec95803ae521bd725afd1d08fa8db9fcf45b8b3bcf92be85e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3cf3eaef6ef6c0f6d9a5102f10fe669b64c62d45a9686c57;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c5b5360f521274262d3f4301f240bf94116928a2c53544c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20da069866aa83ad4e52e69f447c5efe3975b5235ee036c1c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc16cf65a8cdbcf551c437ce624f3e97135d27f803729bbb3c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb39b494b50e7f2a3acc8141e74e193424726d1e4a43033754;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74e01ce8b97a06dff09611c6a212339a11b1fa11ed52e9de4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1818d88d6cd05b4641de39db3a406e3bc1c61803cb2993f7b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haccca4b1c9f0171b4412e092de3222ac6a3923b83b1e94669;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he8e9908dc28310d9debc6d2cbe2e10b85b248d891ad0a2ffb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he85d389e200047b09c4dc55576e2215fdd4d02d32955fce6b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha25a84e1f0cc0f765661f474dbdef068d2c236c57a73d30ca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45e51596488cefb593b93e262fbf58f2865531f1c40f07df1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h539739dc2b0f20a8a13922c577ffb8e3724a9b99ee7a17964;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe6b02e5231f40dc0def6c38eff80c93ba581d9e7ca445e44;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h23bd3401fd8e74f35f68f70f819dc86fd20f6f268310d739e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb1227c1a64ecd6d7179b9a66e8498c42fb6f86bee559bf49;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he38321d2dba32edc6d6b604661aba70b052b09c07625ea15d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb5fe9cdba674dafa1cb99d682f799140c7cdf4bd96a1bd4b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d90f1a6ff43de0b4b1c09b5b60e68c3a2ca20a20bea76141;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49971de4b4807046d3aa8be0341e824f80aa488ae0b3bb2e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4326b16e9dd4cb20fcf321b28499db65bc8e03095f49cb9d5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60f4dffaddbe09b20e0c4c03dbca3a2c945ca1a7339c48634;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa29712f144f933f22bf2b883dd219a0c8707d241a190de5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1962faa9090fa370b8bace0c5dfe9f0b6f02c4146a686fe52;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6aa0a64cb662609259ec3e6e8f0fc8dbb868622a487061364;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha78e18cbd4a282b50f6a4add49b76e306a6facedadc3ed790;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bb80dd56fb23ecca52356f888799b7060e185203f6ac2511;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9b129baabf740539a3010ced8dcc13a5f61d2df90cfb1734;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9450bdb62d54e8470b42577c8b0ef164bf6f2f7579aec2236;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe21affb2bb2c6059a8339e26d12f513edd30580a4f2d6084;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77ba5a944949f4a48cb47d5878e8bb625fcc06baa72f54996;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6651731fcb36720725d2415dd714999a696ad6164686e5f6f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h319e2f11085f264a045bd2ab4b5a79dd755972d3b3f3584d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4b7371cd44995546e3b0f13e0ad0bcecf384f34ca877e16e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d36d38cc2270840a0df7ba00aca58c290dbc0a71cbd6bd84;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h360ceaea214a41839ad11e602ba874fa7dc0d4ce1f9e87f70;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25a85a1ac0ff7210d6cecd8d1966dec44712ea46af39a8be5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h340ddbc88e3167df6e9d011aa53fa30f84f3b647bbdebe533;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37a5fd7c39f506568105b35a8f4b29eb5e1cdcb5c7b57a52;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c9b92045196f892d8bd76ca31f5243c266e8b33145b8e84;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc8165f134ce439c5ac3f0bbaac1d3e4de4b071db23497546;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0c8655615da0d28b061181688a00b7595151fdc41d7b35db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60e0b4e53d366a8c4017f780ba2cb318e0cf4ee8d3c4d39c5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h237c7250a62973803031c2d341c31d3f91a63d1c7b5a4dc82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9da7e04aa516040b9d7f52fe9a022f8ecc6cc0721f531d3a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9de97b1a036dec3d3a196e8b264728d57523dadcee61839e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hacc1b8d77f03263ca3564066a2659e2e06283ee8a919377af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2ecc9e52aa33b34b0c61f124653bde08666c682f4956a88b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'habeb0f754d0c9f918b2d59f175c4817270c92f5b558590827;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1677de255b65cd58729bb05272674b3558d4d519ebd2e4d10;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e7f50653cf894eea7776d618e924d7cd075a0853083303bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc4fcc5a72754862ad20d6f02bd7b6765a23352a6490f741b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b97374ef855e3e707c79145e86b4889a71ef7fe8be97bb69;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28e157d64d9848c846c1278401fd2f4208bc247e04a08537e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf364054fc5d5e63eb3c3d3a521a729c5bcb8d9ad4281e0ca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h564fc4acb33b2823d10470726908f846d41f9ac4eabddc66;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2182372c54d0d1251bb41f5b4c1d457d2d21e00d9273efacd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3eb6c0207ba3fdd9522f31bb8bfa0ff3300c74ea40e1a22d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95241921d7bec939acbd7668eb064790f2b3c1ab39f981add;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54452ae92cd4a6ca4c109e2d64a624adfe4d4f27a3c9bd089;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2d49e683962f9131e2decd619f9affa56c93ae8fcc4814af9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21297b32ec1ad93d3e439e7133f3564baead820fc5712ecd4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d3bb84fd85f60afaa79bc4ec6004bb9d7cfa53d5d90100e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfd071a5057abe1aa243f53257da1cf774a615e69c9de48fb5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29a99c52cfdeb3e4ea7084af589081f9c45243421947d1cf3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hacf94e5ba254b17880a222e2199d78721e753a9c2120a01e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h421379e7b36e84217b7781da7a59993ec14757f76a9bb0d5d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd1e12e43d391d305a99508bee09622afd6e7fb8a43f58548;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75fcbe5f912ce9e54cd6be4b6249a31dead7524cbd95e5db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h85c62ca56d632535553f98797d6afedfa2765a3c208cf37f3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a4749a2747342939fa48bd9a27d91a946111486880b6589d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd46e1fe94847a8da240e0b02156aa29e9360464092068a9f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9aea2307f19148159b96f91c5a9d094cc8db00b4775e8bc27;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58b81e03fe346c2df3c8f48c6e10734ca11e0c32ed5c078e4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4dbb8579941a6c4827fb6ea0c5ff8cd1fcc1be6cc070e5b6d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8fc86465eb32cf0dc01ce9e82d1b2ec31bb2566d79701d6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7bb59ae08d1689e16410e3d11e757ea68e6c6731a57583102;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc3cd341489df9620d55ed0cc888189aaa083678fa2c79e1a4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1639b89dd3a3f66b6c186f8ab67f3ed9362b331e20d5be6fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf90c7a30262f0f1ee87f95e90ff198b8b357846853997908b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb32cb460b4965cce78830fdeb086167b0e94c5f0c93b10f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2fb08a9780106ed50116633cfb98bb1b5029d72de366492c3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbc2e4b08f9adde7b3e016a5130b2ddd54d0a11f3ff5299f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9eb4cf17f093db6bde94b63017ae89c065a1f61597ec8cc14;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h653f0954ac3ac854fc60bf75a77356faf5eb9b068d90b3e10;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf03117824df81f1eb1c9c7bea5c0560359ee362aae4edc6ce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e2f1529125b6dc64f9fa1d741d16afd0c80ee1b4ce6b317c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c5dff644c9be78ffeae817fcebd8717412a29004cef509a1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha550393096ab222d9c35722cc5100761531eaaeaeece19728;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha194b550afd5d61071650ac24e0e7eaf6a952fe875a22d009;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c8a8694b576696761553884b449d0be0f9022c65bfac5d01;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haca636f581e4a71dae1932529560b408b78d7c752af766833;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb69d9ce81479a177e518e110580984f1f5e4e8f427639771;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76dfbbc550baf68ceef4bd470e06012da9d6774d584c755cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e1f7b3c8460ca25721c50e28ae70154e39834bba83bd8ea3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf2a598baeaadbdf0b9697aa3d9666a7332063df59a5415f7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h841f9d1e5fc70575a05cfa6e04f1631470078f8698485f7e6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7bbfd5e9f03e9b151ba6c5d1a3e151428c49486dffe43fcae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he59992977b074a75e7e9d94378d264c1e60dbde31cf01951b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c6de3381c231bb15648c7ecacd2e44cb47bf9bd9ed13898;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf84b3d6ef54c3a57be40825e89d1e43775d7fd2c2bddc0441;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbaed1ef213553e0313344062a40aa6067c92ee1ee9b4fe645;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf65378146be21d3d17156a41182bfce0d12fbdf9f2f3f4573;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f6443906008448f348b24f695fba5821642a9749948f548f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6634b07c90791f6415b4d196990c94b8d00ab386f56f82393;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93942fe3f71f77a49077ede36799c6463250a7beb6de1b25c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h367250f6934f86d5b32d9c7ff56706bebabc336b1487f1ce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49d16b93756090a5bf18e8db84f841495ae90ba9c1c324640;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf2b277f4cddd651e36a73a62374de729b021b5a2e32896b7f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8182f715c670e83d1e0041c634de99315d59f34d00ad2afb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5122b09020259f90a5483f1379046037500d04652decf1bbe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd616ea6585d024915b768773726621fa4a93eb0001567f5a8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17ebb43d3d3a3457e4fc878d11e611e61bb3aa06bcd1669c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6eb57b3c70500c3c6d89d6703c69e600c8ac57c7dce2f029b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h902867102b6e816bbfa372470923df4c742800ceaf3fbcef3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7084eacdc8b980b0fc79df35d8593f89ec00db13fa2949151;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb81f5385b80e9099d0d02b930877941d18a73177d4be910d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc63102c75670b6694ba21cc6c86f40120b92e1f32e176768;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d942666852d68f7b05d1876a677e525c27ffd50b48b01a44;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h45844eb368d91b6a89f0aed85e8509014465c6f59e0e77afe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ed63e66e6bd3c39870e3fb7a087782f4b416bc2238e64c6f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4738281e564a7b17b8ae72c06ed7474c2e43952504d70f0d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98d925ca5deed242850bcdd06d71d916f0c9322a58c14fa95;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h668d00ed369f09634b3b357d3e669ff46a5dfe1d18d112712;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h64275c118fa5ec29ab9f3d134e6af11b6e6509adcb80c2c06;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8d7bacc5518fbb5aa0148d642d7906fa84a6183474dcf136;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he62ebfeb351713a8a92b38d0eecb2be4213548790aeb19056;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ae8ab4e48293c32986714260f79079148320328e172ba31b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haf6796d3a5dec30f309b980b540e02bdd70b9f78d9377e010;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc50118732810f3f886e292271eb2431c23ef7cb3c75634d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b76f8d7978d3a6f36c14ac7f5096cadfee4a23e5d39dc83c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'habb09d0305ccb69d72f80dcc70096f4cd7129dca0f82af3e4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3ad310c6e5e74c4d9fa878b6bf6402fab6af511053f154ad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc81ca7f206fc21e7c7e09714af721bc44a66f4697df355b8a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50959bdde00b08a2335c190b6dfc3abdf9ffb68617acfbee8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef332e2af0af7d13397d842bf5516883a8b9d303c017519a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6dc50fcce2b4d32e85dd0ce47ec9d29b7848b6cfdb5a4140;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf51490cee7ec0196b2187aed83fd31467b993a9db806e238;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7c562ee7e863af687b92b282f351efc64e46c2a097658e7fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3282e5d8ae8f25e7bee50508005a75caeddfcf3fa53f5c8a4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4149cb658da3d248f5d8964c3a76552f9673885acbaf9de5c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h884652bf541dd807ed0d41b1c649178651164f7eb4e552824;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60c1265912a18ee63f43fefa1d6b2906b82187a0079e3075c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7f650fde522585a62f3d447f837786be3cfcb12acbe61ccf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce02196649c6e323fee0b8264193a613a822496b0422c29f2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb566917556393d1befe2267dc155124affcba41c7d653d788;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab381abf5a29dc1635fcd298e35fa79b377dc35d7641ff53a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b83986300fd73e7002e330bb19cb193fc41fdbb89da92f62;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h15cdddce4bdfdf9463c7914bbf491b28fbe177e43f96162d1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba8abcddec535a754b6c1e5178e3430847ca6944decef5fa7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he08d7649296fb4ad4066c97ad00a8bb8a99ff16815f8ff52a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha43922f9d6e8007286fd044d0ff0c2753cf30c8fe737acfba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae7751e3b5e157dca554836777f3b0a3467a33c42b916727a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d9f557b2a4b5429493628cf1ae1bf904091eb51585def7d5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe2a6afd212ae7a37cc97197889b599009dda420513ed140;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8883158372c000243e21dfe8b1e5b625c04c8bc09b905af4e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73122c940fcc9d58138115f615abd533d8bb3b8acb1699ea1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d2d821ecdbd9d04900df63b7775d96a7356d6426a570483b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5789e22274ad8ed76dba08ea91b2753479ad656a69485001;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5dda482192462db8d0135fa8386058df58d46eec500e7ec4a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37b7028d392f8478d6c9406a5e9dce1ae15b0162698d5659f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e721ab93bc60d7b8b57f9c6e1875ceaa8456233b8327f387;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f2dced3bfbeb1b5022c8cb0e6d3bfd39835bb84f29c80a21;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c4a63caff9823878d9b4c8f9e9bd812f140912784d11fc0a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70856487da5ed67a368db71b00994e2d10c42380c1bf855fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he51899166620f514d380d04909f8103608ae074ede2198057;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h732555284dd3e818e861b58321832cb3426d42ea7b6093f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he670e23ee3cf3f008e32de6524bb39e6a8c60864a8031b21e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29eb23697cdfef1ef9e1a88a3cf832bb6a6ffaa7f8d26ac1d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc59a4789b402b0990cc9d467c0ce3db12f9afd20c2a78adc5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h696fd1f9af1a013a0b4356962cdd81238f22a87c3b3481120;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h779700a41e049d0c7b468f9971bfffb60e0b065885d31ef52;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf48b43e79373ac786ab4a36a7a223e15785b75dfd2923ea7b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h541479a36c56422402e7488d592c04ac1779cb289c2f39a2f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf1b737fd54d58f84119a95a64e1c7ba7bc00af4448bb7e38;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7dba487f3c9c70bce3fe60a7da8aa9f0da1068f11601c6d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h668f0a4eb8e1db2fde793ced1c197fb94c35bea9ef406a7b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h802428ad68002d93fa8294033dd954f4cd3f8d8dcc7960a35;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ec914a16893e2fcff612f79f1db3672712e05fda5447729;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbf55947018dafa4ae3859a4fc59c58a6ecfce1e2a8d8d11;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f6254dba1a6576ac5266f9662b9dfac0d1e790b368e1289e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heed37299493781d9db929b6fce0deeadecedac2de2cefdc11;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22870276bbaaecedefb684cd82546573f579ee69db93165e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'habcf89dec404a7619eb4552ca9c8ac0dc7797e183dd3b299a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hedc3b9356cb654db7bf7b23c99e161070bf47710d7408c7ff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h52d1c2ad7ec8ee867f0c18e2bb65a857bdfd4ab7a5a202e55;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf20bb7b048f409cd939d1a8a64da0183c2e4f5fc162ffec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3e4ff746aa9a12673a697e23f9f7b7d74eb4580e9e5fe435;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h43313fd8d8df0a15a4290507b7931e33845ba069d03e17e7d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8c61d9b5d0ad6251d99e5fd346db54e0636bb966e5a7a6103;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59f9e333c1dd6b616b85caccf030f25be8f2058c873edde21;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2f27a85ebd2e024deb4921adbb4c9b73aafbb3e107461878a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf721f13ad194fd83a62b0bc243f390c9e6bb93fcf8e9dcce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc67a478cb86c8dfd4b062b45fadfd807c29014e5275cf0047;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he03e1b543cd19af7ea23387de7d95c1c6b87f3610a7d7d2f2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h333ac522d7eeb6e56772803b9c8d524a11f74f491a98c2ef4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4d81d72910148c1a8575bae648b614b4fb0e729f67a1b62c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h97f99473d44421a850fb06ad467e0fb33e7beaf377a84b89a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24fe0a59361b0f930e5741f2618d0a539bfee90120854cfcb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc528e3320ac2f627aff0442cdd50567e2ffd69190f0b31354;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6ab650d89856ac20ee0249817a0fb7b69e3d0c93ec90184f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75c1199f03d8e3f9a9b87ba55fa7b34045a60a810dd670bb3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb4c7d6fdbd8181d08438936c4270210f74fc336954983257;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1cf5c5c7b918be2fb9a0a3fdf2fe94d585683bdccb7fa668d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h57759be8ac2c3e27c78093fe07d6f029d64c895ff7082608e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89605c092d2106eab6cc4482446a3628c9818986244fce3f7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8203c52717d90194f84f9431acceebc7ad47713191365631;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h799e523a625e3d6a9a92b71e619dd13547af2ea016def7396;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7fbdc1030ea2611e14f6f67d54feb7c171c117ac63dfce7b9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1914aa43aaacdc82168e4c220203c84b6cf9ec7bdcd5ac3a4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha74c93ff0eeb27a7a259b33b4433832d9092a6491cd6562e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ad8cd062ad1f2e4af12af84d129c49f96dee4184acab45e6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f7e6162bfb425a6d9ea656cd9bef6ed37be8a86d307fc481;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb1fa7fa150c5c7a11c3a9fe7724298e9716669f046bf5e53;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd20c4e6d37f590256ff816989c95205d9d7a5a2c1200224f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h678ae8204e47bb4026e7c643c17df5ed286224a6ad10f7009;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb664454dd4e2d30a99a90f92ccb1d8aa933ac395b6a523066;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ef86b563c5c10b1d38c3ce41b0672ac4eb64e13842ad4f29;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc630de3dfb44ca70f5e78dab20180388393579feac524010;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24003457391e931c50405ddc4d802735ec1ccfc184541a112;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1159e51023eb92fb1067e0bcf4f9c8ea424813ff0f764e62;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3acfc393eb47bc7f66e8aa4aef233d28987c640e912cff64e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h82deda4df385fbc64e0e06e1f75a2e115ca1f3bbfe393c4de;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb7de36c0f6e89a6de5ab6012e8b539412e8ef3a45302a332;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h29388e5713393c67501e612da01f5e93a7b85f32d32108a50;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf39367e51281418c4d526193ce20d42c26aa9054244f4ecd4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heca0b231789ef6f094091010dc56d1504e72c04695b705487;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h156842abe8a9f2333ef1449c660e48905b6c721a8056cb166;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hafde9313335917320787a787d013b46242c8372880b0b447;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d640dff3d6ee39dcb11c0eec69404b8ccd4900306dd68adf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf9b8299c23f67af23e37091e33a4af7b586e9b44833c8c451;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e9f8c7aa89bdd4586f0af6b78454595b34e61c316e26fffb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e00f0a810910c13527afdb035a0db60d1300048e7161fb52;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5fb809765c028c57ca8b1d1dc06117631be216615f302f877;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdc4e505c505477d3a4252634d1d5f12e11fcd27a5285c3586;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb390013cfe25a016765c09d7ba83c48daafd074ec348ad3c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27394861a767a823c62d491914d571a77bf6fdc5f15213d17;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8a486b29a6aa54821a29e904a3d41f262595333bf384f649;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99ae63bb9102891c418656f77332433a2728374b046fc3d62;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6f666688b6d3bd23991ab37e04ffd1fd95b70fe756011f259;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce31b3be2bd68b430cb7caf3283f0c427dd73acd0e4436edf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8e45306fc04302f1dc6ebd8be85c04403926ca96a0778f76d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3cc7ffaf83d43186f8ebe62d411804c0eaf777bb3c8c04d96;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9078406a19d55b6c7772f96d972e3b66eff978576d14aeffa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbca549a553c094296812bd5d188dbc71d9270c257bec030f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24ea528e70da516b6f94196e8e01e88df2e3227d50919ebd8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha35d516e8ba3b6138d5a40ff20e48c65573c95416d7bbe7e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3453ccc72de0b3fa6f2c46c78c2e80b6fd1a4ddb2a419c529;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde6d22aa1f7cb8559fdad6e343c4bfe7012ea635ef602585c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h288360addba69e4bd549b79fe8427a41e1650e41e4baa0888;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50c22ef848a2763e487e71eda8e8a764de4844c337d65bda9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9428e63ec8f3ed06b1b15b6e33e23a3381c9e8f80341d1f3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h523bb1c0cb1eee97005caafa7aa1320e8f34a525e530bdcc7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6da9ec29c11fcc0327a07a089cfdaf980575c3236783c2eb2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d491ab227f9c6b065ee199f534e58ff66f0c2d81e60f496a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d1c44ff1912e15f34f5bf64f95a25fb24493afb59a604fe6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0ff578a3055051cfc4baebc95f5a4b917bce7e512c0f0d35;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5736116d2035e3c021f6cbcfd4d2c4d236410b78e126b8b76;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc118c2b2dd19299c5334e01934f42e1aebaa874c06c0f17fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9665fb824684573a15755c8d4e7dd4e229bd1a65483d06eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7776a57c87fb6603524fbe928ea4eb8d66b7f01aaa7ce63d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc8b5e6af24e5d0535a9073daeb20c71354f1dc52c84ef9abc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf36221d57add05110d1131b7657bbb19f20c8d4e33386904;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1c7fe8622ca17e436fff4072c063eddcaaed58a1f978f9a77;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8206cd358a7e1e0587d28f407b57d94f07242a9852da9612a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0540aeda67da8166dbcde9288874bd7eadb4cf8c24a39737;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6b5cd769d0be3a3fc8bac4b772712ef1c4551252f9dd57e0a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65f6553cd44bd97123cf94f7b6bc65feac1422c2a714834ac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb6283a7d7a0e4d5b316581f815169e7cf0c5682f2cf8f46b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haab7770831c82894e766e4a0d1c5b6a865d2bc6e16b0c5990;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17f55675a71f68632c54ef4a598bf9888e138116b0e85d831;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he829f4660e46b4fba584545a3b48e190866a2a0efa593b823;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f7192418ce99203e4c1f0c19a7d6801f07e8b3797775dec5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9fd26d184ad44f895040e4f1a8ff39139d2acfb1729db2aa1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h669f9e12fbc73d7824e00f1b0db1dd4ce3bb6cffa7c841e67;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e4c8dbabe3af2fb2f36a58d2d5b270f35d2e742d6208fb04;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b96c03ec7fffcbad6fed1cab89cbdad4f325278e39f0299f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf0d194b899ea4d137cab8dcf39cec0fd7bd295c113d2ed7dc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf54660f8c8bc4340863ea8b777fc73f0037ed40523cedf571;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed2996755928ad9febbca677f128a5e452d6127546c970ae5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4389e4b35a8286685100cd1598e688b497eb82b873121e1b3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14743e30c3ad2730bcff24ec5f36810d918d9f56fe1bf54e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4dceb9f628e8bf9f776bca9e7941095e65ded3dce9222d099;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h82a17f9b52056f83ce5381ab40568c2e41a51ee1b50f4c1c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3540d12a48550eb9c36ff7851ef76d19a5c6d752cd4890dbd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa2623f3967a82a24020754ce6e23e82b79ade9090bbc60f7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haeb8cb17cc09d69d8e5d9c50ce373a0ecc663fb888d93b7c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h15d58a7d2395f63fbfd54d158e2ea693380713256490c359b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcca4d2fe6baf83a76141f47b4e3a045f4c3508a4e72b35d9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h14b4ff9a459636241013df9ebf41f497692a2ce30cf7dcc9d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he2b03cf35667180e6fad176bce4ee845ae6f311c204560544;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7098a0d3361e1286e6479915c7998a565ee47ef251f9c61e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h120f74de7afb64430ec3992c451363df21c71f13ca79e6b96;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda2f2401c67991e99e13b8ef159126fdea520700b3f6c7914;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89aa89522dfe658984457d5dcc1dc3ca67631b78ed3fa7bdc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b352afe94eb7d4ec898ac807835438cc0ab2f0e7a911d52;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc10021154d75add85b625ed0c8ded1cc98c87f8ca481b4b97;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47a4bac1251b01c3dbf6e1c32d292c3e66b22920f6128a6b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32afc53c880cc80102f2cc677e88f47125395110e8ca5e418;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h217e83915bf134be04963a5e226e19e1905a11711d33e3e57;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9ae0cb9f5c93c7cbc3bf5f560af5b009eb3a74ebd85770b4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9dc0183864d712e39fd597d0896414192d5dd0765b0dc33eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd3b36bb8939c14a82af73e74ed6bd45f3c1368585258892d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h81a42d0de3bc44acb2bea5783c8a6e4d1b7416863091f99c8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he8614a80d459096f420b65212dd1b5d17be14a0ce3d0f34fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd81e30f6c795756b9093c1f9c3fb5cb4a660aa6af10c7c86a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h593f47d419008f0480749689f320ddf7abac18175f0df4f82;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4721097f3987f17ebaf489ad7d85a7a3f0f2be6d87630034;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he39cffd36eba15a979940e10f554fbae1bc7f8d7bcbb5c685;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3fde76461335f272bbcd6fc20b87a8042989d5c3a27d5f23c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8485dbf9b7149d8acb565de0608fb31baa5753461fc85fa43;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ddeb28c34bb70b8f8d3a644a2f6dd3890327ce9338a2e881;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0e08900d8112018b7e87f0d22930162a2f01a22824013d52;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h251e78770762b317ff4da239cbd18c559cfd386d32a358a3f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf3267d5b3e648137f0286b902ca91c629354e8d980d429bfc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4cc0e8f66ead6a714c5476a470012db2f46a66c6356f37d3a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20f06481ac5dd47d7a70070270cb49bc0798e7501742e1317;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a815d01664e59e908932070607425889cca857aede7a5bd8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ed6ad004740f55a4a9cc0a1ef63b22e65254013074f856c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6a8c5c3ece6d9c321867aa54a5792248bfbfacc672765fb61;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haba7fa37cfddd5124f97aa73071b99097384e976f22385ec7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc6764cfd4547c77348b1cf680569fa4296e597a806334dc65;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d479fb51912d905bf5b8bd715c5276870d928cd54ee3c10e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71cf90913e7cd44ba79243b08ef5e813318c24547c6072769;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e4ffe22a022a59cb454e0257634fd7287cbb62b6ac2ba44;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he8d0410c53d4ccb9b8ac95d50e28eacf95a73f097b5a5bfc7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8117d7e65ce23e2d1d67e9d9938a5a1767c909c46050b54e6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h97515abe03336b8aa21f01ddebacec63f9e235df498ac85ca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c83b8ba8357fe0989e2df3dd0abf9c6e09baaae5b51c18c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86fc0ae90b60038b1add057b278ece5a8e52725b8109636a6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3fdfc6c8f3a91046769caf1286758ee08e6c67fc9dafe6c3a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa01cb2f661d787abd38a25d2655a69f28192a2f2000563c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1824d5ce1ee4b17f9de275053120d1f417e79d82e8a3daab6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h96fd9d21e9a2792f39c7c10a5ba4b32246b25a66c5f831a47;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef94cda5a6f11275ca64efa40685a64e3f3bbc4727dbf909;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31be3cf1903fe7972995d7acabf2aa9b486e88a004b09b4a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha02659bdc4b0225119e3f2da237de28c80a6ce051f1fc187a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2dc1d1a78344c4509bf198cc852cd45a0547cce2483bf224e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h98312a3a1ca67c44c5eb43dcf508e3015ad38f6da6e878683;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90bd2e7ba8c16f5d2980cd1e989e483d0fa2babf7054736b1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e237176022a733bd3112146c4bf87b9f4a8ef081e90d453d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd063542e43a5b63b8d70148ea31b2239201760d1814e4ea08;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbf13294a4398836124e66f160bc8e1c76ba5f7f26416df5df;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48c478581a8912e3d2a150541c7e9fc430f40abce467a559d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58321fcdc7e83ae622d189bb9478e1b365103acb7b63ae7b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d0c486fa7519d931b44f2ccfeb11e735210e9db2883d2228;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb077e87b4af66aefeb4a9dc12db6f3280dee92e647c49c806;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35d0d7026bcc0e067d901614ea03c452f7e2f228c0de543e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d4921f21573b4209e1d4b14845637ce1c875338f7c37d3b5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h299dcd8a451f290356f1099e73c0c190b7e8034ef9be9fefc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha48b8c16d78b5b9552ae030acaf09a64d3948fdb1adc2c01f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h71a2b76e197430f0e2ddffad8318d2f3692525018ca7bbed3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d4e09e75e9a43494c0b9cbb90fc4e22090ebe6355089f844;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70e8b1b133d0765735a111fe4f064a2257aaf0925700fb352;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6be385fc100e62177b5dc9ed67a7d4f54a4b7cfc2e64dfdf8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4715fba743f62418e5836176ef720d92816a0b8c51fed41fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfb932a45e93de0a53c23f6ceced92bd2f8ef35a0638d2bed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd7dbd7e093fe6acfc26a8fdada824a521ae40622a1e5a5fe8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf15a5eff2dddfb82c1a49eef05a85f1d7bcc037614060b753;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc91648ae8e8cd1194365e67d3058ff016bacd305bad96f83b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa37d2ce74fe3d8d4a964685b4537b314569363e4cc608e8b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf65ce32a629d2524501b841fb56b2f6e0ad2db59b5757e9cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcaf11b92b33035899ae53ab06e9f4d48736e3157de73df578;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a0bd7a4a270d3124e3734c31113367b5c75bf7b6ccb39dc5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfaebc9c2e72aa3c6b51e6a494ff1ab7eb490f68cb93ce90ce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h188b4558a41c1d3a919c32b5cc7e8d7021e6840f258cefe13;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc9fd87903c4956edeb1c1bf132ff3b6a9ba5e3804ec845a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5146bedc6764c022abb2948c3cd88f04efb3367cb786e190;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha10ab04869ea66402bb9ea0f38301d86083e432f41dce05bd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he41b1fabb41c40d4c6ce489b8209e4827e550b16ce3ada9a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8c6f8e5836f7bed587d868389d44a96a712546a562b26581;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda2916d80592dc66b3e82f38e222d4e524c04bda6f6be6089;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc444711f14ff31e00ff089075148c9690506246f46f35cddf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd3b578a3ac0f2224bde2897601c519b6cc7f86e2b006e59f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb2c401639d86a3943b2bc936d4405c7b3f2ccfa2fce9c3548;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf74f15b03aa91c0f53534bc0f7942319a458e40d68a7e3358;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc7d859fd2e8e22eab61b2a9c86d0035b2cd6e2dea1967030;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf21c52f2d7cb6ae36bc9da9c0cabe99e3912e7de44e337833;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha18975222f87f0bb6ae94fda2110ca98310eafca2abfb4801;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h77f81ee5e9e6364a8d45f6a30d6ce4e6362b2ed3109a0c588;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb89faab778f99ba13e8b98c35cc298603b527861e5a74aac;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9319471ddcc251b37a56cf2a9c1cafd2c22a8d5b3bc836c4c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h741e46518ce1207941a19488be98542f076550de2e7e9cc6f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd79f65f9a154b71a94ebcf9d90af7355e07981aae20605fb1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0603f44e516765e605dac8c7c0abf248ba25e878e74a5f2c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8b38b04fd1e81d6fae8f59cc352eae08e5df981a66b803d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a0973dc90bc1572ef171d9c169e7b24362c188d8a557a7da;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h31754228c68554012d8fa6f4dfd680544e0c500fed6897566;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f328b68749ac31aa3402f3399d298085b04f2b3bb6c8f47d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff107f928465a30053b77039ab9524de57d1c47ffa5525eff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7bf00dbc79bb287bad6619e138a2ba58d1724708cc8be2d6c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1bb5505f54ca60eb69c84924b098c1491986ca26fa3e74357;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee6c1342c60c919416212ce84223c82e05a76df62d0da6327;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d386ac2dbe548d97a998946397f921504cefd75bd76541db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3006b2dbd9ba4797242c5b6268274e7a7339e3d1f7c6ef706;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22f58247f9bec0283a238814857f5c9fee8714a1147c646f8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he49cc45534f6b3aaf7cf2e849019c91483f85d2ef76d0725a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3a0c7327ee65e1b126f9f6d8b4574ff98783d3d4edad438d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hae3ed2c82cece73150bbefa3fc0a12a2e4ef4b708fa22d93e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h683346d954bf1a58f7378c8d806418f2f43900f493e718cbf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h894ca922a1df3519a7e1b7f744f66fb21e55c1265b685e79f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6ef20417c8d3dce91326829d4dbdf500e281fe483a9d485a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9fb96c6f3589f1dedcf15f7c36b6300fbfcfd4456cf2ed6fd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf659ca79e6c52aa66f5961c5d45a44463af4ca4b9f95dfc74;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7cc9215ae866629db3bcd0f274ec048e49f6b791b0facf3b8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h73ca1b9b18025740bef2ba3327d10541e1f79cec2651c321b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5b9fffbb151fa2b817ebfb91ace5740f370bf22a4bfbfa53;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb834a47428560120b8fa31d47139df077fb8ecbf218afdb7e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47f1e186b7aebce3bec615a22b3514bf4d7e48c87d5a0d156;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba4f55308d4cfffdcac80df0567fbaee4a500b63f71c3e4ad;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b4868d3d81d2396ce439f944d189dfc713880103dbba5992;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h97ad590185fbb6a70e3eb7ec713608fe5bc7dec4942b96e0d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e811440dae37167623b097ae8dab869a203351b3930ed0de;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h559902649077a1537133b053de8f69ede0545add69a3f06af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e3b86a1e963f9fe7f6aec978bfef9a2aa1994492fa805839;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcdd5b550c75fed90fe06199b82cbb32e1967d2190ac288425;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc81cb2873163d894b6eb92738413792de267117d4b57a58ed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26d28d919d8e0deb513ebc81f5aac05b795f1b3997c6d3bbc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87a99c573292a444880afea29edb99333bce4b2b50ede8417;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd5df98da6afbe11cab16d1b05c0a6e3d0c025a2c5641eb11f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c64681bcdc313e317c9544ceca5ae3e8713d0fa550757e6d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e4799f52ae449256ccc02a55e69385d93ce5eca934cf527a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h30f4ddf373cd469b2d64a8a5923f53c529d39ab47072916b5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e198751da93d53f3bf78f1f9e93a677aa9c180542740ad54;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5da662df900c6ecbafa7d7bb090391e9489772de67684b5e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0c42cb93f139ed791dbf8ecab2f1659359daa359ec83c55c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd8937f75e14a4e629f7c26bcb1951e65e0c8a58d7b2af49cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h48c1b72a937acb67f779b1bda1b79ed7d459036c9783d644a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d616a10ab736033bd7bd87cc5fd4b1b58628d15a9f3c45e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb909a45c1e0adb9c79a55e88c23b0cd7ddbf0886c145a98c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d230d92926b997a5d3fc2423052d50159ed9206374da6f05;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde61e3636107565f0fd8d9d15e1130cb41d4f83db752bf1a7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2bcc63bd15ffeda560e8b295fc2597dac5c0a0551cf815532;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9489208b66fb60bd2ca078944ffa460ffba4fff851bef8272;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h402eae1f5ee12e208a4c39fa9aaf11c6f880566e6d965e52c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0079cc842399806600f704a16c220196ea33c17802900486;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h771078872c10b450a1457be7431effba74386acae934759d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4e4dda037e83433fcf5cd25c4667314b017692899e155e83;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f1dcb29d9450ed8b7232539f6b741e406390295dac879841;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h19bf22c585650cab7a81373b73583d24dd068fe79ebada8e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9b6f250111398b3fd17c549e45c8eda28294b9526dad148ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haed3bcebea17ae53bbd75e54d23781834ccb5c853ef20b561;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8bddba3903ff9099671d5fc5bafe7c0d6331f03a9604fe810;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0d4afad4074e91cfb2e9fb9a0f693455b8c4a4fc2e2771b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h511169b402377cda3862904d58d354491b1e1ff7faea8ca62;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8e573dbc6e12e8c03e640848937d9d425ca9edd8e7ab506;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3d888a44c3563544dff7e135ebef075c7c8d222b02db3a350;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40777aa6b03f3060ebf5abceed81b0b5e8c6233d78e571573;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49886c9a3b4ebcbc42374d75cabc2a365934d91bd36e055f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha5090442cd5ffc576e91ae1e91d6b115b821a7408e15a9940;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d563afec8b8d93c8b2b0e7cd1c7bb807fd767433daff4329;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he1b0c2d73df2ea59c7714dec92f5fe93900f5bc2cd1c3a12d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb6b77d4fe74a735f4ccf75b77e8df3736c06d14bd819eb8b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1cd8ff2e33533552e8a70a69fa2e72112df4271f669d80e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a2ef2ba66c795f25e8a9ca7acd65053f922e4f4dc6e18c43;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef268ce02004c665af346dc7c10b9ff774cf8319dc4a690be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5e880113e813d3f5cd8c4a89b52fc776bbad8503c9706dfa8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h160b478f7cfe5b2023392d34698ffd09524b4260c4596295a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c8d9fdc58aeb884f313e75c87abeeeeb912576650dc27c97;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9698b018793e79df8df989863670f8ef6ada6ddfd03d76570;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h20efaa586e53a5a04f35ee67af0befe0f9c302f66a2ff7208;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h205f2cb7d272642c3b9acf3d8d1bc08df2fd041ce7a0b7ef5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbe33a419a48b8b826af9da8ef8fbb96823b666aa0277b6c58;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1191181c0af227e2882f9f800740e01e3fb98be280f92c7e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6144064f9b8df8f63d11dc2347d815f0d2de8ae1f32797c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68b8ea5334d36d4be9bd82e8d7b26e31c6222ec90e1f60277;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc0bc565eeae8e3568e8410780e9854eb9c4341e387e5ec86;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e3e1f6b73371ae6c3358593cd2b394754190b6441f6531eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3b0ddd9b6359cbc55b42718ef3a23e149f415327902f7bb3b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf34b6d8915dc86a65d75534de59dc72110b20484b1ddf78f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h59ee448aefd43005e2c7e66e8b9616e47af7297d51d79553b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h133f772896e3920c7e2194b17769091d830dbcb246538b868;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2856dc7a54c73157ac4a49726cc35d1fca906d2cc2fe3d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2782c2f2a62e889874d652adf25ace31f6af8e955d9ba01eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h61ba3861958990fa5db947213f73c329989ef49c2a9048196;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h35d1eb255baf6342c059527ae1cd3db5dde1523545669ad3e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a9088030971971c289aef04481e3ad74230242a4ec001b5f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf35c503a8ece6abea4c6e620508a4bf1c39389b15df771095;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c040361230d2305be8eee6fb54bd576e5fb4354cf81527af;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4fac32740750851bca61e262a061b42898f19fc18d215bd94;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h37e0c832634ff99d00a6c3ef6c6201cc6f78123c522fecffe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h90b6f0c5c6e3bfa0a1aea9d1e19a3e1e610fdc2cd1eeece02;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5d2c39dc282b4b169e462d8ed16cc1df0fc6f9c48731102d5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed21ee2febd602f0d1819b3756469745c96f574b76d315379;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28710d05f31d47b431ef6fe0a20acd1e35b2bff024d9dc4ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10efe156544c8cc564f9f9d31e5dd8d99382048ff7d48816a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h36d9ecbac0bc8989df98c528a1a7f36153db75a46c5d6c840;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8087d3c66d0720945966f7be323403f5cd474220bf9700d48;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hce2b9f9d5491f0af185b397e92552b4ca76bb226f9e0d5466;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1b6ebdf1119c478d60ab7882f7f2aa2bace11cdd5177e103e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5dd43b40c4821caa5e4e63f3c4de419e8c8c1bf3b3c1dd336;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1bf73f441b3c00f02cc5701c97353ce548f9f3e1d71df554e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6fd783a1451ded216ca3f04903d84893a00b0c75283dfac4b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb03b3c2881da22742f55341a02fa55db1d7e4290565814c91;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3813a3a655b80477387ea09d6a51549845324e946f5219b0e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc9446be3bd6bec470ffcb48e0de4c89890dc63b5d02ee9eca;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf26cec6e82ef91898e80c0f820d96ac79c77047494fe86960;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9ad229d60288572b626c46e2dd46263e161524752015571b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9fc4f52d5bb9178ab9c7b72748c8053b3b13e12cbfb8590a1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bf0d7b132c7c760550b618ac03d97d1d48f7d203b94b1d8a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfbea1c8f2ffb39f1723509b97323d8bee76e2bff2d20f72;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8a2fc718ca18564fc46890c3ee12e76908436dd2155e70647;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ba5cf0f2185ac4e6b0e975d3c7e2940d9ca739771ffc5bef;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h17640344767a41914583a2b0a1a575a57e507b8fe70a9f8eb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h67a0c7c04380ed9d5e2749b940b561c797b764c3c757e63ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb7579ab2c1c280a4c8dfb7ecb6d39cc452fd4f7223498a0c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5ca20d63ea573ad6493d443e8447f91bee304cab003178c05;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0423e1cf6625921470aecd504778734971d31cb159f468d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32969bea3d8a315ed4ca4ab6c90dacdc251dd6f31bee7f45d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ecd081c4a6c41481424ffb791d347f89a7f9916a0da06d74;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h89653a9b35e16221aaa1a42d6fa7b5c4c6780c48a14ebcfde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7aa66e37ffb9e04f2471e8c99bd3b476287bc4e9322fa9d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heed14464fbd1cb1186d10365c50976eff827ea7506b71a2f7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba03d42c10ca07f700f05e2d6e4ca7b7051527002aa4ca9c7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h823c465bee3f57364ab1b18d2b54cd9426bba96a179b35218;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff17ea1acc35bcbdaa1fd88e7bd8adb97e721eecc5dc10ab1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6862a92df851bed52bb258c5fffb701308ee1cf47af4604bc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8bedc3253ff761e764f712f752817990d0b8dbb0908d7b8d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2432c3d56b8fe08dd45c6740e6650117743cf2bd83f20630b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf128ca570ab4ef3a5e37bc1b4659286f9030e9499e3cbbbdf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5752e3a851c912f20eaa01c026808b0102648fb0f4a3c7403;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ee32803f9674bb2835b976e081c2ba15e24bc1c30b29aaba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h645a1d90c0953a20ba71cdc0b3d52575dc816bbdc3ceb3e24;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8ce5297c22879fe21df9c0e61988db5562793926cc94d9cec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb292b70f797e8f78885d08aae756c055edbe27b0de2d1161a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h92aa5f0bc38a34bff7d0190dd8acc64d595f5f1e09b23c6f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7e06ca789cf5ff290f43e92f7e188b5ecf5db93f70fcd383;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a850f4a004c4c9437b45b287f2b7c43a6738c3883c938ab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9e1a197e6096b3c3f70679c6ee1949de33246631e0c455246;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h333f851c12ad7e06d6ffb23f1857483ff43a790f343eb24c3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h99df39d3979e6fd161f14fd21508b69f7b3be1b14ba84ac57;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3da07f650be0ba36c2a5c836f5f87b6e4a374c1ac6dbc80cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h74e5aefece1f6a8585457393f0a9101e91cf601741b5da5fd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5471997c6290900de7dce55890a5a17d60700ed660211af79;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1feb9efbccedb32c0da59d1086b682e9ccc818ec53c3238c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2768bc2c4c9919ce11bc61c0d19cd98a7979bcadc71e0a26;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h68db715a8850027e96dabf618b1a5cd51d0e332b0c364b64c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc18f7bc567d696d45fa22b57573703bcbfe7d277c12b7e3b0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd5b0db4511f3c240344da57296dc517d857e5106ea5de423;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcbc883d8c31e31b457cd4cb9816f0b38df60473991280323c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10144a44d2588b9839245c8c1f8a369b0824bdbdcb2252b77;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h64287e138d56ca6599dc043bfd5dd19ac7d66df904b70fce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h277dfe06423d3e36a8544d35d1af37682a100be7fd6a1348b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5c085a583a6ecf7b205144ace14c43a1ce2c540929d394333;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha43c0f0de8c83d76f16bd14c6dfa7a21efcae7b7f1c4f68b5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he867cafbfa74060b523c0bc027c30412396b08216483e9349;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h924dc8776f8f3b9b8d9e5a962482f4eeb8393cb72a42acd94;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6865646eac0f3899a64f9741108a411af07d208c455f4630a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcda75d89b75fbe64683a668d5a5e363dfbfd247c6d589c4aa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7794f5705b0976c6868e8c199894d0d76b275171c8b97c7e0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b2bca10d57f197dc21f0e7bd6d25682deae721b738ac22d5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h846e245da29633772e6a8638b75c8eb8bf4bd9d9de69b4d09;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0f7cb5ef5a194767a646b652a1e49685df5aa998b4acec66;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6cab87c3938096dc77d607eab70a2710b1c9d3c8221760347;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8534d1d6e4b6150d704523542300b7b6f4697a7ac8e18be2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47faba8ad5c64bb720733a325e40d3fec4188a235c786af23;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26c8f1d263e4664281db709fb0a0cf5ca9bc627bcd5d90393;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h225d514de3e252774f33a06ece28ab900b62f8723091f5301;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hded2cc7bf4ac8f238585decb866cd0cb4bd56019d4db9386b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h801c489ecccad93576af13a1dd57b1a9bf707b16757f14773;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hca8c0bfb1ccb7e5b8b5f47c9c94c1fb812427bcb742993d47;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd096009d2722f69fb992df449ba3860eff360638f27f7e650;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2380acd1cb80e2268b02cf4af26c54e8437fdd5a41aaad2dd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h64b95c7abc0ccca3ee47ca076c3e0e85f5da7e2c12c9e6d0f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h49df178af8f8257f827889f1bbead5e97abb7123f1861129f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he93dfc3f5e39dbb0477b50369bd5d485312ccbd0a8bc33995;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b57274ecf4496de532d54aeea844b2791a82653e1f0eb008;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c5782f3b68392917be7d31bf7a13bc44e8b4511b4bf11ceb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c7ffb09b1a8bd84d46491aa69268058ef3a2209838e97d11;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfc9c77b5deeed4f375e033febbccc887b6e6ba5c496356aa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h689500fa33dc69b3148f37dd116b10ad9e83d3dc2d83b5481;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfce3c87aec7c7f50f3a39496126711eb58129ada9bf0fe7cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfa40f570557a239f48f87c50c351a3e76a692478103c035cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1e72ba34d49765a887a67187bfb90a923087a0337fdd5b11b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hba13573d292d0f61bf600de25b2ab21a01b5798d8abf7a48b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbfd850b8cf3c45c3690317a7463e53bfcf310c9815d6c19bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1739a6062c11c1d8f32891f05223be28eb9c95a753007cdea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb24242069481341419d58f602cdc3731b3fffcbfa049b9ee6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a72b743493dcf365ee0cd0f6875b5b061bc1561fcb019ac6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4c45793154a210b5991045272a1c7e2e96b59c0006400f4c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbac8e35dc7fe131cdff097d0c99b09d723062fb5141c787e5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'habfd7da1dee80fc4680395d508ac4bbee5c275cdfe2e488bd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5468479f192630dfc24cef0d60dd565bcd5adeef9a0b7922f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c5181d6ae3441e6e06386ef9990f96c950f39644114f28c8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf5a1df91427e1282e3ac89e50fc5f381b5b832e0e3d7e3673;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0330a1e2eaa42acae172ad08f302c035008676191cfd18a3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc09445416d1c9b1d478ce71a380f57e7dcbfaff406f767129;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7efc83be09f144061d3e24d345632e8cca8f3e28a6bd1dc45;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he8b5a8a02ef7bc48f2407733d49212b5e98bbe338f8fa7bf7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4e649c0b8d0b544bfc8ec4a211b4b9ba63149598eafff6c1b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1d71c25c9bee55040b6a1ab264873a01c7feaf1c5bfa0abfc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb6a1a09ae8f97dc39327a46ee14951a0194ae2e78116e83b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h64ab162b318f1ae222ce1abd01e4daa669db15acc3bdd76a5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h63d3222e45557d9c5fda0e902594bd21b3efaa9fc7a5cd9f5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he5eb90c8549d93ca3d36f3aaaa7318c7c9e55b2de9c4d5ad6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94cf2e95e2e468a92369f3f2836ac305e9af8e9acb6833d70;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5acde26fff702f722166e1dd1912ff703279b611eab1d23b5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hef1d97575a647d081becb182ec7905840dcceeb345ea7148a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7f6f2674a62afd7a131dd7e2aa14aadd77277423f604196ab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4cf1efb0cb357a9478cd2e9c49f4622cccc445202721f04bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9d986f4d0eaaaa71d1a4e9a677900aba82d23e22c2b36f015;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heaf4b63ced9b786382eca5467b0446f2710345450bf489e51;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b26f65b450155be7dc6f2e3d68066ca314f66a545e37f1e6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a2446f8822734597b9713550605c82995b737802609ac02d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h40a7d78135d3a94870ba9405e22cabaab10cf857793cf6835;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee87e0a4efcd621ba02499ba71b146d0607a8f2605c78a27f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd4b08a6fda765a5f18f2ddc3a15cc053f079bc37a64eb0729;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7148bd45a1bffb006cf7370250b8022f09a1a854d52402e49;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa0e1fcadf51f5311fc5da458d8909f17179d07a07bb888db;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd50b9778b2affc383548da83e406989c565294f7caa681382;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2021beee863d153daa29ff60f6cd2ef181a6bd05e1ae061e4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd141082b3a830c8cb74c705a0da013f57eec98ed91ca1523;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h94360ef4481d1617baf08a62fb187c50cfe87507f1df3d667;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1dc5ded910453eae0341ea7289870afd17e3532df9b13268;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bbc4a4668f7a497c4df7c212bc3ed3e2c8b22f246e80584b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h628e8a14feb7ddfd26d540efdaad3a58a5368a8e69f0dbb1b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h26188cbc2e1ad483e86d7752f402bfd5aeb5ca7681ac08f88;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa3ccfe540cfa3391a86e0c7589d0095891f56b0c73bb4155;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h715ca8d9a5d7506b0bba9bce27ab5838900473caf22447095;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha7a03b961649524f53d75757c40c705016d40d5bf70b6ca1b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32a6bc10cd951172f185f3030d4862d912162a346be36c57b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16b09dd5c5be829cc03c80a4397f6569a06bf6571e3c7cce6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h201b054b93b40aadb4c891544375d378b4cf91860b5cae946;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a4b4ea5f3d611ca678b74d2bda7db7b71fa5281551b62070;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1ef0220eb42bf89a322b40fd31416923ef060b47a8c4075ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7b8ca104159330b5eaeb3068bb448b720b079e193bb13f610;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h726b319e05d7927a04abef4a9886402c4aff545650a248b5c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd9ca04d7d65f843732fa2cceecce94a3cd6ab460c352a04c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8525c939d7c7c07ffed7a252ccdb0aeaa3aa255ebf9df068d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h50be8e09a6d1eb21647b99d7372bebde39aa9e9987ace54b7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a7eb00cbdbee43c5096442d0637d8e71c445385822ace2f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4db90ca36401035610f00fcac60ce03247b70808784f740fd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h58e6536b66e44f6964ccda78dff3edf3e585c5cf735a346a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h947ac1aaa59a5a821dfcd03ec0f6f14d576d32da04fc82537;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd0952ea858ae2e2e5413b0a81ace89925e10537ad2f4ff7c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hff3dd3144c00543de006787bbd41c43068371a334c5288189;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h32d647b6f53cfe7b9337230eb2aaa0a3087af8bea00308c40;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h36cd2f3e6f09eae38a87959d689062075a72f8c18762d5811;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2270b68a1c3303cbf9e30b8d3e68a3cc05ab740e2592ecdab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee3e3b54692988e1369627d0d78274e5bccb6d356840b5bdd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h115bc6b2ccecedbc4db769c4b7dde9dc8d46c048e3b52adc4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd11120006b8f42632cc8b7ed8e1030a1ca640810087d702fb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha17500cc85ac83856a3cf3ca29b1a969cbc1c532456f1d5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76703dcf361b75add6afd90bd176e7cda53436c8e2e4aa0bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h93e660d9bc1e6f3a7f5fc7b21954a167ae5bc67a61de357b4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h905b6ce64570d9e9d9b6d18b6aa49c8637f557f5b44a40a25;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb727509961084109b98f65bb7f606021a535467c486cbcc8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h270f5e24a40c8daa65bf098ba172ac75a0fbb217c421e4c78;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc81ffffde55500db99fca94bc9564e74d7a2cc56f16e256c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1f47cd76b080624f137ec02b291396834099f31c42ffe7bce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0349d6f4ad721a9af368922bae3d9511f9b0fc38a09394a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h767859fd8809450b20e4121f8f2524afe452c838a244167d6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc63e21426316c120b03be7e7c1a9c3f49ddaa057ee0560bb6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h24deb2de60d0cb91b8fe33f4c5d83ea6739663ce9e46c18e3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he4fc98679563b5021be161d7cf50bf5d4521b0bd3458a11c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ce9e2c131bf30b357d0e49b8240977080910ae6825db6d4c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8207c6bde210d304ce7aa127c93f6b3202fd5acdecdd708bd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1bd3e5df4787cedfb2a4463260eacbfa5ad56b4da60c4690b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha9ddac908bf43e1adab6b8a56ba16f5ab608031d509951762;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1d037b23f092b26e239f8bce00d2797d4763287856ebb18e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd421a26ee261131299323b10920f3b0c92c4cd83cf46920cd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb8b64ea3300c7e3416abf17734c3183b3754424f4cbe86a74;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb753ee52d18a9e2fcc7af1f0bc420bdc487a75fb36c376273;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6c5551fe1135840b306c51c7ea92f39fa5aabf8d2db1cb4a8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6f356ad97e849f8474db124b0508a8ab4151d06f1e78b48e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfe0aed9130905d73a6690108a499f0ea15f75348792c62cfa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75e5ab1a64662ea4ad4b8388b8dd378787cda92312956cd73;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7cd7ca0bccda9c8cad19f83fca929369e8757d9dee538c5a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he7df393876849717cf8ca40649fb11061e114918e8ddf6470;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21055a540ca3cb93cb2d9143e6e9b7e6e94e7afca388f3f67;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1a4d8fb2bf0d040e06b2640401f51c3c28270a365836e9df;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86b5762cd232f53b5525e38a028fa9de34b572fb2492820d8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h64b23343862381b7c759f166a4b44c04ae17c66b9ece9bcee;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8b30977f2cfb37a7b09e6e95feb5b4e387a332663c0b430e7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8336a201ca77d3092c2ac7e62b3fee26f86af6993d9e52ad6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb56dcb4ea3c12d308822aacb94ce5f6ae39913153fb94b78a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hde165d42bb077437e82c8e0f2172a9219fabcfcf71fffd63;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h461793c470a695f0fd327c2e4c942af415a049691e483bda5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbb8cc5115e69aab9709316a0a9bc41015324635c623d657bb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h108c4b231392e972918d89b637da46b11b85c0599986dc6c0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7d653a481f8ad5f034abd7ed8b5756e21afe64fd00f7a3306;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4adea6a651bf53d1156a244f4805da920573746bdf0ce458e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6217c4625b8ff500ac5093505157c8d122f963c9df6ebda35;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6d22b2e414ce35db750d08363eb1608fbfaf477fc38678e39;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69e15fe89c660ec60521d11ceef02b05a37bcea8cdd3f4f5d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd506737b960e14462a95f0469833e076b0a53ae77a7675948;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he8b0cfcafffcabdc03f5fc7940bcbec4399be536a1a0bd70e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hccfcef6daea80f1451872d76b1c86860e0db497e13a76e882;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4f863d540f619627560fa9a304e99c44604bd78886b522f63;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h27f2a1d6bfe82332ae0e16d34ed349538c8ed1c034b4a7cf4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18459bdfd0d01737435e92d54c9a2e4af92580aa19d7a9b84;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he3e804da7db121cc5bf077bc0d8de30eb965cb13086fe0ec2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he52c2faf3f6b55e53e01e4a0d7d7c58aa9fbe0216cc19355d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa6cfa830b9f980de1f58e0e29bd03f42531b29ae57c77f1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd479415f1e022e2f0ac34afbea0c211ce06498621b353d0ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf4321db0969e025217566ac9d5f305ff33d73ec481c6e1798;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc41c47fe0918f6c3bc578a623462835abb20ba19d9ff1c28c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'had49140ed937f15e7f2aaea3e824483f66c2db8025f4b5d14;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h881ec5c13b2dd20c9123abde72d25b7fd9cf420e94561c2e8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h888aec01519b9e92995e7a952a63ca9d8a26927cdc4f5f867;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8bce67fdd5faf880e0e1cb41ab5e1d36c5ddeec1411b4b710;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h953b4c1f8286d6ed43d7314f2bfbfec9dcd06d13318a8ad2a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h36318f9e3de25dfdd071b8892d203e46c062198f40e99c7c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3ca5998492b723ac1d717320ed3b721bd9a711ecb996b957;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha0c67403d0880024a80990c702e16c82bcbb3a5be8ffee9d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h47e62c8b3f059b1a92ef91673d01bac44a9301166422e059;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he92fdc7fcd23e5f0b48e1c4fd6cc9549d9c39991d8b820234;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h201710902c2b7fddb53209f5a011a8cd4225d7c70a8d391d2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha228471503687c3fbb9a3d13351041dc0a30ee47e47b81ae0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he74955509b9835d067bb9816e4d131fdf3b709699f2b0531b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heacc0f0983f3be3fbdfc123df2a6ae20e2a2b0ff039c79404;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb35b38887e463c4956c9e0003424d2fb53adaa41d41c0e540;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h214dcd67516bf74874b1183db0419676ed090cec3fee7865d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h60798d156e9e7b5d2b5a7efa83c057b53fcf3289500ef3195;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c94a1b1b74d133cb56fa5fde177177fdff932c4be20a7c4b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5a2f85e542ba9f24c72404c51f4c13b5ca1d3d272791d64ed;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86e22d5c8ecad5eff25804f4834c4b8c5a4bf168d5c127fb8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h730d915ab70dc4b3633f0bcea66c120a4af7d3784190880d5;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h81f929efc70caa0de6d10e00c1c476858ff04560a3a14a4e9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4422db380641427fbba0faa43132ff74cb64a91a48741059c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha953f2a5e418e0c5f7081a817ac139585226d3087720694c6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he8831c421c979cdb6d5b14a8aa250e7474ec0669df33d56bd;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3aae886f6d8781f066dc596696c6f13b46427d0ded92ea57f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha4b062c595391e1035c239ed4c2b3c6d7ad12fa4d39cd3474;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c55f183f3abd94798f1df2834e66fddeb1a889e16f33092b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbc6b72f0a7331219e47668f905e59450ae59262b7aabdbae2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h876265414150b1bb5da62d5b09d163a3e507da776c2141cba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h87f59c25c4b27d9b8ba477256a0c6af72ac7b5b8e5a2306d9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h178bd11795793fbe1c28181cb1686c166d2b4f0cad94b193e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h95cdd6568928aa791ca93b4fd3b8168ee5fdf83d7642f4dde;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hfdbfc39834a68ce59d0e3705d9d322795d465aaae614ce928;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3bca24c693c2285b025382d2cc006835d8a1cbbffdd557057;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c01880b36ae781946d3225a9000981b323e6a778ef58e22b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0b5c8286f560d4f6fe8e5ecd0a874cfeda04f1e1e790a72b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c33465ed90639b1b53d2927a4423c3a920dbcdafa925a438;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22e9df0b820816bc15d902d3a15ddbf58ec327ed66114b63;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h41b8ba6ffec231b21ff40c9ef7f0c8e27ed7eab98ddcd4d43;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd2e70ed2681d534448116d4086b82f344a7c2a8f31097b148;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha2658f44d8f81eb619f1ab6622891fe7c4674af4bf95d8b52;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha1ad5f45ebd27203d77fb35977d64b0ee4f43d585120881fe;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha280e3ec74d78c03babee0902e3f81ab65d12865131156444;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h16aa97a5091405a2de970707aa028bc83447b23fa3372929b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf068b161a7f980ff0257963a5443b2a9b5ff7d6448a23653d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e234bd4fb6664fba951aa3c4a854bb154ad670cb41d4a0a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9901dc715102741a384f1f69cc343e75830be00b96ac0e3d9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2dfaac6de640aa4319d9eeb768c7e3f5c4338783d8d17e475;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h25e580da6351260bb75bdb3176eed35db076284b855711c6e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h75dab96e0d8ba1cb931d026544d2a924adc7f6a56cbcf233;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d95391acda4679a8ef9b4fa6608f9a9a07e343efe2d20e2d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70b3cfc65b1c90f04d3066c1c4660c4251884733ff9dbdb7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb0f1db8c267dc1d713f4ecb67d903602c09ed693ccdf0896;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7edb2406be4e5b089058f79e1c76a68c931335b215a5baacb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h843d8ea335d97323ee9d8150142a05b99d261c0ce6839461;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdd25bdcc24a902b646f7bf6118499be27b58009779aeb9240;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haa3f96987ad4c60ce277cd038afb2d39bd5f9ce3439a75fa2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf110247477bb53ac473fdcccffcd501f79fc493fe0a25ca2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9fd8cb14a683c3ebbd317dfee1fd52c660f8b09e6955478d0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h587b9dab1da4576695180fd947c45c868c2e4228d314878f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcbc681c73e7324911800cbbc2cfa6f360b9ca3425577e05f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h468aac994602d2f952eaaa144f3525c9ac346360e13424f83;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8323dd942de5e14a472155377d65bc46ce78b00bcd1abb886;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h69b576984540d85fb0400821ddd5f42dcb2b0255586422375;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10533539fd7eb9c48ba4b93b2004db07b3e90abc27322a870;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha6ac40bb36b11a9b7a7661376b450cecbd85603676bbacd9f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he01675e2b6fb51b28f4cea5be04aa9f747817942bea5dde1d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he17fcf7ccdaab73099aa16978a910b2fa2248861fe82cfc7e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcd91ccc2f38024467bb6f9acc1fb3e3de467e6fba0ecbe855;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h872ea208c9bb56ecde634f72ab72c38602b33d53dc898208c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdb41007660f3d027dc9979f5f3686829f02fe532aa565483;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3cd00040d12bbc56ef142fea1d40103f5bd8e0ad4d5380dda;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34193ae246e892aae0f92834b3930eb8bb31813d9fbfecad7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c24941c2c841cd3adc10431c5481e348c5e5097c49b91293;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb96cbf5a9b48ee9550be70367ccce9dc8515673ba44697c65;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1edbd6d321491e6ef813c9dfaf4cae55c161dc5e63e7e72b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'he9be072d877456edac5a22bf6e50df713f03dc229cf38b974;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdf18e391ed6bd7acd98260beeaa217bf4da7cd8726126e82c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h44f532680fd1148040aef9a93d7ae3e3b91c2acef41f884ba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac18722dde7c6395e3df2547d1f74437a98f6a87339a0be;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4b62791b0468acb35d5b4d5593ba07f290a441481350a99d1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf25dd5e96e64a294a4bb5e676d4464429699ce47c7c4bce5e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1cab7f175db406ebfdb77b773f25cfb81c4daef0ff11b24ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h778523498234966193ddf9f2088d5e55d09d533363974cb91;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a50f929214b382f4d9afe6f9ea887dd058d7729a95d4fe62;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h28eb58fef6ac39bce39dcb13f2170f9c42c638300cd9c2c1c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8026b35951cc91eb12e38566664ff8a825f661b192618d751;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd9a6e4ce2ece9a824eaa2c1d1dd8127064a9189f9bf5bab61;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb676fa8cc8f871b08ff060277bd375cf2dbf09843c8ad105;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hffbcf33b400170e0b5db545e8c54149ed166e99df6768fa50;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h18417c0907024adb661ff3c1893d4d95aa4b52f1f7f739fa7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h822b815e9cbe557aafddd2782b52877db7350e68a3d5a12f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ec385aa2820740326c653b837a1a4bb4f1b7c28767ad4634;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcc12f250b8a1877f96c8790c298665f1477b7c16c81af8648;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54f5fd240e600e71fc486d323ec0df13015c4ccb7ac673d1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h854ca3092e377d20485a4d39a6bd330488a21b922f9544bc3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h246bb0028a9f63158d0553b1ab31b495a6d013a0fc3f56fbc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4ce93c2e433ae844bc729dfd1edb1cd4361539c7f93b97f6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3be4dcb77f5886507118b1f7e0b9540ee21b558a6d3855d99;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb0d0e77925183e2e073fc9539dc75d3098bd797966ee3ed9d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h11f12e674e050f6b4ec49cca2aa83d16271a4fd1ef21cf8da;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h65136ac3ec32a6a8942e1a9e9ecb708c83c0cff32689b9c80;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h380272466b80bc6fa2aeb49c8c9de6190e0bf031d9470d980;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heb0fadcece76839e2eaa7d0d9456637406211e7f6f5c9ab8a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6967d3d7049fda4a6befca24ed1e010ff8f6d27438d3c936e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hca85b6aaf240dea968b58b39c89050fcdede8572ebf858630;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'haaa808f31a082d1b794130ec982f5f9556b39dc2616ef68d7;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h439308df07f3b73e3738ef741f195e99b10c76e2e360a5bd6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h10a0a978bdefb3a625fa93a2f14cd0ce76523974d5baa7e41;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h394fd2c0519cd67e153db7548eae06327e6aaa70fbe5f06a8;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0397787484b436f256cb9ee4dda3df1001b20922cfdeb07d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h701f8f1cc0f4ec23aa8610e66f8800f5965945734cee38e58;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc896deac496834aea9ef0cce49a2fcaa66962b8ba602ccb5d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4f525ac539a4fa9aefb999531896c30d4465937d2a4bf09c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf1d7f93890ac98bbd2f6198ed492e1912b414ca6d32896fab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h917c48fa1072b72f10fcc34eaed7b0068457918759f2e67fc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h932df3336a9356ea29e346babb22f7c5ed7f56a8eff40ebf1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5b079461868e5961e276ccb4b362d80cdfe27e2242762b30e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf8d7dcd90e5fa5e93e65e6d08a1365f2f2d226b1e5fbc49d4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h70837af2ff5719d5a10b33270c3bcbae9d931311d9cca792a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h742bacddf94a948752cf72c3bac3de61b09a024def454bdc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb79134002150b7dcaed595b6144900490a0a6cc37cc67b1ec;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb5bf5a8493dd18cf36d4b147b134b023e59a968ea7bc98d51;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4bc135e2c52cff8f0df1a0fa638dc8c0952de8cafdd3e35b2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h88060db907b262d0eac4d3ea200fe25fde3cfa9d067cb73bf;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2c98714b0515b5edc1c08faded5f34929374da15db1e47341;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9893ea9fa54d77ac7ea5bfbfcbef0ce4a7d48a308709171f9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf934cf4386fa5f90b2bf57de24369980993315cb67f252e0f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4dabbd6a55502a285b452211afde062ab20dc57a2c3f9c882;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4a61e441feec61745df6793b92b566a1f0b9a14a9d0aefef6;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h76780e6255b79fc4a89e0fe8a153462d5816711e7c4d683a1;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h103b2eb5d470fc3ce69aa0ffc9baff8fd0fb1f88f04ffcbb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3af57577a5abc7e6a4ca727d4976eb1063dc8507cd4ac85c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ef9314d7eb0d4099a9aec5e65f66e93631a6af09ebfdc7a0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8f926a28b2d27f9b5aab2fd92192af2922f4899baea388834;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hac8558437628e3a48cb2fb8ce97bd9d1af8050d68109da28c;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd1d949cf0fc469612c6b4bd3838cf85dcc975360b44b699d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9601181a3bb63778072ed5a86d0de72437aed973375a054f0;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf93514e236be44552214851f9fa8e57db70e32c9d2cf916de;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6dc502b939382ef6842d7848eff586d991556153a3a8ce00;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha8e808d7f5a12e6cf95c2ee3173ec1951dc2a4623fd2db450;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc043b33e2fecc53cad76bb53da02e91006fa8a22203650a6f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h54652b76f0fef7588d617e469d69550cc792d378f2f0fb663;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcbd0a7307d6e1533e2068d6ce132194c16108d672ad55ecba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7bdb80a57a998f5adcb6a4395ec57c235f74e87773739768b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha33289eb5daa679a1d05027a70505a9efd74b603d4ab15107;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3f0f45dd82b283e15858e0971e771275cb26fbcfe44ebeab;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h693e009baa060011461e5a46ade5ef94abaac14259e1e7062;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9303c233d11b91ae6bd898f106ec6eccfbfbebae731d57b7f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2a30dd40d9972dcb656a40a44b981721ff4ff91170754d157;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc482ceae6261d7c24b1e664ebb12111a6353fc2f306f3fe2a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h938b73568850a5ee1b815e890a10d1ff5e8173c139d8e6013;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'heba99c1fb7f18977c00617351e41f592b6e612becb289b50f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h810f4c7e55947c9b42a0753c45cd0ec678144e64ccb59f407;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hd0bab3b1a5a8afd37283dd427dd8bdfdb50f429aa60d595fa;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4c189efaaefebb0811c621047b8d17cace8884e96c3b071c4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h22d315c7b962b462114e5b21a3da16c25e8e022b32428bba;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc0deea993d4bcd00dc5afad1d1e66d23e387e03660981a85;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h6e0508d27b50dd0eda9a8618be524310d39907c8f73134956;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h952e778182cc0d72d1fe8a0a119c86e22ba867f9f0b3f98ce;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h34f63c3b0f3b333f2ef128be40b461c539c94da90e53fc6ae;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'ha3775c12784656419cbb9172d0fd4b1699b181e07ee4b257d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h1295fee5eb16a72ae996c93792d807739c9384852bb31143f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdeaa78a83fbfc50dff478872b2c07b86cbdb98c8a697fa4c2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4d047d02ac0a164ca29df5786bd20a92869a39129085bf18f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h4da0cb21116b5a222060bafc8ae5f3b9bd2d723a31589eff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbd1ee66c419413196694eb9066aac958f3aa895becaf31c30;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hbed95e8352eced0df8380d750a51cb455351f35dd61f11776;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee169259afa5c2ac09bb801b5b722507cfb6ccfaef2f7c6c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h458f7ecc8b8476d986af9210dd0f9dffdbc8ac5b8d6497c9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h2e5077f12162700458ac1f94c5cf13508e5f67706edf44a36;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9a385543530f397fba1b2d9df1a83183fcc6ceff3cf0c1b7a;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7ec8419821bcd7d8c03430b488e1f103a54712b5cac07030;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3c99ef7b8d4aa25a15763154281e8df8a82ea82e9856fcad4;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h5db7d25c33748439935a7b791b3375a35dbc6069051cd461d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4ffd92ae3f6012baf53bddf87a021f167badcdf551458825;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h390418ad784b36eb5efcd3e7d9d4062f258ae864572a2bde2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h8d0b62bd74ef1b6edda7c49a2f4cae0b15ae9d5970f1f29ff;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hf7f509b874c0dc1039a3bf85a51ca6cc464ab48ed2f92b0ea;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hdbcf0d7f8aced7e605207f5da5abf935b59d9509381a54247;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb4c340f99de11c0cac05987758c05085ec8cf425411efa58f;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h3ec573a4e1a25b06989b3d1915c4aa7aec2247f5ade5c91d3;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hed23a4d35f9a5040d1386f25d9119dff81a08a6e2c3704787;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc1913e6bd9f0add756a77741b453e22784dd4b111997ea7f2;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hcf9c1384a131ee348fac8b25f9273ac076f4444271719d1f9;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h33c442590c8ce7e860827e8ff768e057ade8c80a6edac125b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb30f8e1d6c60a24b74214232a0b5cf015afb17787a6373735;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h7857d111719f31b2cb479dd31776a9a3be63d61926366804d;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hee551fe229a9375dd5e52b34ec46068a99831490d20f94058;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hda736d0266dab89a6e04bd4fff4104c5179144bb5ca94a851;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc11dcb17d8a6d141f0f7862008e9d8a08aaa4cde138b8c700;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hab03b86a5434912281dc11607a0d6fe71f438b1bbadf6fe81;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h443dec22c850568ae387a4d5d728cdf2c5321fe4e071fbbdb;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h21941d11ebd98adcae51efb7985fe65636755fa741682fc3e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb05d821453711adbcb410c629cd4b0d59f482de7627f3686b;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hb56f90e3496205905d74495cb2bb45b115acc396139bca9cc;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h9c229ec297aa8d4c4e9fabeb21e1a0336b7945d365459124e;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'hc4a55737ec6e5729c08e3504e4feabf91860de441260d2e00;
        #1
        {src13, src12, src11, src10, src9, src8, src7, src6, src5, src4, src3, src2, src1, src0} <= 196'h86f41e2a59a44114df28bc490ae8adfe28c9621fd3956a3ed;
        #1
        $finish();
    end
endmodule
